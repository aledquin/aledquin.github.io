# LEF OUT API 
# Creation Date : Tue Apr 30 11:34:03 IST 2019
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_se_io_ns
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_se_io_ns 0 0 ;
  SYMMETRY X Y ;
  SIZE 41.04 BY 90 ;
  PIN TxStrenCodePU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1428419375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 131.308 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 17.442 0 17.518 0.114 ;
    END
  END TxStrenCodePU[1]
  PIN TxStrenCodePU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1812219375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 128.392 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 23.218 0 23.294 0.114 ;
    END
  END TxStrenCodePU[2]
  PIN TxStrenCodePU[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.14288 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 132.068 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 16.682 0 16.758 0.114 ;
    END
  END TxStrenCodePU[3]
  PIN TxStrenCodePU[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.109212 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 23.066 0 23.142 0.114 ;
    END
  END TxStrenCodePU[4]
  PIN TxStrenCodePU[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.109212 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 16.986 0 17.062 0.114 ;
    END
  END TxStrenCodePU[5]
  PIN TxStrenCodePU[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.109212 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 24.282 0 24.358 0.114 ;
    END
  END TxStrenCodePU[6]
  PIN TxStrenCodePU[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.109212 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 16.834 0 16.91 0.114 ;
    END
  END TxStrenCodePU[7]
  PIN ZQCalCodePD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087932 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 398.009 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 38.418 0 38.494 0.114 ;
    END
  END ZQCalCodePD[0]
  PIN TxSlewPU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0857659375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 3326.87 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 15.466 0 15.542 0.114 ;
    END
  END TxSlewPU[1]
  PIN TxSlewPU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0857659375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 3249.46 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 15.314 0 15.39 0.114 ;
    END
  END TxSlewPU[2]
  PIN TxSlewPU[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0857659375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 2778 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 15.162 0 15.238 0.114 ;
    END
  END TxSlewPU[3]
  PIN TxSlewPD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0857659375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 14.706 0 14.782 0.114 ;
    END
  END TxSlewPD[0]
  PIN TxSlewPD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0857659375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 14.098 0 14.174 0.114 ;
    END
  END TxSlewPD[2]
  PIN TxSlewPD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0857659375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 3446.17 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 14.402 0 14.478 0.114 ;
    END
  END TxSlewPD[1]
  PIN TxSlewPD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0857659375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 13.946 0 14.022 0.114 ;
    END
  END TxSlewPD[3]
  PIN TxBypassDataInt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.070452 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002176 LAYER M5 ;
      ANTENNAMAXAREACAR 178.313 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 5.738 0 5.814 0.114 ;
    END
  END TxBypassDataInt
  PIN TxModeCtl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2177399375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 843.974 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 10.298 0 10.374 0.114 ;
    END
  END TxModeCtl[0]
  PIN RxModeCtl[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.634144 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 10.906 0 10.982 0.114 ;
    END
  END RxModeCtl[3]
  PIN RxModeCtl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.634144 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 11.818 0 11.894 0.114 ;
    END
  END RxModeCtl[2]
  PIN RxModeCtl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.78668 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03488 LAYER M5 ;
      ANTENNAMAXAREACAR 56.937 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 2.85 0 2.926 0.114 ;
    END
  END RxModeCtl[1]
  PIN RxModeCtl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.643492 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 767.321 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 21.242 0 21.318 0.114 ;
    END
  END RxModeCtl[0]
  PIN PwrOkVDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.22 LAYER M6 ;
    ANTENNADIFFAREA 0.02048 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.026016 LAYER M6 ;
      ANTENNAMAXAREACAR 1330.53 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0.3 20.27 40.74 20.77 ;
    END
  END PwrOkVDD
  PIN TxBypassDataExt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.105146 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002176 LAYER M5 ;
      ANTENNAMAXAREACAR 169.218 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 5.434 0 5.51 0.114 ;
    END
  END TxBypassDataExt
  PIN RxDfe1ClkC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.692208 LAYER M5 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 20.33 0 20.406 0.114 ;
    END
  END RxDfe1ClkC
  PIN RxDfe1ClkT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.680048 LAYER M5 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 22.61 0 22.686 0.114 ;
    END
  END RxDfe1ClkT
  PIN RxDfe0ClkT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.692208 LAYER M5 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 19.114 0 19.19 0.114 ;
    END
  END RxDfe0ClkT
  PIN RxDfe1DataClkT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.670092 LAYER M5 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 27.778 0 27.854 0.114 ;
    END
  END RxDfe1DataClkT
  PIN RxDfe0DataClkT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.670092 LAYER M5 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 13.186 0 13.262 0.114 ;
    END
  END RxDfe0DataClkT
  PIN OdtEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.106628 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 584.311 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 4.826 0 4.902 0.114 ;
    END
  END OdtEn
  PIN RxBypassData[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.692208 LAYER M5 ;
    ANTENNADIFFAREA 0.0037239375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 27.474 0 27.55 0.114 ;
    END
  END RxBypassData[2]
  PIN RxBypassData[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.692208 LAYER M5 ;
    ANTENNADIFFAREA 0.0037239375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 28.082 0 28.158 0.114 ;
    END
  END RxBypassData[3]
  PIN RxBypassRcvEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.692208 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002432 LAYER M5 ;
      ANTENNAMAXAREACAR 748.255 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 20.482 0 20.558 0.114 ;
    END
  END RxBypassRcvEn
  PIN TxBypassModeInt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.095228 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 448.218 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 3.61 0 3.686 0.114 ;
    END
  END TxBypassModeInt
  PIN IOPAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1502 LAYER M6 ;
    ANTENNADIFFAREA 0 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 11.0233 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 18.823 18.22 40.74 18.82 ;
    END
    PORT
      LAYER M6 ;
        RECT 5.601 87.075 35.439 87.525 ;
        RECT 5.601 85.275 35.439 85.725 ;
        RECT 5.601 83.475 35.439 83.925 ;
        RECT 5.601 81.675 35.439 82.125 ;
        RECT 5.601 79.875 35.439 80.325 ;
        RECT 5.601 75.375 35.439 75.825 ;
        RECT 5.601 73.575 35.439 74.025 ;
        RECT 5.601 71.775 35.439 72.225 ;
        RECT 5.601 69.975 35.439 70.425 ;
        RECT 5.601 68.175 35.439 68.625 ;
    END
    PORT
      LAYER M6 ;
        RECT 22.7705 64.975 40.385 65.475 ;
        RECT 22.7705 55.825 40.385 56.325 ;
        RECT 0.655 55.825 18.2695 56.325 ;
        RECT 22.7705 46.815 40.385 47.315 ;
        RECT 0.655 46.815 18.2695 47.315 ;
        RECT 0.655 37.665 18.2695 38.165 ;
        RECT 0.655 64.975 18.2695 65.475 ;
        RECT 22.7705 37.665 40.385 38.165 ;
    END
  END IOPAD
  PIN TxBypassModeExt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.086868 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 199.05 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 3.762 0 3.838 0.114 ;
    END
  END TxBypassModeExt
  PIN TxBypassOEExt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.335578 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002176 LAYER M5 ;
      ANTENNAMAXAREACAR 195.969 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 6.65 0 6.726 0.114 ;
    END
  END TxBypassOEExt
  PIN TxBypassOEInt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.335844 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002176 LAYER M5 ;
      ANTENNAMAXAREACAR 198.575 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 6.042 0 6.118 0.114 ;
    END
  END TxBypassOEInt
  PIN ZQCalCodePD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0970519375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 416.287 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 38.57 0 38.646 0.114 ;
    END
  END ZQCalCodePD[1]
  PIN ZQCalCodePD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1244119375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 456.003 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 38.722 0 38.798 0.114 ;
    END
  END ZQCalCodePD[2]
  PIN ZQCalCodePD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133532 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 476.044 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 38.874 0 38.95 0.114 ;
    END
  END ZQCalCodePD[3]
  PIN ZQCalCodePD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.160892 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 516.246 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 39.026 0 39.102 0.114 ;
    END
  END ZQCalCodePD[4]
  PIN ZQCalCodePD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.170012 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 536.044 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 39.178 0 39.254 0.114 ;
    END
  END ZQCalCodePD[5]
  PIN ZQCalCodePD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.197372 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 564.799 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 39.33 0 39.406 0.114 ;
    END
  END ZQCalCodePD[6]
  PIN ZQCalCodePD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.206492 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 596.105 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 39.482 0 39.558 0.114 ;
    END
  END ZQCalCodePD[7]
  PIN ZQCalCodePD[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.233852 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 624.482 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 39.634 0 39.71 0.114 ;
    END
  END ZQCalCodePD[8]
  PIN ZQCalCodePU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.278084 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1182.48 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.482 0 1.558 0.114 ;
    END
  END ZQCalCodePU[0]
  PIN ZQCalCodePU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.259844 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1197.79 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.634 0 1.71 0.114 ;
    END
  END ZQCalCodePU[1]
  PIN ZQCalCodePU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.223364 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1232.4 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.786 0 1.862 0.114 ;
    END
  END ZQCalCodePU[2]
  PIN ZQCalCodePU[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.132164 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 779.21 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.938 0 2.014 0.114 ;
    END
  END ZQCalCodePU[3]
  PIN ZQCalCodePU[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.159524 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 802.78 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 2.09 0 2.166 0.114 ;
    END
  END ZQCalCodePU[4]
  PIN ZQCalCodePU[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.323684 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1073.89 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 2.242 0 2.318 0.114 ;
    END
  END ZQCalCodePU[5]
  PIN ZQCalCodePU[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2963239375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1155.57 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 2.394 0 2.47 0.114 ;
    END
  END ZQCalCodePU[6]
  PIN ZQCalCodePU[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.186884 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 925.747 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 2.546 0 2.622 0.114 ;
    END
  END ZQCalCodePU[7]
  PIN ZQCalCodePU[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1686439375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1029.45 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 2.698 0 2.774 0.114 ;
    END
  END ZQCalCodePU[8]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.3 22.27 40.74 22.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 18.22 18.196 18.82 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 16.27 40.74 16.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 14.27 40.74 14.77 ;
        RECT 0.3 10.27 40.74 10.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 12.27 40.74 12.77 ;
        RECT 0.3 8.27 40.74 8.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 64.075 40.74 64.525 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 6.27 40.74 6.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 2.27 40.74 2.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 0.27 40.74 0.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 61.375 40.74 61.825 ;
        RECT 0.3 51.765 40.74 52.215 ;
        RECT 0.3 41.315 40.74 41.765 ;
        RECT 0.3 38.615 40.74 39.065 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 26.27 40.74 26.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 24.27 40.74 24.77 ;
    END
  END VDD
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.3 88.875 40.74 89.325 ;
        RECT 0.3 78.075 40.74 78.525 ;
        RECT 0.3 76.275 40.74 76.725 ;
        RECT 0.3 74.475 40.74 74.925 ;
        RECT 0.3 72.675 40.74 73.125 ;
        RECT 0.3 70.875 40.74 71.325 ;
        RECT 0.3 69.075 40.74 69.525 ;
        RECT 0.3 67.273 40.74 67.723 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 59.348 40.74 59.798 ;
        RECT 0.3 57.548 40.74 57.998 ;
        RECT 0.3 54.525 40.74 54.975 ;
        RECT 0.3 52.725 40.74 53.175 ;
        RECT 0.3 49.965 40.74 50.415 ;
        RECT 0.3 48.165 40.74 48.615 ;
        RECT 0.3 43.342 40.74 43.792 ;
        RECT 0.3 40.415 40.74 40.865 ;
        RECT 0.3 62.275 40.74 62.725 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 36.27 40.74 36.77 ;
        RECT 0.3 45.142 40.74 45.592 ;
    END
  END VDDQ
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M6 ;
        RECT 0.3 21.27 40.74 21.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 17.27 40.74 17.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 15.27 40.74 15.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 13.27 40.74 13.77 ;
        RECT 0.3 9.27 40.74 9.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 87.975 40.74 88.425 ;
        RECT 0.3 86.175 40.74 86.625 ;
        RECT 0.3 84.375 40.74 84.825 ;
        RECT 0.3 82.575 40.74 83.025 ;
        RECT 0.3 80.775 40.74 81.225 ;
        RECT 0.3 78.975 40.74 79.425 ;
        RECT 0.3 77.175 40.74 77.625 ;
        RECT 0.3 66.373 40.74 66.823 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 63.175 40.74 63.625 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 11.27 40.74 11.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 7.27 40.74 7.77 ;
        RECT 0.3 5.27 40.74 5.77 ;
        RECT 0.3 3.27 40.74 3.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 1.27 40.74 1.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 60.475 40.74 60.925 ;
        RECT 0.3 58.448 40.74 58.898 ;
        RECT 0.3 53.625 40.74 54.075 ;
        RECT 0.3 50.865 40.74 51.315 ;
        RECT 0.3 49.065 40.74 49.515 ;
        RECT 0.3 44.242 40.74 44.692 ;
        RECT 0.3 42.215 40.74 42.665 ;
        RECT 0.3 39.515 40.74 39.965 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 33.77 40.74 34.27 ;
        RECT 0.3 28.77 40.74 29.27 ;
        RECT 0.3 35.27 40.74 35.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 27.27 40.74 27.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 25.27 40.74 25.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 23.27 40.74 23.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 19.27 40.74 19.77 ;
    END
  END VSS
  PIN CoreLoopBackMode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.647748 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001696 LAYER M5 ;
      ANTENNAMAXAREACAR 1132.27 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 21.85 0 21.926 0.114 ;
    END
  END CoreLoopBackMode
  PIN RxDfe0ClkC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.642048 LAYER M5 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 18.354 0 18.43 0.114 ;
    END
  END RxDfe0ClkC
  PIN RxDfe1DataClkC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.670092 LAYER M5 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 27.17 0 27.246 0.114 ;
    END
  END RxDfe1DataClkC
  PIN RxDfe0DataClkC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.670092 LAYER M5 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 13.794 0 13.87 0.114 ;
    END
  END RxDfe0DataClkC
  PIN RxBypassDataPad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.667888 LAYER M5 ;
    ANTENNADIFFAREA 0.0148959375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 22.458 0 22.534 0.114 ;
    END
  END RxBypassDataPad
  PIN RxClkC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.74916 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.024736 LAYER M5 ;
      ANTENNAMAXAREACAR 1259.98 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 20.919 0 21.033 0.114 ;
    END
  END RxClkC
  PIN RxClkT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6723599375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.024736 LAYER M5 ;
      ANTENNAMAXAREACAR 1250.43 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 19.703 0 19.817 0.114 ;
    END
  END RxClkT
  PIN RxStandby
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.667888 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1444.77 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 18.81 0 18.886 0.114 ;
    END
  END RxStandby
  PIN RxPowerDown
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.657932 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1246.09 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 18.658 0 18.734 0.114 ;
    END
  END RxPowerDown
  PIN RxBypassData[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.680048 LAYER M5 ;
    ANTENNADIFFAREA 0.0037239375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 13.49 0 13.566 0.114 ;
    END
  END RxBypassData[0]
  PIN RxBypassPadEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7043679375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.016432 LAYER M5 ;
      ANTENNAMAXAREACAR 60.15 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 22.306 0 22.382 0.114 ;
    END
  END RxBypassPadEn
  PIN RxVrefCtl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.705394 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 1760.16 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 20.634 0 20.71 0.114 ;
    END
  END RxVrefCtl[0]
  PIN RxVrefCtl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.692208 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 20.026 0 20.102 0.114 ;
    END
  END RxVrefCtl[1]
  PIN TxSlewPU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0857659375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 15.618 0 15.694 0.114 ;
    END
  END TxSlewPU[0]
  PIN RxVrefDAC0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.369284 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 925.893 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 5.13 0 5.206 0.114 ;
    END
  END RxVrefDAC0[0]
  PIN RxVrefDAC0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.351044 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 910.557 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 4.522 0 4.598 0.114 ;
    END
  END RxVrefDAC0[1]
  PIN RxVrefDAC0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.332804 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 900.646 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 4.218 0 4.294 0.114 ;
    END
  END RxVrefDAC0[2]
  PIN RxVrefDAC0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.305444 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 883.986 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 3.914 0 3.99 0.114 ;
    END
  END RxVrefDAC0[3]
  PIN RxVrefDAC0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.241604 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 827.085 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 3.002 0 3.078 0.114 ;
    END
  END RxVrefDAC0[4]
  PIN RxVrefDAC0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.341924 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 795.033 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.33 0 1.406 0.114 ;
    END
  END RxVrefDAC0[5]
  PIN RxVrefDAC0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.396644 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 820.984 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.178 0 1.254 0.114 ;
    END
  END RxVrefDAC0[6]
  PIN RxVrefDAC1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.405764 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 882.638 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 0.114 0 0.19 0.114 ;
    END
  END RxVrefDAC1[0]
  PIN RxVrefDAC1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.396644 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 874.408 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 0.266 0 0.342 0.114 ;
    END
  END RxVrefDAC1[1]
  PIN RxVrefDAC1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.387524 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 859.159 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 0.418 0 0.494 0.114 ;
    END
  END RxVrefDAC1[2]
  PIN RxVrefDAC1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.378404 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 849.697 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 0.57 0 0.646 0.114 ;
    END
  END RxVrefDAC1[3]
  PIN RxVrefDAC1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.369284 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 835.461 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 0.722 0 0.798 0.114 ;
    END
  END RxVrefDAC1[4]
  PIN RxVrefDAC1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.360164 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 829.984 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 0.874 0 0.95 0.114 ;
    END
  END RxVrefDAC1[5]
  PIN RxVrefDAC1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.405764 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 843.24 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.026 0 1.102 0.114 ;
    END
  END RxVrefDAC1[6]
  PIN RxVrefDAC2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.424004 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 887.312 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 37.05 0 37.126 0.114 ;
    END
  END RxVrefDAC2[0]
  PIN RxVrefDAC2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4148839375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 891.607 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 37.354 0 37.43 0.114 ;
    END
  END RxVrefDAC2[1]
  PIN RxVrefDAC2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.387524 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 870.428 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 37.81 0 37.886 0.114 ;
    END
  END RxVrefDAC2[2]
  PIN RxVrefDAC2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.396644 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 874.588 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 37.962 0 38.038 0.114 ;
    END
  END RxVrefDAC2[3]
  PIN RxVrefDAC2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.031882 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 664.569 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 38.114 0 38.19 0.114 ;
    END
  END RxVrefDAC2[4]
  PIN RxVrefDAC2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.060192 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 758.171 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 38.266 0 38.342 0.114 ;
    END
  END RxVrefDAC2[5]
  PIN RxVrefDAC2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.072314 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 695.26 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 39.786 0 39.862 0.114 ;
    END
  END RxVrefDAC2[6]
  PIN RxVrefDAC3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.405764 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 885.253 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 40.85 0 40.926 0.114 ;
    END
  END RxVrefDAC3[0]
  PIN RxVrefDAC3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.396644 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 873.574 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 40.698 0 40.774 0.114 ;
    END
  END RxVrefDAC3[1]
  PIN RxVrefDAC3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.387524 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 859.751 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 40.546 0 40.622 0.114 ;
    END
  END RxVrefDAC3[2]
  PIN RxVrefDAC3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.378404 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 850.225 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 40.394 0 40.47 0.114 ;
    END
  END RxVrefDAC3[3]
  PIN RxVrefDAC3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.332804 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 820.793 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 40.242 0 40.318 0.114 ;
    END
  END RxVrefDAC3[4]
  PIN RxVrefDAC3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.351044 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 827.496 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 40.09 0 40.166 0.114 ;
    END
  END RxVrefDAC3[5]
  PIN RxVrefDAC3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.405764 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 846.751 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 39.938 0 40.014 0.114 ;
    END
  END RxVrefDAC3[6]
  PIN VrefDacRef
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.3415 LAYER M6 ;
    ANTENNADIFFAREA 4.4494 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 0 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 6.057 31.27 40.74 31.77 ;
    END
  END VrefDacRef
  PIN OdtStrenCodePD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.099294 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 96.8758 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 35.226 0 35.302 0.114 ;
    END
  END OdtStrenCodePD[0]
  PIN OdtStrenCodePD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.142006 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 119.631 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 29.146 0 29.222 0.114 ;
    END
  END OdtStrenCodePD[1]
  PIN OdtStrenCodePD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19038 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 135.937 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 35.53 0 35.606 0.114 ;
    END
  END OdtStrenCodePD[2]
  PIN OdtStrenCodePD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.184034 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 136.817 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 29.45 0 29.526 0.114 ;
    END
  END OdtStrenCodePD[3]
  PIN OdtStrenCodePU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.142234 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 132.96 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 22.002 0 22.078 0.114 ;
    END
  END OdtStrenCodePU[0]
  PIN OdtStrenCodePU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.109212 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 122.748 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 17.29 0 17.366 0.114 ;
    END
  END OdtStrenCodePU[1]
  PIN OdtStrenCodePU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2204 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 155.707 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 23.674 0 23.75 0.114 ;
    END
  END OdtStrenCodePU[2]
  PIN OdtStrenCodePU[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.14288 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 138.602 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 16.378 0 16.454 0.114 ;
    END
  END OdtStrenCodePU[3]
  PIN OdtStrenCodePU[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.092112 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 23.826 0 23.902 0.114 ;
    END
  END OdtStrenCodePU[4]
  PIN OdtStrenCodePU[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.109212 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 16.226 0 16.302 0.114 ;
    END
  END OdtStrenCodePU[5]
  PIN OdtStrenCodePU[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.092112 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 23.978 0 24.054 0.114 ;
    END
  END OdtStrenCodePU[6]
  PIN OdtStrenCodePU[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.109212 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 16.074 0 16.15 0.114 ;
    END
  END OdtStrenCodePU[7]
  PIN VDD_TIEHI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 0.3 31.27 5.457 31.77 ;
    END
  END VDD_TIEHI
  PIN RxBypassData[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.680048 LAYER M5 ;
    ANTENNADIFFAREA 0.0037239375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 12.882 0 12.958 0.114 ;
    END
  END RxBypassData[1]
  PIN TxClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.159087 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 339.034 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 6.403 0 6.517 0.114 ;
    END
  END TxClk
  PIN TxData
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.118522 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002432 LAYER M5 ;
      ANTENNAMAXAREACAR 88.586299938 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 7.41 0 7.486 0.114 ;
    END
  END TxData
  PIN TxModeCtl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.256158 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 6.802 0 6.878 0.114 ;
    END
  END TxModeCtl[1]
  PIN TxModeCtl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.124868 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 7.106 0 7.182 0.114 ;
    END
  END TxModeCtl[2]
  PIN TxOE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.161728 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.004864 LAYER M5 ;
      ANTENNAMAXAREACAR 87.1377 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 7.714 0 7.79 0.114 ;
    END
  END TxOE
  PIN TxStrenCodePD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.124716 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003808 LAYER M5 ;
      ANTENNAMAXAREACAR 107.973 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 34.922 0 34.998 0.114 ;
    END
  END TxStrenCodePD[0]
  PIN TxStrenCodePD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1429179375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003808 LAYER M5 ;
      ANTENNAMAXAREACAR 109.907 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 28.842 0 28.918 0.114 ;
    END
  END TxStrenCodePD[1]
  PIN TxStrenCodePD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.182704 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003808 LAYER M5 ;
      ANTENNAMAXAREACAR 118.474 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 34.618 0 34.694 0.114 ;
    END
  END TxStrenCodePD[2]
  PIN TxStrenCodePD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.180614 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003808 LAYER M5 ;
      ANTENNAMAXAREACAR 115.73 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 28.538 0 28.614 0.114 ;
    END
  END TxStrenCodePD[3]
  PIN TxStrenCodePU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1427279375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003264 LAYER M5 ;
      ANTENNAMAXAREACAR 130.893 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 23.37 0 23.446 0.114 ;
    END
  END TxStrenCodePU[0]
  OBS
    LAYER M1 ;
      RECT MASK 1 0 0 41.04 90 ;
      RECT MASK 2 0 0 41.04 90 ;
    LAYER M2 ;
      RECT MASK 1 0 0 41.04 90 ;
      RECT MASK 2 0 0 41.04 90 ;
    LAYER M3 ;
      RECT MASK 1 0 0 41.04 90 ;
      RECT MASK 2 0 0 41.04 90 ;
    LAYER M4 ;
      POLYGON 41.04 0 41.04 90 0 90 0 47.941 21.08 47.941 21.08 47.315 0 47.315 0 0 ;
      RECT 9.8465 0.8 38.2005 0.86 ;
      RECT 4.2125 0.92 34.3475 0.98 ;
      RECT 35.161 1.04 35.531 1.1 ;
      RECT 38.374 1.058 40.0995 1.118 ;
      RECT 1.415 1.16 4.23 1.22 ;
      RECT 4.5255 1.16 7.055 1.22 ;
      RECT 7.299 1.16 7.9715 1.22 ;
      RECT 8.9465 1.16 10.871 1.22 ;
      RECT 17.742 1.16 21.712 1.22 ;
      RECT 8.595 1.171 8.733 1.209 ;
      RECT 38.374 1.178 40.0995 1.238 ;
      RECT 4.5945 1.28 4.9645 1.34 ;
      RECT 5.1715 1.28 5.564 1.34 ;
      RECT 6.0625 1.28 6.56 1.34 ;
      RECT 9.684 1.28 38.0385 1.34 ;
      RECT 38.374 1.298 40.0995 1.358 ;
      RECT 38.374 1.418 40.0995 1.478 ;
      RECT 38.374 1.538 40.0995 1.598 ;
      RECT 1.891 1.64 3.621 1.7 ;
      RECT 3.7345 1.64 6.0565 1.7 ;
      RECT 7.793 1.64 8.912 1.7 ;
      RECT 9.014 1.64 10.872 1.7 ;
      RECT 16.0785 1.64 16.485 1.7 ;
      RECT 16.609 1.64 17.081 1.7 ;
      RECT 17.2635 1.64 17.6335 1.7 ;
      RECT 21.965 1.64 22.724 1.7 ;
      RECT 28.537 1.64 28.949 1.7 ;
      RECT 29.066 1.64 29.464 1.7 ;
      RECT 38.374 1.658 40.0995 1.718 ;
      RECT 2.055 1.76 3.6835 1.82 ;
      RECT 4.077 1.76 33.757 1.82 ;
      RECT 38.374 1.778 40.0995 1.838 ;
      RECT 2.643 1.88 3.7405 1.94 ;
      RECT 5.8975 1.88 7.705 1.94 ;
      RECT 7.813 1.88 9.6745 1.94 ;
      RECT 9.8465 1.88 38.186 1.94 ;
      RECT 38.374 1.898 40.0995 1.958 ;
      RECT 2.051 2 4.4465 2.06 ;
      RECT 4.7555 2 6.052 2.06 ;
      RECT 6.255 2 7.831 2.06 ;
      RECT 8.049 2 9.556 2.06 ;
      RECT 38.374 2.018 40.0995 2.078 ;
      RECT 2.667 2.12 9.3 2.18 ;
      RECT 38.374 2.138 40.0995 2.198 ;
      RECT 2.375 2.24 8.498 2.3 ;
      RECT 8.963 2.24 10.872 2.3 ;
      RECT 11.961 2.24 21.116 2.3 ;
      RECT 22.9945 2.24 23.4115 2.3 ;
      RECT 30.013 2.24 33.983 2.3 ;
      RECT 38.374 2.258 40.125 2.318 ;
      RECT 2.515 2.36 8.0045 2.42 ;
      RECT 8.12 2.36 9.556 2.42 ;
      RECT 10.3355 2.36 33.396 2.42 ;
      RECT 38.374 2.378 40.0995 2.438 ;
      RECT 2.895 2.48 7.588 2.54 ;
      RECT 9.811 2.48 38.033 2.54 ;
      RECT 38.374 2.498 40.0995 2.558 ;
      RECT 3.118 2.6 9.556 2.66 ;
      RECT 9.811 2.6 38.033 2.66 ;
      RECT 38.374 2.618 40.0995 2.678 ;
      RECT 2.215 2.72 6.3895 2.78 ;
      RECT 6.488 2.72 6.909 2.78 ;
      RECT 7.081 2.72 10.405 2.78 ;
      RECT 10.922 2.72 21.075 2.78 ;
      RECT 22.3415 2.72 23.8545 2.78 ;
      RECT 24.295 2.72 28.265 2.78 ;
      RECT 38.374 2.738 40.0995 2.798 ;
      RECT 1.731 2.84 9.44 2.9 ;
      RECT 9.659 2.84 38.1895 2.9 ;
      RECT 38.374 2.858 40.0995 2.918 ;
      RECT 1.895 2.96 8.222 3.02 ;
      RECT 8.398 2.96 10.872 3.02 ;
      RECT 38.374 2.978 40.0995 3.038 ;
      RECT 3.311 3.08 38.1895 3.14 ;
      RECT 3.332 3.2 38.191 3.26 ;
      RECT 38.374 3.2 40.0995 3.26 ;
      RECT 3.1195 3.32 39.9065 3.38 ;
      RECT 1.735 3.44 7.833 3.5 ;
      RECT 11.978 3.44 22.278 3.5 ;
      RECT 23.459 3.44 33.759 3.5 ;
      RECT 34.516 3.44 39.465 3.5 ;
      RECT 1.394 3.56 7.671 3.62 ;
      RECT 9.811 3.56 39.9065 3.62 ;
      RECT 1.575 3.68 6.5225 3.74 ;
      RECT 11.978 3.68 22.278 3.74 ;
      RECT 23.459 3.68 33.759 3.74 ;
      RECT 34.516 3.68 39.465 3.74 ;
      RECT 2.306 3.8 7.363 3.86 ;
      RECT 9.811 3.8 39.9065 3.86 ;
      RECT 4.911 3.92 9.247 3.98 ;
      RECT 9.811 3.92 39.9065 3.98 ;
      RECT 2.7175 4.04 7.8545 4.1 ;
      RECT 9.6715 4.04 19.541 4.1 ;
      RECT 20.9215 4.04 38.8555 4.1 ;
      RECT 2.154 4.16 3.165 4.22 ;
      RECT 4.911 4.16 9.247 4.22 ;
      RECT 38.984 4.16 40.128 4.22 ;
      RECT 8.231 4.28 39.465 4.34 ;
      RECT 3.1525 4.4 39.465 4.46 ;
      RECT 9.0895 4.52 39.396 4.58 ;
      RECT 3.105 4.64 4.619 4.7 ;
      RECT 4.911 4.64 9.247 4.7 ;
      RECT 11.978 4.64 22.278 4.7 ;
      RECT 39.132 4.64 39.965 4.7 ;
      RECT 11.6015 4.76 22.3815 4.82 ;
      RECT 38.534 5.24 39.815 5.3 ;
      RECT 19.691 10.148 19.829 10.228 ;
      RECT 22.109 10.148 22.179 10.228 ;
      RECT 18.7195 11.068 22.3195 11.493 ;
      RECT 18.752 13.438 22.288 13.863 ;
      RECT 18.7195 15.778 22.3195 16.203 ;
      RECT 14.192 16.569 26.848 16.96 ;
      RECT 18.72 19.051 22.32 19.437 ;
      RECT 13.362 37.888 16.498 38.313 ;
      RECT 16.698 37.888 20.234 38.313 ;
      RECT 20.806 37.888 24.342 38.313 ;
      RECT 24.542 37.888 27.678 38.313 ;
      RECT 0.655 37.907 13.155 37.945 ;
      RECT 27.885 37.907 40.385 37.945 ;
      RECT 0.655 38.059 13.155 38.097 ;
      RECT 27.885 38.059 40.385 38.097 ;
      RECT 0.655 38.211 13.155 38.249 ;
      RECT 27.885 38.211 40.385 38.249 ;
      RECT 0.655 38.363 13.155 38.401 ;
      RECT 27.885 38.363 40.385 38.401 ;
      RECT 0.655 38.515 13.155 38.553 ;
      RECT 27.885 38.515 40.385 38.553 ;
      RECT 13.674 38.5495 19.694 38.9405 ;
      RECT 21.346 38.5495 27.366 38.9405 ;
      RECT 0.655 38.667 13.155 38.705 ;
      RECT 27.885 38.667 40.385 38.705 ;
      RECT 0.655 38.819 13.155 38.857 ;
      RECT 27.885 38.819 40.385 38.857 ;
      RECT 0.655 38.971 13.155 39.009 ;
      RECT 27.885 38.971 40.385 39.009 ;
      RECT 0.655 39.123 13.155 39.161 ;
      RECT 27.885 39.123 40.385 39.161 ;
      RECT 0.655 39.275 13.155 39.313 ;
      RECT 27.885 39.275 40.385 39.313 ;
      RECT 0.655 39.427 13.155 39.465 ;
      RECT 27.885 39.427 40.385 39.465 ;
      RECT 0.655 39.579 13.155 39.617 ;
      RECT 27.885 39.579 40.385 39.617 ;
      RECT 0.655 39.731 13.155 39.769 ;
      RECT 27.885 39.731 40.385 39.769 ;
      RECT 0.655 40.076 20.2375 40.256 ;
      RECT 20.8025 40.076 40.385 40.256 ;
      RECT 0.732 41.125 4.2835 41.185 ;
      RECT 4.609 41.125 19.995 41.185 ;
      RECT 21.045 41.125 36.431 41.185 ;
      RECT 36.7565 41.125 40.308 41.185 ;
      RECT 0.7575 41.365 40.2825 41.425 ;
      RECT 0.729 41.485 4.2835 41.545 ;
      RECT 4.609 41.485 19.995 41.545 ;
      RECT 21.045 41.485 36.431 41.545 ;
      RECT 36.7565 41.485 40.311 41.545 ;
      RECT 0.729 41.725 20.015 41.785 ;
      RECT 21.025 41.725 40.311 41.785 ;
      RECT 4.03 41.845 16.937 41.905 ;
      RECT 24.103 41.845 37.01 41.905 ;
      RECT 0.369 41.965 21.1695 42.025 ;
      RECT 0.7185 42.085 20.015 42.145 ;
      RECT 21.025 42.085 40.3215 42.145 ;
      RECT 0.068 42.205 21.1695 42.265 ;
      RECT 0.7185 42.325 20.015 42.385 ;
      RECT 21.025 42.325 40.3215 42.385 ;
      RECT 1.1635 42.445 21.1695 42.505 ;
      RECT 0.2275 42.565 40.2825 42.625 ;
      RECT 6.2355 43.425 17.7635 43.485 ;
      RECT 23.2765 43.425 34.8045 43.485 ;
      RECT 0.734 45.105 18.5435 45.165 ;
      RECT 22.4965 45.105 40.306 45.165 ;
      RECT 0.734 45.345 18.5515 45.405 ;
      RECT 22.4885 45.345 40.306 45.405 ;
      RECT 1.739 46.199 17.185 46.499 ;
      RECT 23.855 46.199 39.301 46.499 ;
      RECT 1.2285 46.915 17.842 47.215 ;
      RECT 23.198 46.915 39.8115 47.215 ;
      RECT 1.071 49.14 17.849 49.2 ;
      RECT 23.191 49.14 39.969 49.2 ;
      RECT 1.64 49.26 17.284 49.32 ;
      RECT 23.756 49.26 39.4 49.32 ;
      RECT 1.071 49.38 17.849 49.44 ;
      RECT 23.191 49.38 39.969 49.44 ;
      RECT 1.0745 52.483 9.1855 52.597 ;
      RECT 32.076 52.483 40.0075 52.597 ;
      RECT 1.071 53.7 17.849 53.76 ;
      RECT 23.191 53.7 39.969 53.76 ;
      RECT 1.64 53.82 17.284 53.88 ;
      RECT 23.756 53.82 39.4 53.88 ;
      RECT 1.071 53.94 17.849 54 ;
      RECT 23.191 53.94 39.969 54 ;
      RECT 1.2285 55.925 17.842 56.225 ;
      RECT 23.198 55.925 39.8115 56.225 ;
      RECT 1.739 56.641 17.185 56.941 ;
      RECT 23.855 56.641 39.301 56.941 ;
      RECT 0.734 57.735 18.5515 57.795 ;
      RECT 22.4885 57.735 40.306 57.795 ;
      RECT 0.734 57.975 18.5435 58.035 ;
      RECT 22.4965 57.975 40.306 58.035 ;
      RECT 6.2355 59.655 17.7635 59.715 ;
      RECT 23.2765 59.655 34.8045 59.715 ;
      RECT 0.2275 60.515 40.2825 60.575 ;
      RECT 1.1635 60.635 21.1695 60.695 ;
      RECT 0.7185 60.755 40.3215 60.815 ;
      RECT 0.068 60.875 21.1695 60.935 ;
      RECT 0.7185 60.995 40.3215 61.055 ;
      RECT 0.369 61.115 21.1695 61.175 ;
      RECT 4.03 61.235 16.937 61.295 ;
      RECT 24.103 61.235 37.01 61.295 ;
      RECT 0.729 61.355 20.015 61.415 ;
      RECT 21.025 61.355 40.311 61.415 ;
      RECT 0.729 61.595 4.2835 61.655 ;
      RECT 4.609 61.595 36.431 61.655 ;
      RECT 36.7565 61.595 40.311 61.655 ;
      RECT 0.7575 61.715 40.2825 61.775 ;
      RECT 0.732 61.955 4.2835 62.015 ;
      RECT 4.609 61.955 19.995 62.015 ;
      RECT 21.045 61.955 36.431 62.015 ;
      RECT 36.7565 61.955 40.308 62.015 ;
      RECT 0.655 62.884 20.2375 63.064 ;
      RECT 20.8025 62.884 40.385 63.064 ;
      RECT 0.655 63.371 13.155 63.409 ;
      RECT 27.885 63.371 40.385 63.409 ;
      RECT 0.655 63.523 13.155 63.561 ;
      RECT 27.885 63.523 40.385 63.561 ;
      RECT 0.655 63.675 13.155 63.713 ;
      RECT 27.885 63.675 40.385 63.713 ;
      RECT 0.655 63.827 13.155 63.865 ;
      RECT 27.885 63.827 40.385 63.865 ;
      RECT 0.655 63.979 13.155 64.017 ;
      RECT 27.885 63.979 40.385 64.017 ;
      RECT 0.655 64.131 13.155 64.169 ;
      RECT 27.885 64.131 40.385 64.169 ;
      RECT 13.674 64.1995 19.694 64.5905 ;
      RECT 21.346 64.1995 27.366 64.5905 ;
      RECT 0.655 64.283 13.155 64.321 ;
      RECT 27.885 64.283 40.385 64.321 ;
      RECT 0.655 64.435 13.155 64.473 ;
      RECT 27.885 64.435 40.385 64.473 ;
      RECT 0.655 64.587 13.155 64.625 ;
      RECT 27.885 64.587 40.385 64.625 ;
      RECT 0.655 64.739 13.155 64.777 ;
      RECT 27.885 64.739 40.385 64.777 ;
      RECT 13.362 64.827 16.498 65.252 ;
      RECT 16.698 64.827 20.234 65.252 ;
      RECT 20.806 64.827 24.342 65.252 ;
      RECT 24.542 64.827 27.678 65.252 ;
      RECT 0.655 64.891 13.155 64.929 ;
      RECT 27.885 64.891 40.385 64.929 ;
      RECT 0.655 65.043 13.155 65.081 ;
      RECT 27.885 65.043 40.385 65.081 ;
      RECT 0.655 65.195 13.155 65.233 ;
      RECT 27.885 65.195 40.385 65.233 ;
      RECT 0.3 66.43 40.74 66.79 ;
      RECT 5.6 68.15 35.44 68.65 ;
      RECT 0.3 69.05 40.74 69.55 ;
      RECT 5.6 69.95 35.44 70.45 ;
      RECT 0.3 70.85 40.74 71.35 ;
      RECT 5.6 71.75 35.44 72.25 ;
      RECT 0.3 72.65 40.74 73.15 ;
      RECT 5.6 73.55 35.44 74.05 ;
      RECT 0.3 74.45 40.74 74.95 ;
      RECT 5.6 75.35 35.44 75.85 ;
      RECT 0.3 76.25 40.74 76.75 ;
      RECT 0.3 77.21 40.74 77.57 ;
      RECT 0.3 78.13 40.74 78.49 ;
      RECT 0.3 78.95 40.74 79.45 ;
      RECT 5.601 79.85 35.439 80.35 ;
      RECT 0.3 80.75 40.74 81.25 ;
      RECT 5.601 81.65 35.439 82.15 ;
      RECT 0.3 82.55 40.74 83.05 ;
      RECT 5.601 83.45 35.439 83.95 ;
      RECT 0.3 84.35 40.74 84.85 ;
      RECT 5.601 85.25 35.439 85.75 ;
      RECT 0.3 86.15 40.74 86.65 ;
      RECT 5.601 87.05 35.439 87.55 ;
      RECT 4.141 88.91 36.899 89.27 ;
      RECT 6.946 0.8 9.629 0.86 ;
      RECT 2.999 1.04 34.3475 1.1 ;
      RECT 6.8525 1.28 9.389 1.34 ;
      RECT 3.0045 1.52 35.7995 1.58 ;
      RECT 6.1755 1.64 7.2475 1.7 ;
      RECT 11.4525 1.64 15.4225 1.7 ;
      RECT 18.0925 1.64 21.6345 1.7 ;
      RECT 23.2615 1.64 23.6315 1.7 ;
      RECT 11.345 2 11.455 2.06 ;
      RECT 15.665 2 15.775 2.06 ;
      RECT 16.145 2 16.255 2.06 ;
      RECT 16.465 2 16.575 2.06 ;
      RECT 16.785 2 16.895 2.06 ;
      RECT 17.105 2 17.215 2.06 ;
      RECT 37.105 2 37.215 2.06 ;
      RECT 11.483 2.011 11.621 2.049 ;
      RECT 12.243 2.011 12.381 2.049 ;
      RECT 18.019 2.011 18.157 2.049 ;
      RECT 18.475 2.011 18.613 2.049 ;
      RECT 19.235 2.011 19.373 2.049 ;
      RECT 20.147 2.011 20.285 2.049 ;
      RECT 21.515 2.011 21.653 2.049 ;
      RECT 22.123 2.011 22.261 2.049 ;
      RECT 22.883 2.011 23.021 2.049 ;
      RECT 23.035 2.011 23.173 2.049 ;
      RECT 25.923 2.011 26.061 2.049 ;
      RECT 26.531 2.011 26.669 2.049 ;
      RECT 29.723 2.011 29.861 2.049 ;
      RECT 30.331 2.011 30.469 2.049 ;
      RECT 30.939 2.011 31.077 2.049 ;
      RECT 31.547 2.011 31.685 2.049 ;
      RECT 32.155 2.011 32.293 2.049 ;
      RECT 37.627 2.011 37.765 2.049 ;
      RECT 11.154 2.12 22.045 2.18 ;
      RECT 30.365 2.72 34.335 2.78 ;
      RECT 11.309 2.96 36.5895 3.02 ;
      RECT 11.978 4.16 22.278 4.22 ;
      RECT 23.459 4.16 33.759 4.22 ;
      RECT 23.459 4.64 33.759 4.7 ;
      RECT 18.909 10.468 18.979 10.548 ;
      RECT 20.907 10.468 21.045 10.548 ;
      RECT 18.7195 12.507 22.3195 12.932 ;
      RECT 18.752 14.877 22.288 15.302 ;
      RECT 18.7195 17.217 22.3195 17.642 ;
      RECT 0.655 37.496 13.155 37.676 ;
      RECT 27.885 37.496 40.385 37.676 ;
      RECT 0.655 37.983 13.155 38.021 ;
      RECT 27.885 37.983 40.385 38.021 ;
      RECT 0.655 38.135 13.155 38.173 ;
      RECT 27.885 38.135 40.385 38.173 ;
      RECT 0.655 38.287 13.155 38.325 ;
      RECT 27.885 38.287 40.385 38.325 ;
      RECT 0.655 38.439 13.155 38.477 ;
      RECT 27.885 38.439 40.385 38.477 ;
      RECT 0.655 38.591 13.155 38.629 ;
      RECT 27.885 38.591 40.385 38.629 ;
      RECT 0.655 38.743 13.155 38.781 ;
      RECT 27.885 38.743 40.385 38.781 ;
      RECT 0.655 38.895 13.155 38.933 ;
      RECT 27.885 38.895 40.385 38.933 ;
      RECT 0.655 39.047 13.155 39.085 ;
      RECT 27.885 39.047 40.385 39.085 ;
      RECT 13.362 39.177 16.498 39.602 ;
      RECT 16.698 39.177 20.234 39.602 ;
      RECT 20.806 39.177 24.342 39.602 ;
      RECT 24.542 39.177 27.678 39.602 ;
      RECT 0.655 39.199 13.155 39.237 ;
      RECT 27.885 39.199 40.385 39.237 ;
      RECT 0.655 39.351 13.155 39.389 ;
      RECT 27.885 39.351 40.385 39.389 ;
      RECT 0.655 39.503 13.155 39.541 ;
      RECT 27.885 39.503 40.385 39.541 ;
      RECT 0.655 39.655 13.155 39.693 ;
      RECT 27.885 39.655 40.385 39.693 ;
      RECT 0.655 39.807 13.155 39.845 ;
      RECT 27.885 39.807 40.385 39.845 ;
      RECT 0.7055 40.436 40.3345 40.55 ;
      RECT 0.7255 40.885 4.2835 40.945 ;
      RECT 4.609 40.885 19.995 40.945 ;
      RECT 21.045 40.885 36.431 40.945 ;
      RECT 36.7565 40.885 40.3145 40.945 ;
      RECT 0.882 43.545 18.4015 43.605 ;
      RECT 22.6385 43.545 40.158 43.605 ;
      RECT 0.882 43.785 18.4015 43.845 ;
      RECT 22.6385 43.785 40.158 43.845 ;
      RECT 0.815 48.653 18.0595 48.767 ;
      RECT 22.9805 48.653 40.225 48.767 ;
      RECT 1.07 48.906 17.8315 49.02 ;
      RECT 23.2085 48.906 39.97 49.02 ;
      RECT 1.07 49.713 17.8315 49.827 ;
      RECT 23.2085 49.713 39.97 49.827 ;
      RECT 0.815 49.97 18.0595 50.09 ;
      RECT 22.9805 49.97 40.225 50.09 ;
      RECT 0.815 53.05 18.0595 53.17 ;
      RECT 22.9805 53.05 40.225 53.17 ;
      RECT 1.07 53.313 17.8315 53.427 ;
      RECT 23.2085 53.313 39.97 53.427 ;
      RECT 1.07 54.12 17.8315 54.234 ;
      RECT 23.2085 54.12 39.97 54.234 ;
      RECT 0.815 54.373 18.0595 54.487 ;
      RECT 22.9805 54.373 40.225 54.487 ;
      RECT 0.882 59.295 18.4015 59.355 ;
      RECT 22.6385 59.295 40.158 59.355 ;
      RECT 0.882 59.535 18.4015 59.595 ;
      RECT 22.6385 59.535 40.158 59.595 ;
      RECT 0.7255 62.195 4.2835 62.255 ;
      RECT 4.609 62.195 19.995 62.255 ;
      RECT 21.045 62.195 36.431 62.255 ;
      RECT 36.7565 62.195 40.3145 62.255 ;
      RECT 0.7055 62.59 40.3345 62.704 ;
      RECT 0.655 63.295 13.155 63.333 ;
      RECT 27.885 63.295 40.385 63.333 ;
      RECT 0.655 63.447 13.155 63.485 ;
      RECT 27.885 63.447 40.385 63.485 ;
      RECT 13.362 63.538 16.498 63.963 ;
      RECT 16.698 63.538 20.234 63.963 ;
      RECT 20.806 63.538 24.342 63.963 ;
      RECT 24.542 63.538 27.678 63.963 ;
      RECT 0.655 63.599 13.155 63.637 ;
      RECT 27.885 63.599 40.385 63.637 ;
      RECT 0.655 63.751 13.155 63.789 ;
      RECT 27.885 63.751 40.385 63.789 ;
      RECT 0.655 63.903 13.155 63.941 ;
      RECT 27.885 63.903 40.385 63.941 ;
      RECT 0.655 64.055 13.155 64.093 ;
      RECT 27.885 64.055 40.385 64.093 ;
      RECT 0.655 64.207 13.155 64.245 ;
      RECT 27.885 64.207 40.385 64.245 ;
      RECT 0.655 64.359 13.155 64.397 ;
      RECT 27.885 64.359 40.385 64.397 ;
      RECT 0.655 64.511 13.155 64.549 ;
      RECT 27.885 64.511 40.385 64.549 ;
      RECT 0.655 64.663 13.155 64.701 ;
      RECT 27.885 64.663 40.385 64.701 ;
      RECT 0.655 64.815 13.155 64.853 ;
      RECT 27.885 64.815 40.385 64.853 ;
      RECT 0.655 64.967 13.155 65.005 ;
      RECT 27.885 64.967 40.385 65.005 ;
      RECT 0.655 65.119 13.155 65.157 ;
      RECT 27.885 65.119 40.385 65.157 ;
      RECT 0.655 65.464 13.155 65.644 ;
      RECT 27.885 65.464 40.385 65.644 ;
      RECT 4.907 67.25 36.133 67.75 ;
      RECT 4.907 69.05 36.133 69.55 ;
      RECT 4.907 70.85 36.133 71.35 ;
      RECT 4.907 72.65 36.133 73.15 ;
      RECT 4.907 74.45 36.133 74.95 ;
      RECT 4.907 76.25 36.133 76.75 ;
      RECT 4.907 78.95 36.133 79.45 ;
      RECT 4.907 80.75 36.133 81.25 ;
      RECT 4.907 82.55 36.133 83.05 ;
      RECT 4.907 84.35 36.133 84.85 ;
      RECT 4.907 86.15 36.133 86.65 ;
      RECT 4.907 87.95 36.133 88.45 ;
    LAYER M5 ;
      POLYGON 0 0 0 90 41.04 90 41.04 66.0715 20.22 66.0715 20.22 19.7315 20.82 19.7315 20.82 66.0715 41.04 66.0715 41.04 0 40.964 0 40.964 0.152 37.772 0.152 37.772 0 37.468 0 37.468 0.152 37.316 0.152 37.316 0 37.164 0 37.164 0.152 37.012 0.152 37.012 0 35.644 0 35.644 0.152 35.492 0.152 35.492 0 35.34 0 35.34 0.152 35.188 0.152 35.188 0 35.036 0 35.036 0.152 34.884 0.152 34.884 0 34.732 0 34.732 0.152 34.58 0.152 34.58 0 29.564 0 29.564 0.152 29.412 0.152 29.412 0 29.26 0 29.26 0.152 29.108 0.152 29.108 0 28.956 0 28.956 0.152 28.804 0.152 28.804 0 28.652 0 28.652 0.152 28.5 0.152 28.5 0 28.196 0 28.196 0.152 28.044 0.152 28.044 0 27.892 0 27.892 0.152 27.74 0.152 27.74 0 27.588 0 27.588 0.152 27.436 0.152 27.436 0 27.284 0 27.284 0.152 27.132 0.152 27.132 0 24.396 0 24.396 0.152 24.244 0.152 24.244 0 24.092 0 24.092 0.152 23.636 0.152 23.636 0 23.484 0 23.484 0.152 23.028 0.152 23.028 0 22.724 0 22.724 0.152 22.268 0.152 22.268 0 22.116 0 22.116 0.152 21.812 0.152 21.812 0 21.356 0 21.356 0.152 21.204 0.152 21.204 0 21.071 0 21.071 0.152 20.881 0.152 20.881 0 20.748 0 20.748 0.152 20.292 0.152 20.292 0 20.14 0 20.14 0.152 19.988 0.152 19.988 0 19.855 0 19.855 0.152 19.665 0.152 19.665 0 19.228 0 19.228 0.152 19.076 0.152 19.076 0 18.924 0 18.924 0.152 18.62 0.152 18.62 0 18.468 0 18.468 0.152 18.316 0.152 18.316 0 17.556 0 17.556 0.152 17.252 0.152 17.252 0 17.1 0 17.1 0.152 16.644 0.152 16.644 0 16.492 0 16.492 0.152 16.036 0.152 16.036 0 15.732 0 15.732 0.152 15.124 0.152 15.124 0 14.82 0 14.82 0.152 14.668 0.152 14.668 0 14.516 0 14.516 0.152 14.364 0.152 14.364 0 14.212 0 14.212 0.152 13.756 0.152 13.756 0 13.604 0 13.604 0.152 13.452 0.152 13.452 0 13.3 0 13.3 0.152 13.148 0.152 13.148 0 12.996 0 12.996 0.152 12.844 0.152 12.844 0 11.932 0 11.932 0.152 11.78 0.152 11.78 0 11.02 0 11.02 0.152 10.868 0.152 10.868 0 10.412 0 10.412 0.152 10.26 0.152 10.26 0 7.828 0 7.828 0.152 7.676 0.152 7.676 0 7.524 0 7.524 0.152 7.372 0.152 7.372 0 7.22 0 7.22 0.152 7.068 0.152 7.068 0 6.916 0 6.916 0.152 6.612 0.152 6.612 0 6.555 0 6.555 0.152 6.365 0.152 6.365 0 6.156 0 6.156 0.152 6.004 0.152 6.004 0 5.852 0 5.852 0.152 5.7 0.152 5.7 0 5.548 0 5.548 0.152 5.396 0.152 5.396 0 5.244 0 5.244 0.152 5.092 0.152 5.092 0 4.94 0 4.94 0.152 4.788 0.152 4.788 0 4.636 0 4.636 0.152 4.484 0.152 4.484 0 4.332 0 4.332 0.152 4.18 0.152 4.18 0 4.028 0 4.028 0.152 3.572 0.152 3.572 0 3.116 0 3.116 0.152 0.076 0.152 0.076 0 ;
      RECT 0.114 0.152 0.19 5.339 ;
      RECT 1.026 0.152 1.102 5.339 ;
      RECT 2.85 0.152 2.926 8.116 ;
      RECT 4.826 0.152 4.902 1.403 ;
      RECT 6.403 0.152 6.517 1.3955 ;
      RECT 7.106 0.152 7.182 1.643 ;
      RECT 7.714 0.152 7.79 2.128 ;
      RECT 10.298 0.152 10.374 2.865 ;
      RECT 10.906 0.152 10.982 8.116 ;
      RECT 11.818 0.152 11.894 8.116 ;
      RECT 13.186 0.152 13.262 8.116 ;
      RECT 13.794 0.152 13.87 8.116 ;
      RECT 13.946 0.152 14.022 1.1285 ;
      RECT 16.226 0.152 16.302 1.437 ;
      RECT 16.378 0.152 16.454 1.88 ;
      RECT 16.682 0.152 16.758 1.88 ;
      RECT 16.834 0.152 16.91 1.437 ;
      RECT 17.442 0.152 17.518 1.8795 ;
      RECT 18.354 0.152 18.43 8.116 ;
      RECT 18.658 0.152 18.734 8.116 ;
      RECT 18.81 0.152 18.886 8.116 ;
      RECT 19.114 0.152 19.19 8.116 ;
      RECT 19.703 0.152 19.817 8.154 ;
      RECT 20.026 0.152 20.102 8.116 ;
      RECT 20.33 0.152 20.406 8.116 ;
      RECT 20.482 0.152 20.558 8.116 ;
      RECT 20.634 0.152 20.71 8.116 ;
      RECT 20.919 0.152 21.033 8.154 ;
      RECT 21.242 0.152 21.318 8.116 ;
      RECT 21.85 0.152 21.926 8.116 ;
      RECT 22.002 0.152 22.078 1.8715 ;
      RECT 22.306 0.152 22.382 8.116 ;
      RECT 22.458 0.152 22.534 8.116 ;
      RECT 22.61 0.152 22.686 8.116 ;
      RECT 23.218 0.152 23.294 2.3845 ;
      RECT 23.37 0.152 23.446 1.878 ;
      RECT 23.674 0.152 23.75 2.9 ;
      RECT 23.978 0.152 24.054 1.212 ;
      RECT 27.17 0.152 27.246 8.116 ;
      RECT 27.778 0.152 27.854 8.116 ;
      RECT 28.538 0.152 28.614 2.3765 ;
      RECT 29.45 0.152 29.526 2.4215 ;
      RECT 34.618 0.152 34.694 2.404 ;
      RECT 34.922 0.152 34.998 1.641 ;
      RECT 35.53 0.152 35.606 2.505 ;
      RECT 37.81 0.152 37.886 5.099 ;
      RECT 37.962 0.152 38.038 5.219 ;
      RECT 38.114 0.152 38.19 0.4195 ;
      RECT 38.266 0.152 38.342 0.792 ;
      RECT 39.938 0.152 40.014 5.339 ;
      RECT 40.85 0.152 40.926 5.339 ;
      RECT 35.682 0.254 35.758 6.77 ;
      RECT 36.29 0.254 36.366 6.77 ;
      RECT 36.898 0.254 36.974 6.77 ;
      RECT 37.506 0.254 37.582 4.019 ;
      RECT 32.338 0.2745 32.414 6.77 ;
      RECT 32.946 0.2745 33.022 6.77 ;
      RECT 33.554 0.2745 33.63 6.77 ;
      RECT 34.466 0.2745 34.542 6.77 ;
      RECT 35.074 0.2745 35.15 6.77 ;
      RECT 3.154 0.2785 3.23 3.446 ;
      RECT 4.37 0.2785 4.446 3.446 ;
      RECT 4.978 0.2785 5.054 3.446 ;
      RECT 5.586 0.2785 5.662 3.446 ;
      RECT 6.194 0.2785 6.27 3.446 ;
      RECT 6.954 0.2785 7.03 3.4425 ;
      RECT 7.562 0.2785 7.638 3.4355 ;
      RECT 8.17 0.2785 8.246 6.77 ;
      RECT 8.778 0.2785 8.854 6.77 ;
      RECT 9.386 0.2785 9.462 6.77 ;
      RECT 10.146 0.2785 10.222 6.77 ;
      RECT 10.602 0.2785 10.678 6.77 ;
      RECT 10.754 0.2785 10.83 6.77 ;
      RECT 11.21 0.2785 11.286 6.77 ;
      RECT 11.362 0.2785 11.438 6.77 ;
      RECT 11.97 0.2785 12.046 6.77 ;
      RECT 12.578 0.2785 12.654 6.77 ;
      RECT 13.338 0.2785 13.414 8.3835 ;
      RECT 14.554 0.2785 14.63 6.77 ;
      RECT 16.53 0.2785 16.606 1.5605 ;
      RECT 17.594 0.2785 17.67 1.515 ;
      RECT 17.898 0.2785 17.974 4.019 ;
      RECT 24.13 0.2785 24.206 2.7615 ;
      RECT 24.738 0.2785 24.814 2.7615 ;
      RECT 25.346 0.2785 25.422 2.7615 ;
      RECT 26.106 0.2785 26.182 6.77 ;
      RECT 26.714 0.2785 26.79 6.77 ;
      RECT 27.322 0.2785 27.398 8.3835 ;
      RECT 27.93 0.2785 28.006 8.3835 ;
      RECT 28.69 0.2785 28.766 6.77 ;
      RECT 29.298 0.2785 29.374 6.77 ;
      RECT 29.906 0.2785 29.982 6.77 ;
      RECT 30.514 0.2785 30.59 6.77 ;
      RECT 31.122 0.2785 31.198 6.77 ;
      RECT 31.73 0.2785 31.806 6.77 ;
      RECT 38.114 0.6975 38.19 4.5 ;
      RECT 23.522 0.7155 23.598 2.22 ;
      RECT 25.802 0.7155 25.878 2.106 ;
      RECT 26.41 0.7155 26.486 5.77 ;
      RECT 27.018 0.7155 27.094 5.77 ;
      RECT 27.626 0.7155 27.702 5.77 ;
      RECT 28.234 0.7155 28.31 5.77 ;
      RECT 28.994 0.7155 29.07 5.77 ;
      RECT 29.602 0.7155 29.678 5.77 ;
      RECT 30.21 0.7155 30.286 5.77 ;
      RECT 30.818 0.7155 30.894 5.77 ;
      RECT 31.426 0.7155 31.502 5.77 ;
      RECT 32.034 0.7155 32.11 5.77 ;
      RECT 32.794 0.7155 32.87 5.77 ;
      RECT 33.402 0.7155 33.478 5.77 ;
      RECT 34.314 0.7155 34.39 5.77 ;
      RECT 34.77 0.7155 34.846 5.77 ;
      RECT 35.378 0.7155 35.454 5.77 ;
      RECT 37.658 0.7195 37.734 5.77 ;
      RECT 36.138 0.724 36.214 5.77 ;
      RECT 36.442 0.724 36.518 5.77 ;
      RECT 36.746 0.724 36.822 5.77 ;
      RECT 37.202 0.724 37.278 4.5035 ;
      RECT 10.45 0.761 10.526 5.7615 ;
      RECT 11.058 0.761 11.134 5.7615 ;
      RECT 11.666 0.761 11.742 5.7615 ;
      RECT 13.034 0.761 13.11 5.7615 ;
      RECT 13.642 0.761 13.718 5.7615 ;
      RECT 14.25 0.761 14.326 5.7615 ;
      RECT 14.858 0.761 14.934 5.7615 ;
      RECT 15.77 0.761 15.846 2.12 ;
      RECT 17.138 0.761 17.214 2.127 ;
      RECT 4.674 1.121 4.75 5.7615 ;
      RECT 5.282 1.121 5.358 5.7615 ;
      RECT 5.89 1.121 5.966 5.7615 ;
      RECT 13.946 1.241 14.022 6.77 ;
      RECT 38.418 1.259 38.494 36.4635 ;
      RECT 4.066 1.2785 4.142 5.7615 ;
      RECT 7.258 1.2785 7.334 5.7615 ;
      RECT 7.866 1.2785 7.942 5.7615 ;
      RECT 8.474 1.2785 8.55 5.7615 ;
      RECT 9.082 1.2785 9.158 5.7615 ;
      RECT 9.69 1.2785 9.766 5.7615 ;
      RECT 38.722 1.739 38.798 36.7145 ;
      RECT 38.874 1.859 38.95 36.8295 ;
      RECT 6.498 2.0295 6.574 5.7615 ;
      RECT 24.52 2.265 24.56 36.048 ;
      RECT 25.72 2.265 25.76 36.048 ;
      RECT 15.2455 2.268 15.2855 36.048 ;
      RECT 16.4455 2.268 16.4855 36.048 ;
      RECT 34.922 2.27 34.998 6.77 ;
      RECT 39.026 2.273 39.102 4.019 ;
      RECT 17.6455 2.274 17.6855 36.048 ;
      RECT 2.09 2.561 2.166 36.9655 ;
      RECT 39.33 2.699 39.406 37.1995 ;
      RECT 15.8455 2.781 15.8855 36.048 ;
      RECT 17.0455 2.781 17.0855 36.048 ;
      RECT 23.92 2.782 23.96 36.048 ;
      RECT 25.12 2.782 25.16 36.048 ;
      RECT 39.482 2.819 39.558 37.322 ;
      RECT 23.32 3.049 23.36 40.808 ;
      RECT 23.52 3.067 23.76 32.4145 ;
      RECT 24.12 3.067 24.36 32.412 ;
      RECT 24.72 3.067 24.96 32.412 ;
      RECT 25.32 3.067 25.56 32.412 ;
      RECT 15.4455 3.088 15.6855 32.412 ;
      RECT 16.0455 3.088 16.2855 32.412 ;
      RECT 16.6455 3.088 16.8855 32.412 ;
      RECT 17.2455 3.088 17.4855 32.412 ;
      RECT 10.298 3.16 10.374 5.7615 ;
      RECT 2.546 3.161 2.622 37.3255 ;
      RECT 39.634 3.161 39.71 37.415 ;
      RECT 35.53 3.259 35.606 6.77 ;
      RECT 38.57 3.273 38.646 4.5 ;
      RECT 39.178 3.273 39.254 4.5 ;
      RECT 35.853 3.401 35.891 3.539 ;
      RECT 35.853 3.641 35.891 3.779 ;
      RECT 1.786 3.761 1.862 36.7135 ;
      RECT 22.781 3.761 22.819 4.019 ;
      RECT 18.962 3.8565 19.038 8.3835 ;
      RECT 22.002 3.8565 22.078 8.3835 ;
      RECT 35.986 3.876 36.062 6.77 ;
      RECT 36.594 3.876 36.67 6.77 ;
      RECT 21.546 3.969 21.622 7.097 ;
      RECT 21.698 3.969 21.774 7.097 ;
      RECT 22.154 3.969 22.23 7.097 ;
      RECT 19.418 3.989 19.494 8.116 ;
      RECT 1.482 4.001 1.558 36.4715 ;
      RECT 1.938 4.001 2.014 36.8395 ;
      RECT 35.834 4.103 35.91 5.77 ;
      RECT 39.026 4.118 39.102 36.9505 ;
      RECT 1.634 4.121 1.71 36.5855 ;
      RECT 2.394 4.361 2.47 37.1955 ;
      RECT 38.266 4.481 38.342 37.415 ;
      RECT 39.178 4.6 39.254 37.0595 ;
      RECT 2.698 4.601 2.774 37.415 ;
      POLYGON 23.2 4.721 23.2 60.5315 23 60.5315 23 20.33 23.124 20.33 23.124 4.721 ;
      RECT 39.786 4.841 39.862 34.869 ;
      RECT 2.242 4.961 2.318 37.0835 ;
      POLYGON 17.9175 5.0165 17.9175 20.3235 18.0375 20.3235 18.0375 60.5315 17.8375 60.5315 17.8375 5.0165 ;
      RECT 38.57 5.201 38.646 36.59 ;
      RECT 37.4845 6.27 37.6845 23.237 ;
      RECT 37.835 7.225 37.915 31.728 ;
      RECT 3.285 8.28 3.365 28.768 ;
      RECT 27.04 10.131 27.12 19.529 ;
      RECT 26.88 18.84 26.96 19.529 ;
      RECT 28.202 19.75 28.282 36.048 ;
      RECT 26.9505 19.763 27.1505 36.048 ;
      RECT 18.7095 23.564 18.7895 29.977 ;
      RECT 19.1 23.564 19.3 29.977 ;
      RECT 19.6105 23.564 19.6905 29.977 ;
      RECT 21.0925 23.564 21.1725 29.977 ;
      RECT 21.6735 23.564 21.7535 29.977 ;
      RECT 22.064 23.564 22.264 29.977 ;
      RECT 22.5745 23.564 22.6545 29.977 ;
      RECT 27.6915 23.564 27.8915 36.048 ;
      RECT 35.1015 23.57 35.3015 36.77 ;
      RECT 35.612 23.57 35.692 31.417 ;
      RECT 36.5835 23.57 36.7835 31.417 ;
      RECT 37.4845 23.57 37.6845 31.417 ;
      RECT 36.193 23.572 36.273 31.417 ;
      RECT 37.094 23.572 37.174 31.417 ;
      RECT 8.7525 24.271 8.8525 24.769 ;
      RECT 11.7165 24.271 11.8165 24.769 ;
      RECT 14.6805 24.271 14.7805 24.769 ;
      RECT 26.2595 24.271 26.3595 24.769 ;
      RECT 29.2235 24.271 29.3235 24.769 ;
      RECT 32.1875 24.271 32.2875 24.769 ;
      RECT 7.752 24.2785 7.79 24.7615 ;
      RECT 9.8145 24.2785 9.8525 24.7615 ;
      RECT 10.716 24.2785 10.754 24.7615 ;
      RECT 12.779 24.2785 12.817 24.7615 ;
      RECT 13.68 24.2785 13.718 24.7615 ;
      RECT 27.322 24.2785 27.36 24.7615 ;
      RECT 30.286 24.2785 30.324 24.7615 ;
      RECT 31.187 24.2785 31.225 24.7615 ;
      RECT 33.25 24.2785 33.288 24.7615 ;
      RECT 34.151 24.2785 34.189 24.7615 ;
      RECT 0.57 28.571 0.646 35.411 ;
      RECT 0.722 28.571 0.798 35.411 ;
      RECT 0.874 28.571 0.95 35.411 ;
      RECT 1.026 28.571 1.102 35.411 ;
      RECT 1.178 28.571 1.254 35.411 ;
      RECT 1.33 28.571 1.406 35.411 ;
      RECT 2.85 28.571 2.926 35.411 ;
      RECT 18.158 30.123 18.198 40.808 ;
      RECT 19.119 30.123 19.159 40.808 ;
      RECT 20.08 30.123 20.12 40.808 ;
      RECT 20.92 30.123 20.96 40.808 ;
      RECT 21.88 30.123 21.92 40.808 ;
      RECT 22.84 30.123 22.88 40.808 ;
      RECT 18.3185 30.372 18.5185 59.007 ;
      RECT 22.52 30.372 22.72 59.001 ;
      RECT 36.5835 31.952 36.7835 38.152 ;
      RECT 36.193 31.971 36.273 38.1275 ;
      RECT 36.353 31.971 36.433 32.77 ;
      RECT 40.062 32.988 40.262 35.79 ;
      RECT 40.462 32.988 40.662 35.79 ;
      RECT 0.114 36.346 0.194 62.5775 ;
      RECT 40.85 36.346 40.926 63.0035 ;
      RECT 40.698 36.436 40.774 63.0035 ;
      RECT 0.274 36.4435 0.354 62.5775 ;
      RECT 0.434 36.5505 0.514 62.5775 ;
      RECT 40.546 36.555 40.622 63.0035 ;
      RECT 0.594 36.6655 0.674 62.5775 ;
      RECT 40.394 36.679 40.47 63.0035 ;
      RECT 0.754 36.7415 0.834 62.5775 ;
      RECT 40.242 36.794 40.318 63.0035 ;
      RECT 0.914 36.886 0.994 62.5775 ;
      RECT 40.09 36.916 40.166 63.0035 ;
      RECT 1.074 36.9995 1.154 62.5775 ;
      RECT 39.938 37.04 40.014 63.0035 ;
      RECT 1.234 37.1225 1.314 62.5775 ;
      RECT 1.394 37.248 1.474 62.5775 ;
      RECT 10.003 40.846 10.061 41.782 ;
      RECT 30.979 40.846 31.037 41.782 ;
      RECT 18.158 41.336 18.198 59.2585 ;
      RECT 39.786 42.639 39.862 62.6135 ;
      RECT 20.081 43.8425 20.119 43.9805 ;
      RECT 20.921 43.8425 20.959 43.9805 ;
      RECT 20.081 44.561 20.119 44.699 ;
      RECT 2.479 50.418 2.537 51.3315 ;
      RECT 2.707 50.418 2.765 51.3315 ;
      RECT 2.935 50.418 2.993 51.3315 ;
      RECT 3.163 50.418 3.221 51.3315 ;
      RECT 3.391 50.418 3.449 51.3315 ;
      RECT 3.619 50.418 3.677 51.3315 ;
      RECT 3.847 50.418 3.905 51.3315 ;
      RECT 4.075 50.418 4.133 51.3315 ;
      RECT 4.303 50.418 4.361 51.3315 ;
      RECT 4.531 50.418 4.589 51.3315 ;
      RECT 4.759 50.418 4.817 51.3315 ;
      RECT 4.987 50.418 5.045 51.3315 ;
      RECT 5.215 50.418 5.273 51.3315 ;
      RECT 5.443 50.418 5.501 51.3315 ;
      RECT 5.671 50.418 5.729 51.3315 ;
      RECT 5.899 50.418 5.957 51.3315 ;
      RECT 6.127 50.418 6.185 51.3315 ;
      RECT 6.355 50.418 6.413 51.3315 ;
      RECT 6.583 50.418 6.641 51.3315 ;
      RECT 6.811 50.418 6.869 51.3315 ;
      RECT 7.039 50.418 7.097 51.3315 ;
      RECT 7.267 50.418 7.325 51.3315 ;
      RECT 7.495 50.418 7.553 51.3315 ;
      RECT 7.723 50.418 7.781 51.3315 ;
      RECT 7.951 50.418 8.009 51.3315 ;
      RECT 8.179 50.418 8.237 51.3315 ;
      RECT 8.407 50.418 8.465 51.3315 ;
      RECT 8.635 50.418 8.693 51.3315 ;
      RECT 8.863 50.418 8.921 51.3315 ;
      RECT 9.091 50.418 9.149 51.3315 ;
      RECT 9.319 50.418 9.377 51.3315 ;
      RECT 9.547 50.418 9.605 51.3315 ;
      RECT 10.003 50.418 10.061 51.3315 ;
      RECT 10.231 50.418 10.289 51.3315 ;
      RECT 10.459 50.418 10.517 51.3315 ;
      RECT 10.687 50.418 10.745 51.3315 ;
      RECT 10.915 50.418 10.973 51.3315 ;
      RECT 11.143 50.418 11.201 51.3315 ;
      RECT 11.371 50.418 11.429 51.3315 ;
      RECT 11.599 50.418 11.657 51.3315 ;
      RECT 11.827 50.418 11.885 51.3315 ;
      RECT 12.055 50.418 12.113 51.3315 ;
      RECT 12.283 50.418 12.341 51.3315 ;
      RECT 12.511 50.418 12.569 51.3315 ;
      RECT 12.739 50.418 12.797 51.3315 ;
      RECT 12.967 50.418 13.025 51.3315 ;
      RECT 13.195 50.418 13.253 51.3315 ;
      RECT 13.423 50.418 13.481 51.3315 ;
      RECT 13.651 50.418 13.709 51.3315 ;
      RECT 13.879 50.418 13.937 51.3315 ;
      RECT 14.107 50.418 14.165 51.3315 ;
      RECT 14.335 50.418 14.393 51.3315 ;
      RECT 14.563 50.418 14.621 51.3315 ;
      RECT 14.791 50.418 14.849 51.3315 ;
      RECT 15.019 50.418 15.077 51.3315 ;
      RECT 15.247 50.418 15.305 51.3315 ;
      RECT 15.475 50.418 15.533 51.3315 ;
      RECT 15.703 50.418 15.761 51.3315 ;
      RECT 15.931 50.418 15.989 51.3315 ;
      RECT 16.159 50.418 16.217 51.3315 ;
      RECT 16.387 50.418 16.445 51.3315 ;
      RECT 16.615 50.418 16.673 51.3315 ;
      RECT 16.843 50.418 16.901 51.3315 ;
      RECT 17.071 50.418 17.129 51.3315 ;
      RECT 23.911 50.418 23.969 51.3315 ;
      RECT 24.139 50.418 24.197 51.3315 ;
      RECT 24.367 50.418 24.425 51.3315 ;
      RECT 24.595 50.418 24.653 51.3315 ;
      RECT 24.823 50.418 24.881 51.3315 ;
      RECT 25.051 50.418 25.109 51.3315 ;
      RECT 25.279 50.418 25.337 51.3315 ;
      RECT 25.507 50.418 25.565 51.3315 ;
      RECT 25.735 50.418 25.793 51.3315 ;
      RECT 25.963 50.418 26.021 51.3315 ;
      RECT 26.191 50.418 26.249 51.3315 ;
      RECT 26.419 50.418 26.477 51.3315 ;
      RECT 26.647 50.418 26.705 51.3315 ;
      RECT 26.875 50.418 26.933 51.3315 ;
      RECT 27.103 50.418 27.161 51.3315 ;
      RECT 27.331 50.418 27.389 51.3315 ;
      RECT 27.559 50.418 27.617 51.3315 ;
      RECT 27.787 50.418 27.845 51.3315 ;
      RECT 28.015 50.418 28.073 51.3315 ;
      RECT 28.243 50.418 28.301 51.3315 ;
      RECT 28.471 50.418 28.529 51.3315 ;
      RECT 28.699 50.418 28.757 51.3315 ;
      RECT 28.927 50.418 28.985 51.3315 ;
      RECT 29.155 50.418 29.213 51.3315 ;
      RECT 29.383 50.418 29.441 51.3315 ;
      RECT 29.611 50.418 29.669 51.3315 ;
      RECT 29.839 50.418 29.897 51.3315 ;
      RECT 30.067 50.418 30.125 51.3315 ;
      RECT 30.295 50.418 30.353 51.3315 ;
      RECT 30.523 50.418 30.581 51.3315 ;
      RECT 30.751 50.418 30.809 51.3315 ;
      RECT 30.979 50.418 31.037 51.3315 ;
      RECT 31.435 50.418 31.493 51.3315 ;
      RECT 31.663 50.418 31.721 51.3315 ;
      RECT 31.891 50.418 31.949 51.3315 ;
      RECT 32.119 50.418 32.177 51.3315 ;
      RECT 32.347 50.418 32.405 51.3315 ;
      RECT 32.575 50.418 32.633 51.3315 ;
      RECT 32.803 50.418 32.861 51.3315 ;
      RECT 33.031 50.418 33.089 51.3315 ;
      RECT 33.259 50.418 33.317 51.3315 ;
      RECT 33.487 50.418 33.545 51.3315 ;
      RECT 33.715 50.418 33.773 51.3315 ;
      RECT 33.943 50.418 34.001 51.3315 ;
      RECT 34.171 50.418 34.229 51.3315 ;
      RECT 34.399 50.418 34.457 51.3315 ;
      RECT 34.627 50.418 34.685 51.3315 ;
      RECT 34.855 50.418 34.913 51.3315 ;
      RECT 35.083 50.418 35.141 51.3315 ;
      RECT 35.311 50.418 35.369 51.3315 ;
      RECT 35.539 50.418 35.597 51.3315 ;
      RECT 35.767 50.418 35.825 51.3315 ;
      RECT 35.995 50.418 36.053 51.3315 ;
      RECT 36.223 50.418 36.281 51.3315 ;
      RECT 36.451 50.418 36.509 51.3315 ;
      RECT 36.679 50.418 36.737 51.3315 ;
      RECT 36.907 50.418 36.965 51.3315 ;
      RECT 37.135 50.418 37.193 51.3315 ;
      RECT 37.363 50.418 37.421 51.3315 ;
      RECT 37.591 50.418 37.649 51.3315 ;
      RECT 37.819 50.418 37.877 51.3315 ;
      RECT 38.047 50.418 38.105 51.3315 ;
      RECT 38.275 50.418 38.333 51.3315 ;
      RECT 38.503 50.418 38.561 51.3315 ;
      RECT 2.479 51.446 2.537 52.252 ;
      RECT 2.707 51.446 2.765 52.252 ;
      RECT 2.935 51.446 2.993 52.252 ;
      RECT 3.163 51.446 3.221 52.252 ;
      RECT 3.391 51.446 3.449 52.252 ;
      RECT 3.619 51.446 3.677 52.252 ;
      RECT 3.847 51.446 3.905 52.252 ;
      RECT 4.075 51.446 4.133 52.252 ;
      RECT 4.303 51.446 4.361 52.252 ;
      RECT 4.531 51.446 4.589 52.252 ;
      RECT 4.759 51.446 4.817 52.252 ;
      RECT 4.987 51.446 5.045 52.252 ;
      RECT 5.215 51.446 5.273 52.252 ;
      RECT 5.443 51.446 5.501 52.252 ;
      RECT 5.671 51.446 5.729 52.252 ;
      RECT 5.899 51.446 5.957 52.252 ;
      RECT 6.127 51.446 6.185 52.252 ;
      RECT 6.355 51.446 6.413 52.252 ;
      RECT 6.583 51.446 6.641 52.252 ;
      RECT 6.811 51.446 6.869 52.252 ;
      RECT 7.039 51.446 7.097 52.252 ;
      RECT 7.267 51.446 7.325 52.252 ;
      RECT 7.495 51.446 7.553 52.252 ;
      RECT 7.723 51.446 7.781 52.252 ;
      RECT 7.951 51.446 8.009 52.252 ;
      RECT 8.179 51.446 8.237 52.252 ;
      RECT 8.407 51.446 8.465 52.252 ;
      RECT 8.635 51.446 8.693 52.252 ;
      RECT 8.863 51.446 8.921 52.252 ;
      RECT 9.091 51.446 9.149 52.252 ;
      RECT 9.319 51.446 9.377 52.252 ;
      RECT 9.547 51.446 9.605 52.252 ;
      RECT 10.003 51.446 10.061 52.252 ;
      RECT 10.231 51.446 10.289 52.252 ;
      RECT 10.459 51.446 10.517 52.252 ;
      RECT 10.687 51.446 10.745 52.252 ;
      RECT 10.915 51.446 10.973 52.252 ;
      RECT 11.143 51.446 11.201 52.252 ;
      RECT 11.371 51.446 11.429 52.252 ;
      RECT 11.599 51.446 11.657 52.252 ;
      RECT 11.827 51.446 11.885 52.252 ;
      RECT 12.055 51.446 12.113 52.252 ;
      RECT 12.283 51.446 12.341 52.252 ;
      RECT 12.511 51.446 12.569 52.252 ;
      RECT 12.739 51.446 12.797 52.252 ;
      RECT 12.967 51.446 13.025 52.252 ;
      RECT 13.195 51.446 13.253 52.252 ;
      RECT 13.423 51.446 13.481 52.252 ;
      RECT 13.651 51.446 13.709 52.252 ;
      RECT 13.879 51.446 13.937 52.252 ;
      RECT 14.107 51.446 14.165 52.252 ;
      RECT 14.335 51.446 14.393 52.252 ;
      RECT 14.563 51.446 14.621 52.252 ;
      RECT 14.791 51.446 14.849 52.252 ;
      RECT 15.019 51.446 15.077 52.252 ;
      RECT 15.247 51.446 15.305 52.252 ;
      RECT 15.475 51.446 15.533 52.252 ;
      RECT 15.703 51.446 15.761 52.252 ;
      RECT 15.931 51.446 15.989 52.252 ;
      RECT 16.159 51.446 16.217 52.252 ;
      RECT 16.387 51.446 16.445 52.252 ;
      RECT 16.615 51.446 16.673 52.252 ;
      RECT 16.843 51.446 16.901 52.252 ;
      RECT 17.071 51.446 17.129 52.252 ;
      RECT 23.911 51.446 23.969 52.252 ;
      RECT 24.139 51.446 24.197 52.252 ;
      RECT 24.367 51.446 24.425 52.252 ;
      RECT 24.595 51.446 24.653 52.252 ;
      RECT 24.823 51.446 24.881 52.252 ;
      RECT 25.051 51.446 25.109 52.252 ;
      RECT 25.279 51.446 25.337 52.252 ;
      RECT 25.507 51.446 25.565 52.252 ;
      RECT 25.735 51.446 25.793 52.252 ;
      RECT 25.963 51.446 26.021 52.252 ;
      RECT 26.191 51.446 26.249 52.252 ;
      RECT 26.419 51.446 26.477 52.252 ;
      RECT 26.647 51.446 26.705 52.252 ;
      RECT 26.875 51.446 26.933 52.252 ;
      RECT 27.103 51.446 27.161 52.252 ;
      RECT 27.331 51.446 27.389 52.252 ;
      RECT 27.559 51.446 27.617 52.252 ;
      RECT 27.787 51.446 27.845 52.252 ;
      RECT 28.015 51.446 28.073 52.252 ;
      RECT 28.243 51.446 28.301 52.252 ;
      RECT 28.471 51.446 28.529 52.252 ;
      RECT 28.699 51.446 28.757 52.252 ;
      RECT 28.927 51.446 28.985 52.252 ;
      RECT 29.155 51.446 29.213 52.252 ;
      RECT 29.383 51.446 29.441 52.252 ;
      RECT 29.611 51.446 29.669 52.252 ;
      RECT 29.839 51.446 29.897 52.252 ;
      RECT 30.067 51.446 30.125 52.252 ;
      RECT 30.295 51.446 30.353 52.252 ;
      RECT 30.523 51.446 30.581 52.252 ;
      RECT 30.751 51.446 30.809 52.252 ;
      RECT 30.979 51.446 31.037 52.252 ;
      RECT 31.435 51.446 31.493 52.252 ;
      RECT 31.663 51.446 31.721 52.252 ;
      RECT 31.891 51.446 31.949 52.252 ;
      RECT 32.119 51.446 32.177 52.252 ;
      RECT 32.347 51.446 32.405 52.252 ;
      RECT 32.575 51.446 32.633 52.252 ;
      RECT 32.803 51.446 32.861 52.252 ;
      RECT 33.031 51.446 33.089 52.252 ;
      RECT 33.259 51.446 33.317 52.252 ;
      RECT 33.487 51.446 33.545 52.252 ;
      RECT 33.715 51.446 33.773 52.252 ;
      RECT 33.943 51.446 34.001 52.252 ;
      RECT 34.171 51.446 34.229 52.252 ;
      RECT 34.399 51.446 34.457 52.252 ;
      RECT 34.627 51.446 34.685 52.252 ;
      RECT 34.855 51.446 34.913 52.252 ;
      RECT 35.083 51.446 35.141 52.252 ;
      RECT 35.311 51.446 35.369 52.252 ;
      RECT 35.539 51.446 35.597 52.252 ;
      RECT 35.767 51.446 35.825 52.252 ;
      RECT 35.995 51.446 36.053 52.252 ;
      RECT 36.223 51.446 36.281 52.252 ;
      RECT 36.451 51.446 36.509 52.252 ;
      RECT 36.679 51.446 36.737 52.252 ;
      RECT 36.907 51.446 36.965 52.252 ;
      RECT 37.135 51.446 37.193 52.252 ;
      RECT 37.363 51.446 37.421 52.252 ;
      RECT 37.591 51.446 37.649 52.252 ;
      RECT 37.819 51.446 37.877 52.252 ;
      RECT 38.047 51.446 38.105 52.252 ;
      RECT 38.275 51.446 38.333 52.252 ;
      RECT 38.503 51.446 38.561 52.252 ;
      RECT 20.081 52.461 20.119 52.599 ;
      RECT 20.921 52.461 20.959 52.599 ;
      RECT 20.081 52.621 20.119 52.759 ;
      RECT 20.921 52.621 20.959 52.759 ;
      RECT 21.881 52.621 21.919 52.759 ;
      RECT 22.841 52.621 22.879 52.759 ;
      RECT 18.325 60.4585 18.383 61.454 ;
      RECT 22.657 60.4585 22.715 61.454 ;
      RECT 17.983 61.356 18.041 62.3085 ;
      RECT 18.439 61.356 18.497 62.3085 ;
      RECT 19.123 61.356 19.181 62.3085 ;
      RECT 20.035 61.356 20.093 62.3085 ;
      RECT 20.947 61.356 21.005 62.3085 ;
      RECT 21.859 61.356 21.917 62.3085 ;
      RECT 22.543 61.356 22.601 62.3085 ;
      RECT 22.999 61.356 23.057 62.3085 ;
      RECT 10.003 61.358 10.061 62.294 ;
      RECT 30.979 61.358 31.037 62.294 ;
      RECT 0.3 66.375 20.28 66.825 ;
      RECT 20.76 66.375 40.74 66.825 ;
      RECT 5.6 68.175 20.28 68.625 ;
      RECT 20.76 68.175 35.44 68.625 ;
      RECT 0.3 69.075 20.28 69.525 ;
      RECT 20.76 69.075 40.74 69.525 ;
      RECT 5.6 69.975 20.28 70.425 ;
      RECT 20.76 69.975 35.44 70.425 ;
      RECT 0.3 70.875 20.28 71.325 ;
      RECT 20.76 70.875 40.74 71.325 ;
      RECT 5.6 71.775 20.28 72.225 ;
      RECT 20.76 71.775 35.44 72.225 ;
      RECT 0.3 72.675 20.28 73.125 ;
      RECT 20.76 72.675 40.74 73.125 ;
      RECT 5.6 73.575 20.28 74.025 ;
      RECT 20.76 73.575 35.44 74.025 ;
      RECT 0.3 74.475 20.28 74.925 ;
      RECT 20.76 74.475 40.74 74.925 ;
      RECT 5.6 75.375 20.28 75.825 ;
      RECT 20.76 75.375 35.44 75.825 ;
      RECT 0.3 76.275 20.28 76.725 ;
      RECT 20.76 76.275 40.74 76.725 ;
      RECT 0.3 77.175 20.28 77.625 ;
      RECT 20.76 77.175 40.74 77.625 ;
      RECT 0.3 78.075 20.28 78.525 ;
      RECT 20.76 78.075 40.74 78.525 ;
      RECT 0.3 78.975 20.28 79.425 ;
      RECT 20.76 78.975 40.74 79.425 ;
      RECT 5.601 79.875 20.28 80.325 ;
      RECT 20.76 79.875 35.439 80.325 ;
      RECT 0.3 80.775 20.28 81.225 ;
      RECT 20.76 80.775 40.74 81.225 ;
      RECT 5.601 81.675 20.28 82.125 ;
      RECT 20.76 81.675 35.439 82.125 ;
      RECT 0.3 82.575 20.28 83.025 ;
      RECT 20.76 82.575 40.74 83.025 ;
      RECT 5.601 83.475 20.28 83.925 ;
      RECT 20.76 83.475 35.439 83.925 ;
      RECT 0.3 84.375 20.28 84.825 ;
      RECT 20.76 84.375 40.74 84.825 ;
      RECT 5.601 85.275 20.28 85.725 ;
      RECT 20.76 85.275 35.439 85.725 ;
      RECT 0.3 86.175 20.28 86.625 ;
      RECT 20.76 86.175 40.74 86.625 ;
      RECT 5.601 87.075 20.28 87.525 ;
      RECT 20.76 87.075 35.439 87.525 ;
    LAYER M6 ;
      RECT 5.495 31.27 6.019 31.77 ;
    LAYER M5 ;
      RECT 3.61 0.152 3.686 1.253 ;
      RECT 6.802 0.152 6.878 3.3705 ;
      RECT 7.41 0.152 7.486 1.5595 ;
      RECT 16.074 0.152 16.15 1.437 ;
      RECT 16.986 0.152 17.062 1.437 ;
      RECT 17.29 0.152 17.366 1.437 ;
      RECT 23.066 0.152 23.142 1.437 ;
      RECT 23.826 0.152 23.902 1.212 ;
      RECT 24.282 0.152 24.358 1.437 ;
      RECT 28.842 0.152 28.918 1.8805 ;
      RECT 29.146 0.152 29.222 1.8685 ;
      RECT 35.226 0.152 35.302 1.3065 ;
      RECT 3.458 1.2785 3.534 4.502 ;
      RECT 3.762 1.351 3.838 3.446 ;
      RECT 23.066 1.802 23.142 3.7725 ;
      RECT 28.842 2.7115 28.918 5.77 ;
      RECT 18.6385 30.123 18.6785 42.7 ;
      RECT 19.5995 30.123 19.6395 42.7445 ;
      RECT 21.4 30.123 21.44 42.7375 ;
      RECT 22.36 30.123 22.4 42.7375 ;
      RECT 18.799 30.372 18.999 59.282 ;
      RECT 19.2795 30.372 19.4795 59.007 ;
      RECT 19.76 30.372 19.96 59.007 ;
      RECT 21.08 30.372 21.28 59.0065 ;
      RECT 21.56 30.372 21.76 59.007 ;
      RECT 22.04 30.372 22.24 59.007 ;
      RECT 13.537 37.806 13.595 39.7865 ;
      RECT 13.765 37.806 13.823 39.7865 ;
      RECT 13.993 37.806 14.051 39.7865 ;
      RECT 14.221 37.806 14.279 39.7865 ;
      RECT 14.449 37.806 14.507 39.7865 ;
      RECT 14.677 37.806 14.735 39.7865 ;
      RECT 14.905 37.806 14.963 39.7865 ;
      RECT 15.133 37.806 15.191 39.7865 ;
      RECT 15.361 37.806 15.419 39.7865 ;
      RECT 15.589 37.806 15.647 39.7865 ;
      RECT 15.817 37.806 15.875 39.7865 ;
      RECT 16.045 37.806 16.103 39.7865 ;
      RECT 16.273 37.806 16.331 39.7865 ;
      RECT 16.843 37.806 16.901 40.5965 ;
      RECT 17.071 37.806 17.129 40.5965 ;
      RECT 17.299 37.806 17.357 40.5965 ;
      RECT 23.683 37.806 23.741 40.5965 ;
      RECT 23.911 37.806 23.969 40.5965 ;
      RECT 24.139 37.806 24.197 40.5965 ;
      RECT 24.709 37.806 24.767 39.7865 ;
      RECT 24.937 37.806 24.995 39.7865 ;
      RECT 25.165 37.806 25.223 39.7865 ;
      RECT 25.393 37.806 25.451 39.7865 ;
      RECT 25.621 37.806 25.679 39.7865 ;
      RECT 25.849 37.806 25.907 39.7865 ;
      RECT 26.077 37.806 26.135 39.7865 ;
      RECT 26.305 37.806 26.363 39.7865 ;
      RECT 26.533 37.806 26.591 39.7865 ;
      RECT 26.761 37.806 26.819 39.7865 ;
      RECT 26.989 37.806 27.047 39.7865 ;
      RECT 27.217 37.806 27.275 39.7865 ;
      RECT 27.445 37.806 27.503 39.7865 ;
      RECT 1.681 40.1685 1.739 41.584 ;
      RECT 1.909 40.1685 1.967 41.584 ;
      RECT 2.137 40.1685 2.195 41.584 ;
      RECT 2.365 40.1685 2.423 41.584 ;
      RECT 2.593 40.1685 2.651 41.584 ;
      RECT 2.821 40.1685 2.879 41.584 ;
      RECT 3.049 40.1685 3.107 41.584 ;
      RECT 3.277 40.1685 3.335 41.584 ;
      RECT 3.505 40.1685 3.563 41.584 ;
      RECT 3.733 40.1685 3.791 41.584 ;
      RECT 3.961 40.1685 4.019 41.584 ;
      RECT 37.021 40.1685 37.079 41.584 ;
      RECT 37.249 40.1685 37.307 41.584 ;
      RECT 37.477 40.1685 37.535 41.584 ;
      RECT 37.705 40.1685 37.763 41.584 ;
      RECT 37.933 40.1685 37.991 41.584 ;
      RECT 38.161 40.1685 38.219 41.584 ;
      RECT 38.389 40.1685 38.447 41.584 ;
      RECT 38.617 40.1685 38.675 41.584 ;
      RECT 38.845 40.1685 38.903 41.584 ;
      RECT 39.073 40.1685 39.131 41.584 ;
      RECT 39.301 40.1685 39.359 41.584 ;
      RECT 17.6775 40.7205 17.7175 59.2585 ;
      RECT 4.759 40.831 4.817 41.7815 ;
      RECT 4.987 40.831 5.045 41.7815 ;
      RECT 5.215 40.831 5.273 41.7815 ;
      RECT 5.443 40.831 5.501 41.7815 ;
      RECT 5.671 40.831 5.729 41.7815 ;
      RECT 5.899 40.831 5.957 41.7815 ;
      RECT 6.127 40.831 6.185 41.7815 ;
      RECT 6.355 40.831 6.413 41.7815 ;
      RECT 6.583 40.831 6.641 41.7815 ;
      RECT 6.811 40.831 6.869 41.7815 ;
      RECT 7.039 40.831 7.097 41.7815 ;
      RECT 7.267 40.831 7.325 41.7815 ;
      RECT 7.495 40.831 7.553 41.7815 ;
      RECT 7.723 40.831 7.781 41.7815 ;
      RECT 7.951 40.831 8.009 41.7815 ;
      RECT 8.179 40.831 8.237 41.7815 ;
      RECT 8.407 40.831 8.465 41.7815 ;
      RECT 8.635 40.831 8.693 41.7815 ;
      RECT 8.863 40.831 8.921 41.7815 ;
      RECT 9.091 40.831 9.149 41.7815 ;
      RECT 9.319 40.831 9.377 41.7815 ;
      RECT 9.547 40.831 9.605 41.7815 ;
      RECT 9.775 40.831 9.833 41.7815 ;
      RECT 10.231 40.831 10.289 41.7815 ;
      RECT 10.459 40.831 10.517 42.0585 ;
      RECT 10.687 40.831 10.745 41.7815 ;
      RECT 10.915 40.831 10.973 41.7815 ;
      RECT 11.143 40.831 11.201 41.7815 ;
      RECT 11.371 40.831 11.429 41.7815 ;
      RECT 11.599 40.831 11.657 41.7815 ;
      RECT 11.827 40.831 11.885 41.7815 ;
      RECT 12.055 40.831 12.113 41.7815 ;
      RECT 12.283 40.831 12.341 41.7815 ;
      RECT 12.511 40.831 12.569 41.7815 ;
      RECT 12.739 40.831 12.797 41.7815 ;
      RECT 12.967 40.831 13.025 41.7815 ;
      RECT 13.195 40.831 13.253 41.7815 ;
      RECT 13.423 40.831 13.481 41.7815 ;
      RECT 13.651 40.831 13.709 41.7815 ;
      RECT 13.879 40.831 13.937 41.7815 ;
      RECT 14.107 40.831 14.165 41.7815 ;
      RECT 14.335 40.831 14.393 41.7815 ;
      RECT 14.563 40.831 14.621 41.7815 ;
      RECT 14.791 40.831 14.849 41.7815 ;
      RECT 15.019 40.831 15.077 41.7815 ;
      RECT 15.247 40.831 15.305 41.7815 ;
      RECT 15.475 40.831 15.533 41.7815 ;
      RECT 15.703 40.831 15.761 41.7815 ;
      RECT 15.931 40.831 15.989 41.7815 ;
      RECT 16.159 40.831 16.217 41.7815 ;
      RECT 16.387 40.831 16.445 41.7815 ;
      RECT 16.615 40.831 16.673 41.7815 ;
      RECT 16.843 40.831 16.901 41.7815 ;
      RECT 24.139 40.831 24.197 41.7815 ;
      RECT 24.367 40.831 24.425 41.7815 ;
      RECT 24.595 40.831 24.653 41.7815 ;
      RECT 24.823 40.831 24.881 41.7815 ;
      RECT 25.051 40.831 25.109 41.7815 ;
      RECT 25.279 40.831 25.337 41.7815 ;
      RECT 25.507 40.831 25.565 41.7815 ;
      RECT 25.735 40.831 25.793 41.7815 ;
      RECT 25.963 40.831 26.021 41.7815 ;
      RECT 26.191 40.831 26.249 41.7815 ;
      RECT 26.419 40.831 26.477 41.7815 ;
      RECT 26.647 40.831 26.705 41.7815 ;
      RECT 26.875 40.831 26.933 41.7815 ;
      RECT 27.103 40.831 27.161 41.7815 ;
      RECT 27.331 40.831 27.389 41.7815 ;
      RECT 27.559 40.831 27.617 41.7815 ;
      RECT 27.787 40.831 27.845 41.7815 ;
      RECT 28.015 40.831 28.073 41.7815 ;
      RECT 28.243 40.831 28.301 41.7815 ;
      RECT 28.471 40.831 28.529 41.7815 ;
      RECT 28.699 40.831 28.757 41.7815 ;
      RECT 28.927 40.831 28.985 41.7815 ;
      RECT 29.155 40.831 29.213 41.7815 ;
      RECT 29.383 40.831 29.441 41.7815 ;
      RECT 29.611 40.831 29.669 41.7815 ;
      RECT 29.839 40.831 29.897 41.7815 ;
      RECT 30.067 40.831 30.125 41.7815 ;
      RECT 30.295 40.831 30.353 41.7815 ;
      RECT 30.523 40.831 30.581 42.0585 ;
      RECT 30.751 40.831 30.809 41.7815 ;
      RECT 31.207 40.831 31.265 41.7815 ;
      RECT 31.435 40.831 31.493 41.7815 ;
      RECT 31.663 40.831 31.721 41.7815 ;
      RECT 31.891 40.831 31.949 41.7815 ;
      RECT 32.119 40.831 32.177 41.7815 ;
      RECT 32.347 40.831 32.405 41.7815 ;
      RECT 32.575 40.831 32.633 41.7815 ;
      RECT 32.803 40.831 32.861 41.7815 ;
      RECT 33.031 40.831 33.089 41.7815 ;
      RECT 33.259 40.831 33.317 41.7815 ;
      RECT 33.487 40.831 33.545 41.7815 ;
      RECT 33.715 40.831 33.773 41.7815 ;
      RECT 33.943 40.831 34.001 41.7815 ;
      RECT 34.171 40.831 34.229 41.7815 ;
      RECT 34.399 40.831 34.457 41.7815 ;
      RECT 34.627 40.831 34.685 41.7815 ;
      RECT 34.855 40.831 34.913 41.7815 ;
      RECT 35.083 40.831 35.141 41.7815 ;
      RECT 35.311 40.831 35.369 41.7815 ;
      RECT 35.539 40.831 35.597 41.7815 ;
      RECT 35.767 40.831 35.825 41.7815 ;
      RECT 35.995 40.831 36.053 41.7815 ;
      RECT 36.223 40.831 36.281 41.7815 ;
      RECT 1.681 41.686 1.739 42.6815 ;
      RECT 1.909 41.686 1.967 42.6815 ;
      RECT 2.137 41.686 2.195 42.6815 ;
      RECT 2.365 41.686 2.423 42.6815 ;
      RECT 2.593 41.686 2.651 42.6815 ;
      RECT 2.821 41.686 2.879 42.6815 ;
      RECT 3.049 41.686 3.107 42.6815 ;
      RECT 3.277 41.686 3.335 42.6815 ;
      RECT 3.505 41.686 3.563 42.6815 ;
      RECT 3.733 41.686 3.791 42.6815 ;
      RECT 3.961 41.686 4.019 42.6815 ;
      RECT 4.189 41.686 4.247 42.6815 ;
      RECT 4.417 41.686 4.475 42.6815 ;
      RECT 4.645 41.686 4.703 42.6815 ;
      RECT 4.873 41.686 4.931 42.6815 ;
      RECT 5.101 41.686 5.159 42.6815 ;
      RECT 5.329 41.686 5.387 42.6815 ;
      RECT 5.557 41.686 5.615 42.6815 ;
      RECT 5.785 41.686 5.843 42.6815 ;
      RECT 6.013 41.686 6.071 42.6815 ;
      RECT 6.241 41.686 6.299 42.6815 ;
      RECT 6.469 41.686 6.527 42.6815 ;
      RECT 6.697 41.686 6.755 42.6815 ;
      RECT 6.925 41.686 6.983 42.6815 ;
      RECT 7.153 41.686 7.211 42.6815 ;
      RECT 7.381 41.686 7.439 42.6815 ;
      RECT 7.609 41.686 7.667 42.6815 ;
      RECT 7.837 41.686 7.895 42.6815 ;
      RECT 8.065 41.686 8.123 42.6815 ;
      RECT 8.293 41.686 8.351 42.6815 ;
      RECT 8.521 41.686 8.579 42.6815 ;
      RECT 8.749 41.686 8.807 42.6815 ;
      RECT 8.977 41.686 9.035 42.6815 ;
      RECT 9.205 41.686 9.263 42.6815 ;
      RECT 9.433 41.686 9.491 42.6815 ;
      RECT 9.661 41.686 9.719 42.6815 ;
      RECT 9.889 41.686 9.947 42.6815 ;
      RECT 10.117 41.686 10.175 42.6815 ;
      RECT 10.345 41.686 10.403 42.6815 ;
      RECT 10.573 41.686 10.631 42.6815 ;
      RECT 10.801 41.686 10.859 42.6815 ;
      RECT 11.029 41.686 11.087 42.6815 ;
      RECT 11.257 41.686 11.315 42.6815 ;
      RECT 11.485 41.686 11.543 42.6815 ;
      RECT 11.713 41.686 11.771 42.6815 ;
      RECT 11.941 41.686 11.999 42.6815 ;
      RECT 12.169 41.686 12.227 42.6815 ;
      RECT 12.397 41.686 12.455 42.6815 ;
      RECT 12.625 41.686 12.683 42.6815 ;
      RECT 12.853 41.686 12.911 42.6815 ;
      RECT 13.081 41.686 13.139 42.6815 ;
      RECT 13.309 41.686 13.367 42.6815 ;
      RECT 13.537 41.686 13.595 42.6815 ;
      RECT 13.765 41.686 13.823 42.6815 ;
      RECT 13.993 41.686 14.051 42.6815 ;
      RECT 14.221 41.686 14.279 42.6815 ;
      RECT 14.449 41.686 14.507 42.6815 ;
      RECT 14.677 41.686 14.735 42.6815 ;
      RECT 14.905 41.686 14.963 42.6815 ;
      RECT 15.133 41.686 15.191 42.6815 ;
      RECT 15.361 41.686 15.419 42.6815 ;
      RECT 15.589 41.686 15.647 42.6815 ;
      RECT 15.817 41.686 15.875 42.6815 ;
      RECT 16.045 41.686 16.103 42.6815 ;
      RECT 16.273 41.686 16.331 42.6815 ;
      RECT 16.501 41.686 16.559 42.6815 ;
      RECT 16.729 41.686 16.787 42.6815 ;
      RECT 24.253 41.686 24.311 42.6815 ;
      RECT 24.481 41.686 24.539 42.6815 ;
      RECT 24.709 41.686 24.767 42.6815 ;
      RECT 24.937 41.686 24.995 42.6815 ;
      RECT 25.165 41.686 25.223 42.6815 ;
      RECT 25.393 41.686 25.451 42.6815 ;
      RECT 25.621 41.686 25.679 42.6815 ;
      RECT 25.849 41.686 25.907 42.6815 ;
      RECT 26.077 41.686 26.135 42.6815 ;
      RECT 26.305 41.686 26.363 42.6815 ;
      RECT 26.533 41.686 26.591 42.6815 ;
      RECT 26.761 41.686 26.819 42.6815 ;
      RECT 26.989 41.686 27.047 42.6815 ;
      RECT 27.217 41.686 27.275 42.6815 ;
      RECT 27.445 41.686 27.503 42.6815 ;
      RECT 27.673 41.686 27.731 42.6815 ;
      RECT 27.901 41.686 27.959 42.6815 ;
      RECT 28.129 41.686 28.187 42.6815 ;
      RECT 28.357 41.686 28.415 42.6815 ;
      RECT 28.585 41.686 28.643 42.6815 ;
      RECT 28.813 41.686 28.871 42.6815 ;
      RECT 29.041 41.686 29.099 42.6815 ;
      RECT 29.269 41.686 29.327 42.6815 ;
      RECT 29.497 41.686 29.555 42.6815 ;
      RECT 29.725 41.686 29.783 42.6815 ;
      RECT 29.953 41.686 30.011 42.6815 ;
      RECT 30.181 41.686 30.239 42.6815 ;
      RECT 30.409 41.686 30.467 42.6815 ;
      RECT 30.637 41.686 30.695 42.6815 ;
      RECT 30.865 41.686 30.923 42.6815 ;
      RECT 31.093 41.686 31.151 42.6815 ;
      RECT 31.321 41.686 31.379 42.6815 ;
      RECT 31.549 41.686 31.607 42.6815 ;
      RECT 31.777 41.686 31.835 42.6815 ;
      RECT 32.005 41.686 32.063 42.6815 ;
      RECT 32.233 41.686 32.291 42.6815 ;
      RECT 32.461 41.686 32.519 42.6815 ;
      RECT 32.689 41.686 32.747 42.6815 ;
      RECT 32.917 41.686 32.975 42.6815 ;
      RECT 33.145 41.686 33.203 42.6815 ;
      RECT 33.373 41.686 33.431 42.6815 ;
      RECT 33.601 41.686 33.659 42.6815 ;
      RECT 33.829 41.686 33.887 42.6815 ;
      RECT 34.057 41.686 34.115 42.6815 ;
      RECT 34.285 41.686 34.343 42.6815 ;
      RECT 34.513 41.686 34.571 42.6815 ;
      RECT 34.741 41.686 34.799 42.6815 ;
      RECT 34.969 41.686 35.027 42.6815 ;
      RECT 35.197 41.686 35.255 42.6815 ;
      RECT 35.425 41.686 35.483 42.6815 ;
      RECT 35.653 41.686 35.711 42.6815 ;
      RECT 35.881 41.686 35.939 42.6815 ;
      RECT 36.109 41.686 36.167 42.6815 ;
      RECT 36.337 41.686 36.395 42.6815 ;
      RECT 36.565 41.686 36.623 42.6815 ;
      RECT 36.793 41.686 36.851 42.6815 ;
      RECT 37.021 41.686 37.079 42.6815 ;
      RECT 37.249 41.686 37.307 42.6815 ;
      RECT 37.477 41.686 37.535 42.6815 ;
      RECT 37.705 41.686 37.763 42.6815 ;
      RECT 37.933 41.686 37.991 42.6815 ;
      RECT 38.161 41.686 38.219 42.6815 ;
      RECT 38.389 41.686 38.447 42.6815 ;
      RECT 38.617 41.686 38.675 42.6815 ;
      RECT 38.845 41.686 38.903 42.6815 ;
      RECT 39.073 41.686 39.131 42.6815 ;
      RECT 39.301 41.686 39.359 42.6815 ;
      RECT 39.634 41.835 39.71 63.0035 ;
      RECT 17.3575 43.63 17.5575 46.8275 ;
      RECT 23.54 43.63 23.74 46.9 ;
      RECT 17.3575 52.419 17.5575 61.33 ;
      RECT 23.54 52.419 23.74 61.33 ;
      RECT 1.681 60.4585 1.739 61.454 ;
      RECT 1.909 60.4585 1.967 61.454 ;
      RECT 2.137 60.4585 2.195 61.454 ;
      RECT 2.365 60.4585 2.423 61.454 ;
      RECT 2.593 60.4585 2.651 61.454 ;
      RECT 2.821 60.4585 2.879 61.454 ;
      RECT 3.049 60.4585 3.107 61.454 ;
      RECT 3.277 60.4585 3.335 61.454 ;
      RECT 3.505 60.4585 3.563 61.454 ;
      RECT 3.733 60.4585 3.791 61.454 ;
      RECT 3.961 60.4585 4.019 61.454 ;
      RECT 4.189 60.4585 4.247 61.454 ;
      RECT 4.417 60.4585 4.475 61.454 ;
      RECT 4.645 60.4585 4.703 61.454 ;
      RECT 4.873 60.4585 4.931 61.454 ;
      RECT 5.101 60.4585 5.159 61.454 ;
      RECT 5.329 60.4585 5.387 61.454 ;
      RECT 5.557 60.4585 5.615 61.454 ;
      RECT 5.785 60.4585 5.843 61.454 ;
      RECT 6.013 60.4585 6.071 61.454 ;
      RECT 6.241 60.4585 6.299 61.454 ;
      RECT 6.469 60.4585 6.527 61.454 ;
      RECT 6.697 60.4585 6.755 61.454 ;
      RECT 6.925 60.4585 6.983 61.454 ;
      RECT 7.153 60.4585 7.211 61.454 ;
      RECT 7.381 60.4585 7.439 61.454 ;
      RECT 7.609 60.4585 7.667 61.454 ;
      RECT 7.837 60.4585 7.895 61.454 ;
      RECT 8.065 60.4585 8.123 61.454 ;
      RECT 8.293 60.4585 8.351 61.454 ;
      RECT 8.521 60.4585 8.579 61.454 ;
      RECT 8.749 60.4585 8.807 61.454 ;
      RECT 8.977 60.4585 9.035 61.454 ;
      RECT 9.205 60.4585 9.263 61.454 ;
      RECT 9.433 60.4585 9.491 61.454 ;
      RECT 9.661 60.4585 9.719 61.454 ;
      RECT 9.889 60.4585 9.947 61.454 ;
      RECT 10.117 60.4585 10.175 61.454 ;
      RECT 10.345 60.4585 10.403 61.454 ;
      RECT 10.573 60.4585 10.631 61.454 ;
      RECT 10.801 60.4585 10.859 61.454 ;
      RECT 11.029 60.4585 11.087 61.454 ;
      RECT 11.257 60.4585 11.315 61.454 ;
      RECT 11.485 60.4585 11.543 61.454 ;
      RECT 11.713 60.4585 11.771 61.454 ;
      RECT 11.941 60.4585 11.999 61.454 ;
      RECT 12.169 60.4585 12.227 61.454 ;
      RECT 12.397 60.4585 12.455 61.454 ;
      RECT 12.625 60.4585 12.683 61.454 ;
      RECT 12.853 60.4585 12.911 61.454 ;
      RECT 13.081 60.4585 13.139 61.454 ;
      RECT 13.309 60.4585 13.367 61.454 ;
      RECT 13.537 60.4585 13.595 61.454 ;
      RECT 13.765 60.4585 13.823 61.454 ;
      RECT 13.993 60.4585 14.051 61.454 ;
      RECT 14.221 60.4585 14.279 61.454 ;
      RECT 14.449 60.4585 14.507 61.454 ;
      RECT 14.677 60.4585 14.735 61.454 ;
      RECT 14.905 60.4585 14.963 61.454 ;
      RECT 15.133 60.4585 15.191 61.454 ;
      RECT 15.361 60.4585 15.419 61.454 ;
      RECT 15.589 60.4585 15.647 61.454 ;
      RECT 15.817 60.4585 15.875 61.454 ;
      RECT 16.045 60.4585 16.103 61.454 ;
      RECT 16.273 60.4585 16.331 61.454 ;
      RECT 16.501 60.4585 16.559 61.454 ;
      RECT 16.729 60.4585 16.787 61.454 ;
      RECT 18.781 60.4585 18.839 61.454 ;
      RECT 19.237 60.4585 19.295 61.454 ;
      RECT 19.465 60.4585 19.523 61.454 ;
      RECT 19.921 60.4585 19.979 61.454 ;
      RECT 21.061 60.4585 21.119 61.454 ;
      RECT 21.517 60.4585 21.575 61.454 ;
      RECT 21.745 60.4585 21.803 61.454 ;
      RECT 22.201 60.4585 22.259 61.454 ;
      RECT 24.253 60.4585 24.311 61.454 ;
      RECT 24.481 60.4585 24.539 61.454 ;
      RECT 24.709 60.4585 24.767 61.454 ;
      RECT 24.937 60.4585 24.995 61.454 ;
      RECT 25.165 60.4585 25.223 61.454 ;
      RECT 25.393 60.4585 25.451 61.454 ;
      RECT 25.621 60.4585 25.679 61.454 ;
      RECT 25.849 60.4585 25.907 61.454 ;
      RECT 26.077 60.4585 26.135 61.454 ;
      RECT 26.305 60.4585 26.363 61.454 ;
      RECT 26.533 60.4585 26.591 61.454 ;
      RECT 26.761 60.4585 26.819 61.454 ;
      RECT 26.989 60.4585 27.047 61.454 ;
      RECT 27.217 60.4585 27.275 61.454 ;
      RECT 27.445 60.4585 27.503 61.454 ;
      RECT 27.673 60.4585 27.731 61.454 ;
      RECT 27.901 60.4585 27.959 61.454 ;
      RECT 28.129 60.4585 28.187 61.454 ;
      RECT 28.357 60.4585 28.415 61.454 ;
      RECT 28.585 60.4585 28.643 61.454 ;
      RECT 28.813 60.4585 28.871 61.454 ;
      RECT 29.041 60.4585 29.099 61.454 ;
      RECT 29.269 60.4585 29.327 61.454 ;
      RECT 29.497 60.4585 29.555 61.454 ;
      RECT 29.725 60.4585 29.783 61.454 ;
      RECT 29.953 60.4585 30.011 61.454 ;
      RECT 30.181 60.4585 30.239 61.454 ;
      RECT 30.409 60.4585 30.467 61.454 ;
      RECT 30.637 60.4585 30.695 61.454 ;
      RECT 30.865 60.4585 30.923 61.454 ;
      RECT 31.093 60.4585 31.151 61.454 ;
      RECT 31.321 60.4585 31.379 61.454 ;
      RECT 31.549 60.4585 31.607 61.454 ;
      RECT 31.777 60.4585 31.835 61.454 ;
      RECT 32.005 60.4585 32.063 61.454 ;
      RECT 32.233 60.4585 32.291 61.454 ;
      RECT 32.461 60.4585 32.519 61.454 ;
      RECT 32.689 60.4585 32.747 61.454 ;
      RECT 32.917 60.4585 32.975 61.454 ;
      RECT 33.145 60.4585 33.203 61.454 ;
      RECT 33.373 60.4585 33.431 61.454 ;
      RECT 33.601 60.4585 33.659 61.454 ;
      RECT 33.829 60.4585 33.887 61.454 ;
      RECT 34.057 60.4585 34.115 61.454 ;
      RECT 34.285 60.4585 34.343 61.454 ;
      RECT 34.513 60.4585 34.571 61.454 ;
      RECT 34.741 60.4585 34.799 61.454 ;
      RECT 34.969 60.4585 35.027 61.454 ;
      RECT 35.197 60.4585 35.255 61.454 ;
      RECT 35.425 60.4585 35.483 61.454 ;
      RECT 35.653 60.4585 35.711 61.454 ;
      RECT 35.881 60.4585 35.939 61.454 ;
      RECT 36.109 60.4585 36.167 61.454 ;
      RECT 36.337 60.4585 36.395 61.454 ;
      RECT 36.565 60.4585 36.623 61.454 ;
      RECT 36.793 60.4585 36.851 61.454 ;
      RECT 37.021 60.4585 37.079 61.454 ;
      RECT 37.249 60.4585 37.307 61.454 ;
      RECT 37.477 60.4585 37.535 61.454 ;
      RECT 37.705 60.4585 37.763 61.454 ;
      RECT 37.933 60.4585 37.991 61.454 ;
      RECT 38.161 60.4585 38.219 61.454 ;
      RECT 38.389 60.4585 38.447 61.454 ;
      RECT 38.617 60.4585 38.675 61.454 ;
      RECT 38.845 60.4585 38.903 61.454 ;
      RECT 39.073 60.4585 39.131 61.454 ;
      RECT 39.301 60.4585 39.359 61.454 ;
      RECT 10.459 61.0815 10.517 62.309 ;
      RECT 30.523 61.0815 30.581 62.309 ;
      RECT 18.667 61.356 18.725 62.3085 ;
      RECT 18.895 61.356 18.953 62.3085 ;
      RECT 19.351 61.356 19.409 62.3085 ;
      RECT 19.579 61.356 19.637 62.3085 ;
      RECT 19.807 61.356 19.865 62.3085 ;
      RECT 21.175 61.356 21.233 62.3085 ;
      RECT 21.403 61.356 21.461 62.3085 ;
      RECT 21.631 61.356 21.689 62.3085 ;
      RECT 22.087 61.356 22.145 62.3085 ;
      RECT 22.315 61.356 22.373 62.3085 ;
      RECT 4.759 61.3585 4.817 62.309 ;
      RECT 4.987 61.3585 5.045 62.309 ;
      RECT 5.215 61.3585 5.273 62.309 ;
      RECT 5.443 61.3585 5.501 62.309 ;
      RECT 5.671 61.3585 5.729 62.309 ;
      RECT 5.899 61.3585 5.957 62.309 ;
      RECT 6.127 61.3585 6.185 62.309 ;
      RECT 6.355 61.3585 6.413 62.309 ;
      RECT 6.583 61.3585 6.641 62.309 ;
      RECT 6.811 61.3585 6.869 62.309 ;
      RECT 7.039 61.3585 7.097 62.309 ;
      RECT 7.267 61.3585 7.325 62.309 ;
      RECT 7.495 61.3585 7.553 62.309 ;
      RECT 7.723 61.3585 7.781 62.309 ;
      RECT 7.951 61.3585 8.009 62.309 ;
      RECT 8.179 61.3585 8.237 62.309 ;
      RECT 8.407 61.3585 8.465 62.309 ;
      RECT 8.635 61.3585 8.693 62.309 ;
      RECT 8.863 61.3585 8.921 62.309 ;
      RECT 9.091 61.3585 9.149 62.309 ;
      RECT 9.319 61.3585 9.377 62.309 ;
      RECT 9.547 61.3585 9.605 62.309 ;
      RECT 9.775 61.3585 9.833 62.309 ;
      RECT 10.231 61.3585 10.289 62.309 ;
      RECT 10.687 61.3585 10.745 62.309 ;
      RECT 10.915 61.3585 10.973 62.309 ;
      RECT 11.143 61.3585 11.201 62.309 ;
      RECT 11.371 61.3585 11.429 62.309 ;
      RECT 11.599 61.3585 11.657 62.309 ;
      RECT 11.827 61.3585 11.885 62.309 ;
      RECT 12.055 61.3585 12.113 62.309 ;
      RECT 12.283 61.3585 12.341 62.309 ;
      RECT 12.511 61.3585 12.569 62.309 ;
      RECT 12.739 61.3585 12.797 62.309 ;
      RECT 12.967 61.3585 13.025 62.309 ;
      RECT 13.195 61.3585 13.253 62.309 ;
      RECT 13.423 61.3585 13.481 62.309 ;
      RECT 13.651 61.3585 13.709 62.309 ;
      RECT 13.879 61.3585 13.937 62.309 ;
      RECT 14.107 61.3585 14.165 62.309 ;
      RECT 14.335 61.3585 14.393 62.309 ;
      RECT 14.563 61.3585 14.621 62.309 ;
      RECT 14.791 61.3585 14.849 62.309 ;
      RECT 15.019 61.3585 15.077 62.309 ;
      RECT 15.247 61.3585 15.305 62.309 ;
      RECT 15.475 61.3585 15.533 62.309 ;
      RECT 15.703 61.3585 15.761 62.309 ;
      RECT 15.931 61.3585 15.989 62.309 ;
      RECT 16.159 61.3585 16.217 62.309 ;
      RECT 16.387 61.3585 16.445 62.309 ;
      RECT 16.615 61.3585 16.673 62.309 ;
      RECT 16.843 61.3585 16.901 62.309 ;
      RECT 24.139 61.3585 24.197 62.309 ;
      RECT 24.367 61.3585 24.425 62.309 ;
      RECT 24.595 61.3585 24.653 62.309 ;
      RECT 24.823 61.3585 24.881 62.309 ;
      RECT 25.051 61.3585 25.109 62.309 ;
      RECT 25.279 61.3585 25.337 62.309 ;
      RECT 25.507 61.3585 25.565 62.309 ;
      RECT 25.735 61.3585 25.793 62.309 ;
      RECT 25.963 61.3585 26.021 62.309 ;
      RECT 26.191 61.3585 26.249 62.309 ;
      RECT 26.419 61.3585 26.477 62.309 ;
      RECT 26.647 61.3585 26.705 62.309 ;
      RECT 26.875 61.3585 26.933 62.309 ;
      RECT 27.103 61.3585 27.161 62.309 ;
      RECT 27.331 61.3585 27.389 62.309 ;
      RECT 27.559 61.3585 27.617 62.309 ;
      RECT 27.787 61.3585 27.845 62.309 ;
      RECT 28.015 61.3585 28.073 62.309 ;
      RECT 28.243 61.3585 28.301 62.309 ;
      RECT 28.471 61.3585 28.529 62.309 ;
      RECT 28.699 61.3585 28.757 62.309 ;
      RECT 28.927 61.3585 28.985 62.309 ;
      RECT 29.155 61.3585 29.213 62.309 ;
      RECT 29.383 61.3585 29.441 62.309 ;
      RECT 29.611 61.3585 29.669 62.309 ;
      RECT 29.839 61.3585 29.897 62.309 ;
      RECT 30.067 61.3585 30.125 62.309 ;
      RECT 30.295 61.3585 30.353 62.309 ;
      RECT 30.751 61.3585 30.809 62.309 ;
      RECT 31.207 61.3585 31.265 62.309 ;
      RECT 31.435 61.3585 31.493 62.309 ;
      RECT 31.663 61.3585 31.721 62.309 ;
      RECT 31.891 61.3585 31.949 62.309 ;
      RECT 32.119 61.3585 32.177 62.309 ;
      RECT 32.347 61.3585 32.405 62.309 ;
      RECT 32.575 61.3585 32.633 62.309 ;
      RECT 32.803 61.3585 32.861 62.309 ;
      RECT 33.031 61.3585 33.089 62.309 ;
      RECT 33.259 61.3585 33.317 62.309 ;
      RECT 33.487 61.3585 33.545 62.309 ;
      RECT 33.715 61.3585 33.773 62.309 ;
      RECT 33.943 61.3585 34.001 62.309 ;
      RECT 34.171 61.3585 34.229 62.309 ;
      RECT 34.399 61.3585 34.457 62.309 ;
      RECT 34.627 61.3585 34.685 62.309 ;
      RECT 34.855 61.3585 34.913 62.309 ;
      RECT 35.083 61.3585 35.141 62.309 ;
      RECT 35.311 61.3585 35.369 62.309 ;
      RECT 35.539 61.3585 35.597 62.309 ;
      RECT 35.767 61.3585 35.825 62.309 ;
      RECT 35.995 61.3585 36.053 62.309 ;
      RECT 36.223 61.3585 36.281 62.309 ;
      RECT 1.681 61.556 1.739 62.9715 ;
      RECT 1.909 61.556 1.967 62.9715 ;
      RECT 2.137 61.556 2.195 62.9715 ;
      RECT 2.365 61.556 2.423 62.9715 ;
      RECT 2.593 61.556 2.651 62.9715 ;
      RECT 2.821 61.556 2.879 62.9715 ;
      RECT 3.049 61.556 3.107 62.9715 ;
      RECT 3.277 61.556 3.335 62.9715 ;
      RECT 3.505 61.556 3.563 62.9715 ;
      RECT 3.733 61.556 3.791 62.9715 ;
      RECT 3.961 61.556 4.019 62.9715 ;
      RECT 37.021 61.556 37.079 62.9715 ;
      RECT 37.249 61.556 37.307 62.9715 ;
      RECT 37.477 61.556 37.535 62.9715 ;
      RECT 37.705 61.556 37.763 62.9715 ;
      RECT 37.933 61.556 37.991 62.9715 ;
      RECT 38.161 61.556 38.219 62.9715 ;
      RECT 38.389 61.556 38.447 62.9715 ;
      RECT 38.617 61.556 38.675 62.9715 ;
      RECT 38.845 61.556 38.903 62.9715 ;
      RECT 39.073 61.556 39.131 62.9715 ;
      RECT 39.301 61.556 39.359 62.9715 ;
      RECT 16.843 62.5435 16.901 65.334 ;
      RECT 17.071 62.5435 17.129 65.334 ;
      RECT 17.299 62.5435 17.357 65.334 ;
      RECT 23.683 62.5435 23.741 65.334 ;
      RECT 23.911 62.5435 23.969 65.334 ;
      RECT 24.139 62.5435 24.197 65.334 ;
      RECT 13.537 63.3535 13.595 65.334 ;
      RECT 13.765 63.3535 13.823 65.334 ;
      RECT 13.993 63.3535 14.051 65.334 ;
      RECT 14.221 63.3535 14.279 65.334 ;
      RECT 14.449 63.3535 14.507 65.334 ;
      RECT 14.677 63.3535 14.735 65.334 ;
      RECT 14.905 63.3535 14.963 65.334 ;
      RECT 15.133 63.3535 15.191 65.334 ;
      RECT 15.361 63.3535 15.419 65.334 ;
      RECT 15.589 63.3535 15.647 65.334 ;
      RECT 15.817 63.3535 15.875 65.334 ;
      RECT 16.045 63.3535 16.103 65.334 ;
      RECT 16.273 63.3535 16.331 65.334 ;
      RECT 24.709 63.3535 24.767 65.334 ;
      RECT 24.937 63.3535 24.995 65.334 ;
      RECT 25.165 63.3535 25.223 65.334 ;
      RECT 25.393 63.3535 25.451 65.334 ;
      RECT 25.621 63.3535 25.679 65.334 ;
      RECT 25.849 63.3535 25.907 65.334 ;
      RECT 26.077 63.3535 26.135 65.334 ;
      RECT 26.305 63.3535 26.363 65.334 ;
      RECT 26.533 63.3535 26.591 65.334 ;
      RECT 26.761 63.3535 26.819 65.334 ;
      RECT 26.989 63.3535 27.047 65.334 ;
      RECT 27.217 63.3535 27.275 65.334 ;
      RECT 27.445 63.3535 27.503 65.334 ;
    LAYER M0 ;
      RECT MASK 1 0 0 41.04 90 ;
      RECT MASK 2 0 0 41.04 90 ;
    LAYER LUP_015U ;
      RECT 1.5635 43.661 17.3605 43.729 ;
      RECT 23.6795 43.661 39.4765 43.729 ;
      RECT 1.5635 45.221 17.3605 45.289 ;
      RECT 23.6795 45.221 39.4765 45.289 ;
      RECT 1.5635 57.851 17.3605 57.919 ;
      RECT 23.6795 57.851 39.4765 57.919 ;
      RECT 1.5635 59.411 17.3605 59.479 ;
      RECT 23.6795 59.411 39.4765 59.479 ;
      RECT 3.944 66.33 37.096 89.49 ;
  END
END dwc_ddrphy_se_io_ns

END LIBRARY
