# LEF OUT API 
# Creation Date : Tue Apr 16 16:13:30 IST 2019
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_vrefdacref
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_vrefdacref 0 0 ;
  SYMMETRY X Y ;
  SIZE 41.04 BY 90 ;
  PIN VDD2H
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.3 70.875 40.74 71.325 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 18.27 40.74 18.77 ;
        RECT 0.3 8.27 40.74 8.77 ;
        RECT 0.3 88.875 40.74 89.325 ;
        RECT 0.3 78.075 40.74 78.525 ;
        RECT 0.3 76.275 40.74 76.725 ;
        RECT 0.3 74.475 40.74 74.925 ;
        RECT 0.3 72.675 40.74 73.125 ;
        RECT 0.3 67.275 40.74 67.725 ;
        RECT 0.3 56.27 40.74 56.77 ;
        RECT 0.3 54.27 40.74 54.77 ;
        RECT 0.3 52.27 40.74 52.77 ;
        RECT 0.3 47.27 40.74 47.77 ;
        RECT 0.3 45.27 40.74 45.77 ;
        RECT 0.3 24.27 40.74 24.77 ;
        RECT 0.3 22.27 40.74 22.77 ;
        RECT 0.3 16.27 40.74 16.77 ;
        RECT 0.3 12.27 40.74 12.77 ;
        RECT 0.3 10.27 40.74 10.77 ;
        RECT 0.3 6.27 40.74 6.77 ;
        RECT 0.3 2.27 40.74 2.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 69.075 40.74 69.525 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 49.27 40.74 49.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 14.27 40.74 14.77 ;
    END
  END VDD2H
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M6 ;
        RECT 0.3 65.27 40.74 65.77 ;
        RECT 0.3 64.27 40.74 64.77 ;
        RECT 0.3 63.27 40.74 63.77 ;
        RECT 0.3 62.27 40.74 62.77 ;
        RECT 0.3 61.27 40.74 61.77 ;
        RECT 0.3 59.27 40.74 59.77 ;
        RECT 0.3 58.27 40.74 58.77 ;
        RECT 0.3 57.27 40.74 57.77 ;
        RECT 0.3 55.27 40.74 55.77 ;
        RECT 0.3 53.27 40.74 53.77 ;
        RECT 0.3 51.27 40.74 51.77 ;
        RECT 0.3 50.27 40.74 50.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 87.975 40.74 88.425 ;
        RECT 0.3 86.175 40.74 86.625 ;
        RECT 0.3 84.375 40.74 84.825 ;
        RECT 0.3 82.575 40.74 83.025 ;
        RECT 0.3 80.775 40.74 81.225 ;
        RECT 0.3 78.975 40.74 79.425 ;
        RECT 0.3 77.175 40.74 77.625 ;
        RECT 0.3 66.375 40.74 66.825 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 48.27 40.74 48.77 ;
        RECT 0.3 46.27 40.74 46.77 ;
        RECT 0.3 33.77 40.74 34.27 ;
        RECT 0.3 5.27 40.74 5.77 ;
        RECT 0.3 3.27 40.74 3.77 ;
        RECT 0.3 1.27 40.74 1.77 ;
    END
  END VSS
  PIN AOBS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.22 LAYER M6 ;
    ANTENNADIFFAREA 0 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 11.0233 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 5.601 79.875 35.439 80.325 ;
    END
    PORT
      LAYER M6 ;
        RECT 5.601 87.075 35.439 87.525 ;
        RECT 5.601 85.275 35.439 85.725 ;
        RECT 5.601 83.475 35.439 83.925 ;
        RECT 5.601 81.675 35.439 82.125 ;
        RECT 5.6 75.375 35.44 75.825 ;
        RECT 5.6 73.575 35.44 74.025 ;
        RECT 5.6 71.775 35.44 72.225 ;
        RECT 5.6 69.975 35.44 70.425 ;
        RECT 5.6 68.175 35.44 68.625 ;
        RECT 0.3 60.27 40.74 60.77 ;
    END
  END AOBS
  PIN AObsIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.5343 LAYER M5 ;
    ANTENNADIFFAREA 77.4158 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 23.992 0 24.192 0.2 ;
    END
  END AObsIn
  PIN VrefDacRef
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 121.32 LAYER M6 ;
    ANTENNADIFFAREA 109.533 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 0 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0.3 17.27 40.74 17.77 ;
        RECT 0.3 43.27 40.74 43.77 ;
        RECT 0.3 41.27 40.74 41.77 ;
        RECT 0.3 39.27 40.74 39.77 ;
        RECT 0.3 37.27 40.74 37.77 ;
        RECT 0.3 31.27 40.74 31.77 ;
        RECT 0.3 26.27 40.74 26.77 ;
        RECT 0.3 23.27 40.74 23.77 ;
        RECT 0.3 15.27 40.74 15.77 ;
        RECT 0.3 13.27 40.74 13.77 ;
        RECT 0.3 11.27 40.74 11.77 ;
        RECT 0.3 9.27 40.74 9.77 ;
        RECT 0.3 7.27 40.74 7.77 ;
    END
  END VrefDacRef
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.3 0.27 40.74 0.77 ;
    END
  END VDD
  PIN InAObsEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.150252 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0872 LAYER M5 ;
      ANTENNAMAXAREACAR 5.90346 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 26.562 0 26.638 0.114 ;
    END
  END InAObsEn
  PIN PwrOkVDD2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.22 LAYER M6 ;
    ANTENNADIFFAREA 0.012032 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.288128 LAYER M6 ;
      ANTENNAMAXAREACAR 89.8455 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0.3 4.27 40.74 4.77 ;
    END
  END PwrOkVDD2
  PIN PowerDown
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.150252 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0872 LAYER M5 ;
      ANTENNAMAXAREACAR 4.01355 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 25.726 0 25.802 0.114 ;
    END
  END PowerDown
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.3 44.27 40.74 44.77 ;
        RECT 0.3 42.27 40.74 42.77 ;
        RECT 0.3 40.27 40.74 40.77 ;
        RECT 0.3 38.27 40.74 38.77 ;
        RECT 0.3 36.27 40.74 36.77 ;
        RECT 0.3 34.77 40.74 35.27 ;
        RECT 0.3 27.77 40.74 28.27 ;
        RECT 0.3 25.27 40.74 25.77 ;
    END
  END VDDQ
  PIN DacRefModeCtl
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136002 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0872 LAYER M5 ;
      ANTENNAMAXAREACAR 3.58615 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 4.142 0 4.218 0.114 ;
    END
  END DacRefModeCtl
  OBS
    LAYER M1 ;
      RECT MASK 1 0 0 41.04 90 ;
    LAYER M1 ;
      RECT MASK 2 0 0 41.04 90 ;
    LAYER M2 ;
      RECT MASK 1 0 0 41.04 90 ;
    LAYER M2 ;
      RECT MASK 2 0 0 41.04 90 ;
    LAYER M3 ;
      RECT MASK 1 0 0 41.04 90 ;
    LAYER M4 ;
      RECT 0 0 41.04 90 ;
    LAYER M3 ;
      RECT MASK 2 0 0 41.04 90 ;
    LAYER M4 ;
      RECT 14.4095 1.82 15.1555 1.9 ;
      RECT 25.477 1.82 26.026 1.9 ;
      RECT 26.485 1.82 29.094 1.9 ;
      RECT 39.4355 1.82 39.957 1.9 ;
      RECT 8.3815 3.43 39.5215 3.65 ;
      RECT 8.3815 3.85 39.5215 4.07 ;
      RECT 3.2985 4.1965 4.6555 4.2565 ;
      RECT 8.847 4.2935 20.0865 4.3735 ;
      RECT 20.8105 4.2935 29.1145 4.3735 ;
      RECT 3.2985 4.3165 4.6555 4.3765 ;
      RECT 3.2985 4.4365 4.6555 4.4965 ;
      RECT 13.276 4.4535 23.5225 4.5335 ;
      RECT 25.5655 4.4535 36.811 4.5335 ;
      RECT 17.502 4.6135 23.554 4.6935 ;
      RECT 29.5595 4.6135 38.376 4.6935 ;
      RECT 3.2985 4.6765 4.6555 4.7365 ;
      RECT 3.2985 4.7965 4.6555 4.8565 ;
      RECT 3.2985 4.9165 4.6555 4.9765 ;
      RECT 8.3815 4.94 39.0755 5.14 ;
      RECT 18.3585 5.698 27.425 5.778 ;
      RECT 18.3585 5.858 28.7215 5.938 ;
      RECT 29.576 5.858 38.399 5.938 ;
      RECT 1.63 6.24 39.421 6.36 ;
      RECT 2.011 6.9185 39.029 6.9785 ;
      RECT 2.011 7.1585 39.029 7.2185 ;
      RECT 2.011 7.8485 39.029 7.9085 ;
      RECT 2.011 8.0885 39.029 8.1485 ;
      RECT 2.011 8.7785 39.029 8.8385 ;
      RECT 2.011 9.0185 39.029 9.0785 ;
      RECT 2.011 9.7085 39.029 9.7685 ;
      RECT 2.011 9.9485 39.029 10.0085 ;
      RECT 2.011 10.6385 39.029 10.6985 ;
      RECT 2.011 10.8785 39.029 10.9385 ;
      RECT 2.011 11.5685 39.029 11.6285 ;
      RECT 2.011 11.8085 39.029 11.8685 ;
      RECT 2.011 12.4985 39.029 12.5585 ;
      RECT 2.011 12.7385 39.029 12.7985 ;
      RECT 2.011 13.4285 39.029 13.4885 ;
      RECT 2.011 13.6685 39.029 13.7285 ;
      RECT 2.011 14.3585 39.029 14.4185 ;
      RECT 2.011 14.5985 39.029 14.6585 ;
      RECT 1.63 15.24 39.421 15.36 ;
      RECT 1.63 15.87 39.3855 15.99 ;
      RECT 2.011 16.5485 39.029 16.6085 ;
      RECT 2.011 16.7885 39.029 16.8485 ;
      RECT 2.011 17.4785 39.029 17.5385 ;
      RECT 2.011 17.7185 39.029 17.7785 ;
      RECT 2.011 18.4085 39.029 18.4685 ;
      RECT 2.011 18.6485 39.029 18.7085 ;
      RECT 2.011 19.3385 39.029 19.3985 ;
      RECT 2.011 19.5785 39.029 19.6385 ;
      RECT 2.011 20.2685 39.029 20.3285 ;
      RECT 2.011 20.5085 39.029 20.5685 ;
      RECT 2.011 21.1985 39.029 21.2585 ;
      RECT 2.011 21.4385 39.029 21.4985 ;
      RECT 2.011 22.1285 39.029 22.1885 ;
      RECT 2.011 22.3685 39.029 22.4285 ;
      RECT 2.011 23.0585 39.029 23.1185 ;
      RECT 2.011 23.2985 39.029 23.3585 ;
      RECT 2.011 23.9885 39.029 24.0485 ;
      RECT 2.011 24.2285 39.029 24.2885 ;
      RECT 1.63 24.87 39.3855 24.99 ;
      RECT 24.7245 25.25 36.354 25.33 ;
      RECT 1.63 25.59 39.421 25.71 ;
      RECT 2.011 26.2685 39.029 26.3285 ;
      RECT 2.011 26.5085 39.029 26.5685 ;
      RECT 2.011 27.1985 39.029 27.2585 ;
      RECT 2.011 27.4385 39.029 27.4985 ;
      RECT 2.011 28.1285 39.029 28.1885 ;
      RECT 2.011 28.3685 39.029 28.4285 ;
      RECT 2.011 29.0585 39.029 29.1185 ;
      RECT 2.011 29.2985 39.029 29.3585 ;
      RECT 2.011 29.9885 39.029 30.0485 ;
      RECT 2.011 30.2285 39.029 30.2885 ;
      RECT 2.011 30.9185 39.029 30.9785 ;
      RECT 2.011 31.1585 39.029 31.2185 ;
      RECT 2.011 31.8485 39.029 31.9085 ;
      RECT 2.011 32.0885 39.029 32.1485 ;
      RECT 2.011 32.7785 39.029 32.8385 ;
      RECT 2.011 33.0185 39.029 33.0785 ;
      RECT 2.011 33.7085 39.029 33.7685 ;
      RECT 2.011 33.9485 39.029 34.0085 ;
      RECT 1.63 34.59 39.9665 34.71 ;
      RECT 1.63 35.22 39.3855 35.34 ;
      RECT 2.011 35.8985 39.029 35.9585 ;
      RECT 2.011 36.1385 39.029 36.1985 ;
      RECT 2.011 36.8285 39.029 36.8885 ;
      RECT 2.011 37.0685 39.029 37.1285 ;
      RECT 2.011 37.7585 39.029 37.8185 ;
      RECT 2.011 37.9985 39.029 38.0585 ;
      RECT 2.011 38.6885 39.029 38.7485 ;
      RECT 2.011 38.9285 39.029 38.9885 ;
      RECT 2.011 39.6185 39.029 39.6785 ;
      RECT 2.011 39.8585 39.029 39.9185 ;
      RECT 2.011 40.5485 39.029 40.6085 ;
      RECT 2.011 40.7885 39.029 40.8485 ;
      RECT 2.011 41.4785 39.029 41.5385 ;
      RECT 2.011 41.7185 39.029 41.7785 ;
      RECT 2.011 42.4085 39.029 42.4685 ;
      RECT 2.011 42.6485 39.029 42.7085 ;
      RECT 2.011 43.3385 39.029 43.3985 ;
      RECT 2.011 43.5785 39.029 43.6385 ;
      RECT 1.63 44.22 39.3855 44.34 ;
      RECT 9.213 44.756 9.489 44.836 ;
      RECT 9.213 44.916 9.489 44.996 ;
      RECT 8.0105 47.16 40.4615 47.28 ;
      RECT 8.6475 47.7 39.764 47.82 ;
      RECT 9.0295 48.3785 39.4075 48.4385 ;
      RECT 9.0295 48.6185 39.4075 48.6785 ;
      RECT 9.198 48.8905 39.3435 48.9705 ;
      RECT 9.0295 49.3085 39.4075 49.3685 ;
      RECT 9.0295 49.5485 39.4075 49.6085 ;
      RECT 9.198 49.8205 39.3435 49.9005 ;
      RECT 9.0295 50.2385 39.4075 50.2985 ;
      RECT 9.0295 50.4785 39.4075 50.5385 ;
      RECT 9.198 50.7505 39.3435 50.8305 ;
      RECT 9.0295 51.1685 39.4075 51.2285 ;
      RECT 9.0295 51.4085 39.4075 51.4685 ;
      RECT 9.198 51.6805 39.3435 51.7605 ;
      RECT 9.0295 52.0985 39.4075 52.1585 ;
      RECT 9.0295 52.3385 39.4075 52.3985 ;
      RECT 9.198 52.6105 39.3435 52.6905 ;
      RECT 9.0295 53.0285 39.4075 53.0885 ;
      RECT 9.0295 53.2685 39.4075 53.3285 ;
      RECT 9.198 53.5405 39.3435 53.6205 ;
      RECT 1.1965 53.638 6.7125 54.063 ;
      RECT 9.0295 53.9585 39.4075 54.0185 ;
      RECT 9.0295 54.1985 39.4075 54.2585 ;
      RECT 9.198 54.4705 39.3435 54.5505 ;
      RECT 8.6475 54.84 39.764 54.96 ;
      RECT 8.0105 55.38 40.4865 55.5 ;
      RECT 7.164 55.765 38.782 56.165 ;
      RECT 1.1965 55.978 6.7125 56.403 ;
      RECT 8.0105 56.43 40.4615 56.55 ;
      RECT 8.6475 56.97 39.764 57.09 ;
      RECT 8.695 57.6485 39.742 57.7085 ;
      RECT 8.695 57.8885 39.742 57.9485 ;
      RECT 9.268 58.1605 39.5035 58.2405 ;
      RECT 1.0465 58.439 6.8625 58.83 ;
      RECT 8.695 58.5785 39.742 58.6385 ;
      RECT 8.695 58.8185 39.742 58.8785 ;
      RECT 9.268 59.0905 39.5035 59.1705 ;
      RECT 8.695 59.5085 39.742 59.5685 ;
      RECT 8.695 59.7485 39.742 59.8085 ;
      RECT 9.268 60.0205 39.5035 60.1005 ;
      RECT 1.0465 60.268 6.8625 60.654 ;
      RECT 8.695 60.4385 39.742 60.4985 ;
      RECT 8.695 60.6785 39.742 60.7385 ;
      RECT 9.268 60.9505 39.5035 61.0305 ;
      RECT 8.695 61.3685 39.742 61.4285 ;
      RECT 8.695 61.6085 39.742 61.6685 ;
      RECT 9.268 61.8805 39.5035 61.9605 ;
      RECT 8.695 62.2985 39.742 62.3585 ;
      RECT 8.695 62.5385 39.742 62.5985 ;
      RECT 9.268 62.8105 39.5035 62.8905 ;
      RECT 8.695 63.2285 39.742 63.2885 ;
      RECT 8.695 63.4685 39.742 63.5285 ;
      RECT 9.268 63.7405 39.5035 63.8205 ;
      RECT 8.6475 64.1095 39.764 64.2295 ;
      RECT 8.0105 64.65 40.4865 64.77 ;
      RECT 0.3 66.43 40.74 66.79 ;
      RECT 5.6 68.15 35.44 68.65 ;
      RECT 0.3 69.05 40.74 69.55 ;
      RECT 5.6 69.95 35.44 70.45 ;
      RECT 0.3 70.85 40.74 71.35 ;
      RECT 5.6 71.75 35.44 72.25 ;
      RECT 0.3 72.65 40.74 73.15 ;
      RECT 5.6 73.55 35.44 74.05 ;
      RECT 0.3 74.45 40.74 74.95 ;
      RECT 5.6 75.35 35.44 75.85 ;
      RECT 0.3 76.25 40.74 76.75 ;
      RECT 0.3 77.21 40.74 77.57 ;
      RECT 0.3 78.13 40.74 78.49 ;
      RECT 0.3 78.95 40.74 79.45 ;
      RECT 5.601 79.85 35.439 80.35 ;
      RECT 0.3 80.75 40.74 81.25 ;
      RECT 5.601 81.65 35.439 82.15 ;
      RECT 0.3 82.55 40.74 83.05 ;
      RECT 5.601 83.45 35.439 83.95 ;
      RECT 0.3 84.35 40.74 84.85 ;
      RECT 5.601 85.25 35.439 85.75 ;
      RECT 0.3 86.15 40.74 86.65 ;
      RECT 5.601 87.05 35.439 87.55 ;
      RECT 4.141 88.91 36.899 89.27 ;
    LAYER M5 ;
      POLYGON 4.066 0 4.066 0.19 4.294 0.19 4.294 0 23.916 0 23.916 0.276 24.268 0.276 24.268 0 25.65 0 25.65 0.19 25.878 0.19 25.878 0 26.486 0 26.486 0.19 26.714 0.19 26.714 0 41.04 0 41.04 90 0 90 0 0 ;
    LAYER M4 ;
      RECT 2.141 0.8 39.5055 1 ;
      RECT 2.1405 1.16 39.504 1.36 ;
      RECT 3.8985 1.66 4.336 1.74 ;
      RECT 17.7715 1.66 39.2425 1.74 ;
      RECT 2.4135 2.13 4.89 2.31 ;
      RECT 5.2375 2.13 8.7305 2.31 ;
      RECT 9.4445 2.13 20.3295 2.31 ;
      RECT 20.7845 2.13 24.5055 2.31 ;
      RECT 25.0145 2.13 29.7645 2.31 ;
      RECT 30.3755 2.13 34.14 2.31 ;
      RECT 34.4375 2.13 39.125 2.31 ;
      RECT 2.414 2.49 4.89 2.67 ;
      RECT 5.2375 2.49 8.732 2.67 ;
      RECT 9.445 2.49 20.331 2.67 ;
      RECT 20.785 2.49 24.507 2.67 ;
      RECT 25.015 2.49 29.766 2.67 ;
      RECT 30.376 2.49 34.1415 2.67 ;
      RECT 34.4375 2.49 39.125 2.67 ;
      RECT 3.794 4.5565 4.6555 4.6165 ;
      RECT 8.3815 5.37 39.0755 5.55 ;
      RECT 2.011 6.7985 39.0985 6.8585 ;
      RECT 2.011 7.0385 39.0985 7.0985 ;
      RECT 2.1645 7.4305 38.8905 7.5105 ;
      RECT 2.011 7.7285 39.0985 7.7885 ;
      RECT 2.011 7.9685 39.0985 8.0285 ;
      RECT 2.1645 8.3605 38.8905 8.4405 ;
      RECT 2.011 8.6585 39.0985 8.7185 ;
      RECT 2.011 8.8985 39.0985 8.9585 ;
      RECT 2.1645 9.2905 38.8905 9.3705 ;
      RECT 2.011 9.5885 39.0985 9.6485 ;
      RECT 2.011 9.8285 39.0985 9.8885 ;
      RECT 2.1645 10.2205 38.8905 10.3005 ;
      RECT 2.011 10.5185 39.0985 10.5785 ;
      RECT 2.011 10.7585 39.0985 10.8185 ;
      RECT 2.1645 11.1505 38.8905 11.2305 ;
      RECT 2.011 11.4485 39.0985 11.5085 ;
      RECT 2.011 11.6885 39.0985 11.7485 ;
      RECT 2.1645 12.0805 38.8905 12.1605 ;
      RECT 2.011 12.3785 39.0985 12.4385 ;
      RECT 2.011 12.6185 39.0985 12.6785 ;
      RECT 2.1645 13.0105 38.8905 13.0905 ;
      RECT 2.011 13.3085 39.0985 13.3685 ;
      RECT 2.011 13.5485 39.0985 13.6085 ;
      RECT 2.1645 13.9405 38.8905 14.0205 ;
      RECT 2.011 14.2385 39.0985 14.2985 ;
      RECT 2.011 14.4785 39.0985 14.5385 ;
      RECT 2.1645 14.8705 38.8905 14.9505 ;
      RECT 2.011 16.4285 39.0985 16.4885 ;
      RECT 2.011 16.6685 39.0985 16.7285 ;
      RECT 2.1645 17.0605 38.8905 17.1405 ;
      RECT 2.011 17.3585 39.0985 17.4185 ;
      RECT 2.011 17.5985 39.0985 17.6585 ;
      RECT 2.1645 17.9905 38.8905 18.0705 ;
      RECT 2.011 18.2885 39.0985 18.3485 ;
      RECT 2.011 18.5285 39.0985 18.5885 ;
      RECT 2.1645 18.9205 38.8905 19.0005 ;
      RECT 2.011 19.2185 39.0985 19.2785 ;
      RECT 2.011 19.4585 39.0985 19.5185 ;
      RECT 2.1645 19.8505 38.8905 19.9305 ;
      RECT 2.011 20.1485 39.0985 20.2085 ;
      RECT 2.011 20.3885 39.0985 20.4485 ;
      RECT 2.1645 20.7805 38.8905 20.8605 ;
      RECT 2.011 21.0785 39.0985 21.1385 ;
      RECT 2.011 21.3185 39.0985 21.3785 ;
      RECT 2.1645 21.7105 38.8905 21.7905 ;
      RECT 2.011 22.0085 39.0985 22.0685 ;
      RECT 2.011 22.2485 39.0985 22.3085 ;
      RECT 2.1645 22.6405 38.8905 22.7205 ;
      RECT 2.011 22.9385 39.0985 22.9985 ;
      RECT 2.011 23.1785 39.0985 23.2385 ;
      RECT 2.1645 23.5705 38.8905 23.6505 ;
      RECT 2.011 23.8685 39.0985 23.9285 ;
      RECT 2.011 24.1085 39.0985 24.1685 ;
      RECT 2.1645 24.5005 38.8905 24.5805 ;
      RECT 2.011 26.1485 39.0985 26.2085 ;
      RECT 2.011 26.3885 39.0985 26.4485 ;
      RECT 2.1645 26.7805 38.8905 26.8605 ;
      RECT 2.011 27.0785 39.0985 27.1385 ;
      RECT 2.011 27.3185 39.0985 27.3785 ;
      RECT 2.1645 27.7105 38.8905 27.7905 ;
      RECT 2.011 28.0085 39.0985 28.0685 ;
      RECT 2.011 28.2485 39.0985 28.3085 ;
      RECT 2.1645 28.6405 38.8905 28.7205 ;
      RECT 2.011 28.9385 39.0985 28.9985 ;
      RECT 2.011 29.1785 39.0985 29.2385 ;
      RECT 2.1645 29.5705 38.8905 29.6505 ;
      RECT 2.011 29.8685 39.0985 29.9285 ;
      RECT 2.011 30.1085 39.0985 30.1685 ;
      RECT 2.1645 30.5005 38.8905 30.5805 ;
      RECT 2.011 30.7985 39.0985 30.8585 ;
      RECT 2.011 31.0385 39.0985 31.0985 ;
      RECT 2.1645 31.4305 38.8905 31.5105 ;
      RECT 2.011 31.7285 39.0985 31.7885 ;
      RECT 2.011 31.9685 39.0985 32.0285 ;
      RECT 2.1645 32.3605 38.8905 32.4405 ;
      RECT 2.011 32.6585 39.0985 32.7185 ;
      RECT 2.011 32.8985 39.0985 32.9585 ;
      RECT 2.1645 33.2905 38.8905 33.3705 ;
      RECT 2.011 33.5885 39.0985 33.6485 ;
      RECT 2.011 33.8285 39.0985 33.8885 ;
      RECT 2.1645 34.2205 38.8905 34.3005 ;
      RECT 2.5005 34.9065 38.1285 34.9865 ;
      RECT 2.011 35.7785 39.0985 35.8385 ;
      RECT 2.011 36.0185 39.0985 36.0785 ;
      RECT 2.1645 36.4105 38.8905 36.4905 ;
      RECT 2.011 36.7085 39.0985 36.7685 ;
      RECT 2.011 36.9485 39.0985 37.0085 ;
      RECT 2.1645 37.3405 38.8905 37.4205 ;
      RECT 2.011 37.6385 39.0985 37.6985 ;
      RECT 2.011 37.8785 39.0985 37.9385 ;
      RECT 2.1645 38.2705 38.8905 38.3505 ;
      RECT 2.011 38.5685 39.0985 38.6285 ;
      RECT 2.011 38.8085 39.0985 38.8685 ;
      RECT 2.1645 39.2005 38.8905 39.2805 ;
      RECT 2.011 39.4985 39.0985 39.5585 ;
      RECT 2.011 39.7385 39.0985 39.7985 ;
      RECT 2.1645 40.1305 38.8905 40.2105 ;
      RECT 2.011 40.4285 39.0985 40.4885 ;
      RECT 2.011 40.6685 39.0985 40.7285 ;
      RECT 2.1645 41.0605 38.8905 41.1405 ;
      RECT 2.011 41.3585 39.0985 41.4185 ;
      RECT 2.011 41.5985 39.0985 41.6585 ;
      RECT 2.1645 41.9905 38.8905 42.0705 ;
      RECT 2.011 42.2885 39.0985 42.3485 ;
      RECT 2.011 42.5285 39.0985 42.5885 ;
      RECT 2.1645 42.9205 38.8905 43.0005 ;
      RECT 2.011 43.2185 39.0985 43.2785 ;
      RECT 2.011 43.4585 39.0985 43.5185 ;
      RECT 2.1645 43.8505 38.8905 43.9305 ;
      RECT 9.0295 48.2585 39.4075 48.3185 ;
      RECT 9.0295 48.4985 39.4075 48.5585 ;
      RECT 9.0295 49.1885 39.4075 49.2485 ;
      RECT 9.0295 49.4285 39.4075 49.4885 ;
      RECT 9.0295 50.1185 39.4075 50.1785 ;
      RECT 9.0295 50.3585 39.4075 50.4185 ;
      RECT 9.0295 51.0485 39.4075 51.1085 ;
      RECT 9.0295 51.2885 39.4075 51.3485 ;
      RECT 9.0295 51.9785 39.4075 52.0385 ;
      RECT 9.0295 52.2185 39.4075 52.2785 ;
      RECT 9.0295 52.9085 39.4075 52.9685 ;
      RECT 1.9795 52.95 7.592 53.341 ;
      RECT 9.0295 53.1485 39.4075 53.2085 ;
      RECT 9.0295 53.8385 39.4075 53.8985 ;
      RECT 9.0295 54.0785 39.4075 54.1385 ;
      RECT 1.1965 55.077 6.7125 55.502 ;
      RECT 1.1965 57.417 6.7125 57.842 ;
      RECT 9.0295 57.5285 39.4075 57.5885 ;
      RECT 9.0295 57.7685 39.4075 57.8285 ;
      RECT 9.0295 58.4585 39.4075 58.5185 ;
      RECT 9.0295 58.6985 39.4075 58.7585 ;
      RECT 9.0295 59.3885 39.4075 59.4485 ;
      RECT 9.0295 59.6285 39.4075 59.6885 ;
      RECT 9.0295 60.3185 39.4075 60.3785 ;
      RECT 9.0295 60.5585 39.4075 60.6185 ;
      RECT 9.0295 61.2485 39.4075 61.3085 ;
      RECT 9.0295 61.4885 39.4075 61.5485 ;
      RECT 9.0295 62.1785 39.4075 62.2385 ;
      RECT 9.0295 62.4185 39.4075 62.4785 ;
      RECT 9.0295 63.1085 39.4075 63.1685 ;
      RECT 9.0295 63.3485 39.4075 63.4085 ;
      RECT 4.907 67.25 36.133 67.75 ;
      RECT 4.907 69.05 36.133 69.55 ;
      RECT 4.907 70.85 36.133 71.35 ;
      RECT 4.907 72.65 36.133 73.15 ;
      RECT 4.907 74.45 36.133 74.95 ;
      RECT 4.907 76.25 36.133 76.75 ;
      RECT 4.907 78.95 36.133 79.45 ;
      RECT 4.907 80.75 36.133 81.25 ;
      RECT 4.907 82.55 36.133 83.05 ;
      RECT 4.907 84.35 36.133 84.85 ;
      RECT 4.907 86.15 36.133 86.65 ;
      RECT 4.907 87.95 36.133 88.45 ;
    LAYER M5 ;
      RECT 19.2545 0 19.4545 5.77 ;
      RECT 4.142 0.19 4.218 1.7895 ;
      RECT 25.726 0.19 25.802 1.977 ;
      RECT 26.562 0.19 26.638 1.977 ;
      RECT 23.992 0.276 24.192 65.8355 ;
      RECT 2.542 0.283 2.742 2.7705 ;
      RECT 3.182 0.283 3.382 2.7705 ;
      RECT 3.822 0.283 4.022 2.7705 ;
      RECT 4.658 0.283 4.858 2.7705 ;
      RECT 25.0945 0.283 25.2945 2.7705 ;
      RECT 25.918 0.283 26.118 2.7705 ;
      RECT 26.766 0.283 26.966 2.7705 ;
      RECT 27.446 0.283 27.646 2.7705 ;
      RECT 28.126 0.283 28.326 2.7705 ;
      RECT 28.806 0.283 29.006 2.7705 ;
      RECT 29.486 0.283 29.686 2.7705 ;
      RECT 2.222 0.7215 2.422 3.7815 ;
      RECT 2.862 0.7215 3.062 3.7815 ;
      RECT 3.502 0.7215 3.702 5.0635 ;
      RECT 4.338 0.7215 4.538 5.0635 ;
      RECT 5.2545 0.7215 5.4545 5.775 ;
      RECT 5.6545 0.7215 5.8545 5.775 ;
      RECT 6.0545 0.7215 6.2545 5.775 ;
      RECT 6.4545 0.7215 6.6545 6.4405 ;
      RECT 6.8545 0.7215 7.0545 5.775 ;
      RECT 7.2545 0.7215 7.4545 5.775 ;
      RECT 7.6545 0.7215 7.8545 5.775 ;
      RECT 8.0545 0.7215 8.2545 5.775 ;
      RECT 20.0705 0.7215 20.2705 4.1815 ;
      RECT 22.0545 0.7215 22.2545 4.1005 ;
      RECT 22.4545 0.7215 22.6545 6.4405 ;
      RECT 23.5925 0.7215 23.7925 4.072 ;
      RECT 30.435 0.7215 30.675 4.187 ;
      RECT 31.235 0.7215 31.475 4.187 ;
      RECT 31.655 0.7215 31.855 5.784 ;
      RECT 10.8545 0.73 11.0545 4.1815 ;
      RECT 12.8545 0.73 13.0545 6.4405 ;
      RECT 14.0545 0.73 14.2545 4.1815 ;
      RECT 25.41 0.73 25.61 1.8115 ;
      RECT 26.237 0.73 26.437 1.8115 ;
      RECT 27.106 0.73 27.306 1.8115 ;
      RECT 27.786 0.73 27.986 1.8115 ;
      RECT 28.466 0.73 28.666 1.8115 ;
      RECT 29.146 0.73 29.346 1.8115 ;
      RECT 29.826 0.73 30.026 1.8115 ;
      RECT 35.2545 0.73 35.4545 6.4405 ;
      RECT 36.503 0.73 36.703 4.047 ;
      RECT 37.6625 0.73 37.8625 4.187 ;
      RECT 39.254 0.73 39.454 4.187 ;
      RECT 17.2545 0.7395 17.4545 4.1815 ;
      RECT 18.4545 0.74 18.6545 4.187 ;
      RECT 9.6545 0.7605 9.8545 6.4405 ;
      RECT 16.0545 0.7605 16.2545 6.4405 ;
      RECT 32.0395 0.8035 32.2695 4.187 ;
      RECT 14.463 1.7145 14.703 5.2345 ;
      RECT 39.618 1.7145 39.858 5.2345 ;
      RECT 10.0545 1.899 10.2545 25.0125 ;
      RECT 10.4815 1.899 10.6815 25.0125 ;
      RECT 11.277 1.899 11.477 25.0125 ;
      RECT 11.6545 1.899 11.8545 25.0125 ;
      RECT 12.032 1.899 12.232 5.582 ;
      RECT 12.4095 1.899 12.6095 5.582 ;
      RECT 13.2545 1.899 13.3745 25.0125 ;
      RECT 13.4945 1.899 13.6145 6.769 ;
      RECT 13.7345 1.899 13.8545 25.0125 ;
      RECT 14.913 1.899 15.113 5.595 ;
      RECT 15.29 1.899 15.49 5.595 ;
      RECT 15.6675 1.899 15.8675 5.595 ;
      RECT 17.6345 1.899 17.7545 25.0125 ;
      RECT 17.8745 1.899 17.9945 7.2055 ;
      RECT 18.1145 1.899 18.2345 25.0125 ;
      RECT 19.6545 1.899 19.8545 25.0125 ;
      RECT 21.2545 1.899 21.4545 25.0125 ;
      RECT 22.8545 1.899 23.0545 25.0125 ;
      RECT 24.312 1.899 24.432 25.0125 ;
      RECT 24.552 1.899 24.672 25.0125 ;
      RECT 34.4545 1.899 34.6545 5.7375 ;
      RECT 34.8545 1.899 35.0545 5.7375 ;
      RECT 35.6545 1.899 35.8545 25.0125 ;
      RECT 36.8545 1.899 37.0545 25.0125 ;
      RECT 37.2545 1.899 37.4545 25.0125 ;
      RECT 38.4515 1.899 38.6515 6.757 ;
      RECT 38.8545 1.899 39.0545 25.0125 ;
      RECT 16.4545 1.9025 16.5745 25.0125 ;
      RECT 16.6945 1.9025 16.8145 7.2055 ;
      RECT 16.9345 1.9025 17.0545 25.0125 ;
      RECT 24.835 3.262 25.075 5.7615 ;
      RECT 25.235 3.262 25.475 5.7615 ;
      RECT 26.835 3.262 27.075 5.784 ;
      RECT 28.035 3.262 28.275 5.784 ;
      RECT 28.44 3.262 28.67 5.784 ;
      RECT 28.8345 3.262 29.0745 6.454 ;
      RECT 30.055 3.262 30.255 5.784 ;
      RECT 3.822 3.7325 4.022 4.7875 ;
      RECT 20.8385 4.253 21.0385 25.0125 ;
      RECT 21.7945 4.253 21.8745 25.0125 ;
      RECT 25.7945 4.395 25.8745 25.3665 ;
      RECT 36.1945 4.395 36.2745 25.3665 ;
      RECT 23.3945 4.4 23.4745 63.8555 ;
      RECT 29.6345 4.4645 29.7145 35.023 ;
      RECT 30.4345 4.4645 30.5145 35.023 ;
      RECT 23.2345 4.5745 23.3145 54.711 ;
      RECT 8.4545 4.789 8.6545 25.0125 ;
      RECT 26.0545 4.789 26.1745 25.0125 ;
      RECT 26.3145 4.789 26.4345 25.0195 ;
      RECT 26.5545 4.789 26.6745 25.0195 ;
      RECT 27.252 4.789 27.372 25.0125 ;
      RECT 27.4945 4.789 27.6145 6.769 ;
      RECT 27.7345 4.789 27.8545 25.0125 ;
      RECT 29.2545 4.789 29.4545 25.0125 ;
      RECT 29.8445 4.789 29.9245 25.0125 ;
      RECT 30.6445 4.789 30.7245 25.0125 ;
      RECT 30.8545 4.789 31.0545 25.0125 ;
      RECT 31.1945 4.789 31.2745 6.768 ;
      RECT 31.4145 4.789 31.5345 15.999 ;
      RECT 32.0575 4.789 32.2575 25.0125 ;
      RECT 32.4545 4.789 32.6545 25.0125 ;
      RECT 32.8875 4.789 33.0875 25.0125 ;
      RECT 33.671 4.789 33.871 25.0125 ;
      RECT 34.0545 4.789 34.2545 25.0125 ;
      RECT 36.0345 4.789 36.1145 25.0125 ;
      RECT 37.8445 4.9025 37.9245 15.999 ;
      RECT 1.6945 5.2605 1.8945 15.4775 ;
      RECT 39.2145 5.2605 39.4145 6.077 ;
      RECT 3.2545 5.271 3.4545 6.4405 ;
      RECT 18.3945 5.637 18.4745 14.961 ;
      RECT 20.0705 5.79 20.2705 25.0125 ;
      RECT 18.5945 5.828 18.6745 25.0125 ;
      RECT 2.6445 6.27 2.7245 15.999 ;
      RECT 5.8445 6.27 5.9245 15.999 ;
      RECT 9.0445 6.27 9.1245 15.999 ;
      RECT 12.2445 6.27 12.3245 15.999 ;
      RECT 15.4445 6.27 15.5245 15.999 ;
      RECT 19.2545 6.27 19.4545 25.0125 ;
      RECT 28.2445 6.27 28.3245 15.999 ;
      RECT 34.6445 6.27 34.7245 15.999 ;
      RECT 2.0545 6.271 2.2545 25.0125 ;
      RECT 3.6545 6.271 3.8545 25.0125 ;
      RECT 4.0725 6.271 4.2725 25.0125 ;
      RECT 4.8575 6.271 5.0575 25.0125 ;
      RECT 5.2545 6.271 5.4545 25.0125 ;
      RECT 6.8545 6.271 7.0545 25.0125 ;
      RECT 7.2555 6.271 7.4555 25.0125 ;
      RECT 8.051 6.271 8.251 25.0125 ;
      RECT 14.4545 6.271 14.5745 25.0125 ;
      RECT 14.6945 6.271 14.8145 6.769 ;
      RECT 14.9345 6.271 15.0545 25.0125 ;
      RECT 25.6345 6.271 25.7145 25.0125 ;
      RECT 24.9945 6.283 25.1145 14.7945 ;
      RECT 2.8545 6.6715 3.0545 25.0125 ;
      RECT 4.4545 6.6715 4.6545 25.0125 ;
      RECT 5.5945 6.6715 5.6745 14.961 ;
      RECT 6.0545 6.6715 6.2545 25.0125 ;
      RECT 7.6545 6.6715 7.8545 25.0125 ;
      RECT 8.7945 6.6715 8.8745 14.961 ;
      RECT 9.2545 6.6715 9.4545 25.0125 ;
      RECT 10.8545 6.6715 11.0545 25.0125 ;
      RECT 11.9945 6.6715 12.0745 14.961 ;
      RECT 12.4545 6.6715 12.6545 25.0125 ;
      RECT 14.0545 6.6715 14.2545 25.0125 ;
      RECT 15.203 6.6715 15.283 14.961 ;
      RECT 15.6545 6.6715 15.8545 25.0125 ;
      RECT 17.2545 6.6715 17.4545 25.0125 ;
      RECT 18.8545 6.6715 19.0545 25.0125 ;
      RECT 20.4545 6.6715 20.6545 25.0125 ;
      RECT 21.5945 6.6715 21.6745 14.961 ;
      RECT 22.0545 6.6715 22.2545 25.0125 ;
      RECT 23.6545 6.6715 23.8545 25.0125 ;
      RECT 24.7945 6.6715 24.8745 14.961 ;
      RECT 25.2545 6.6715 25.4545 25.0125 ;
      RECT 26.8545 6.6715 27.0545 25.0125 ;
      RECT 27.9945 6.6715 28.0745 14.961 ;
      RECT 28.4545 6.6715 28.6545 25.0125 ;
      RECT 30.0545 6.6715 30.2545 25.0125 ;
      RECT 31.6545 6.6715 31.8545 25.0125 ;
      RECT 33.2545 6.6715 33.4545 25.0125 ;
      RECT 34.3945 6.6715 34.4745 14.961 ;
      RECT 34.8545 6.6715 35.0545 25.0125 ;
      RECT 36.4545 6.6715 36.6545 25.0125 ;
      RECT 38.0545 6.6715 38.2545 25.0125 ;
      RECT 22.4575 6.687 22.6575 25.0125 ;
      RECT 28.8575 6.687 29.0575 25.0125 ;
      RECT 35.2575 6.687 35.4575 25.0125 ;
      RECT 3.2575 6.752 3.4575 25.0125 ;
      RECT 6.4575 6.752 6.6575 25.0125 ;
      RECT 9.6575 6.752 9.8575 25.0125 ;
      RECT 12.8575 6.752 13.0575 25.0125 ;
      RECT 16.0575 6.7595 16.2575 25.0125 ;
      RECT 31.1945 6.997 31.2745 14.961 ;
      RECT 38.4575 7.6895 38.6575 25.0125 ;
      RECT 13.4945 8.271 13.6145 8.769 ;
      RECT 14.6945 8.271 14.8145 8.769 ;
      RECT 16.6945 8.271 16.8145 8.769 ;
      RECT 17.8745 8.271 17.9945 8.769 ;
      RECT 27.4945 8.271 27.6145 8.769 ;
      RECT 13.4945 10.271 13.6145 10.769 ;
      RECT 14.6945 10.271 14.8145 10.769 ;
      RECT 16.6945 10.271 16.8145 10.769 ;
      RECT 17.8745 10.271 17.9945 10.769 ;
      RECT 27.4945 10.271 27.6145 10.769 ;
      RECT 13.4945 12.271 13.6145 12.769 ;
      RECT 14.6945 12.271 14.8145 12.769 ;
      RECT 16.6945 12.271 16.8145 12.769 ;
      RECT 17.8745 12.271 17.9945 12.769 ;
      RECT 27.4945 12.271 27.6145 12.769 ;
      RECT 13.4945 14.271 13.6145 14.769 ;
      RECT 14.6945 14.271 14.8145 14.769 ;
      RECT 16.6945 14.271 16.8145 14.769 ;
      RECT 17.8745 14.271 17.9945 14.769 ;
      RECT 27.4945 14.271 27.6145 14.769 ;
      RECT 2.3845 15.288 2.4645 25.0125 ;
      RECT 5.5845 15.288 5.6645 25.0125 ;
      RECT 8.7845 15.288 8.8645 25.0125 ;
      RECT 11.9845 15.288 12.0645 25.0125 ;
      RECT 15.203 15.288 15.323 25.0125 ;
      RECT 18.3545 15.288 18.4745 25.0125 ;
      RECT 21.5845 15.288 21.6645 25.0125 ;
      RECT 27.9745 15.288 28.0945 25.0125 ;
      RECT 31.1845 15.288 31.2645 25.0125 ;
      RECT 34.3845 15.288 34.4645 25.0125 ;
      RECT 37.5845 15.288 37.6645 25.0125 ;
      RECT 24.792 15.797 24.912 25.0125 ;
      RECT 13.4945 16.271 13.6145 16.769 ;
      RECT 14.6945 16.271 14.8145 16.769 ;
      RECT 16.6945 16.271 16.8145 16.769 ;
      RECT 17.8745 16.271 17.9945 16.769 ;
      RECT 27.4945 16.271 27.6145 16.769 ;
      RECT 2.5945 16.3015 2.6745 25.0125 ;
      RECT 5.7945 16.3015 5.8745 25.0125 ;
      RECT 8.9945 16.3015 9.0745 25.0125 ;
      RECT 12.1945 16.3015 12.2745 25.0125 ;
      RECT 15.443 16.3015 15.523 25.0125 ;
      RECT 25.032 16.3015 25.112 25.0125 ;
      RECT 28.2445 16.3015 28.3245 25.0125 ;
      RECT 31.3945 16.3015 31.4745 25.0125 ;
      RECT 34.5945 16.3015 34.6745 25.0125 ;
      RECT 37.7945 16.3015 37.8745 25.0125 ;
      RECT 13.4945 18.271 13.6145 18.769 ;
      RECT 14.6945 18.271 14.8145 18.769 ;
      RECT 16.6945 18.271 16.8145 18.769 ;
      RECT 17.8745 18.271 17.9945 18.769 ;
      RECT 27.4945 18.271 27.6145 18.769 ;
      RECT 13.4945 19.271 13.6145 19.769 ;
      RECT 14.6945 19.271 14.8145 19.769 ;
      RECT 16.6945 19.271 16.8145 19.769 ;
      RECT 17.8745 19.271 17.9945 19.769 ;
      RECT 27.4945 19.271 27.6145 19.769 ;
      RECT 13.4945 20.271 13.6145 20.769 ;
      RECT 14.6945 20.271 14.8145 20.769 ;
      RECT 16.6945 20.271 16.8145 20.769 ;
      RECT 17.8745 20.271 17.9945 20.769 ;
      RECT 27.4945 20.271 27.6145 20.769 ;
      RECT 13.4945 21.271 13.6145 21.769 ;
      RECT 14.6945 21.271 14.8145 21.769 ;
      RECT 16.6945 21.271 16.8145 21.769 ;
      RECT 17.8745 21.271 17.9945 21.769 ;
      RECT 27.4945 21.271 27.6145 21.769 ;
      RECT 13.4945 22.271 13.6145 22.769 ;
      RECT 14.6945 22.271 14.8145 22.769 ;
      RECT 16.6945 22.271 16.8145 22.769 ;
      RECT 17.8745 22.271 17.9945 22.769 ;
      RECT 27.4945 22.271 27.6145 22.769 ;
      RECT 13.4945 24.271 13.6145 24.769 ;
      RECT 14.6945 24.271 14.8145 24.769 ;
      RECT 16.6945 24.271 16.8145 24.769 ;
      RECT 17.8745 24.271 17.9945 24.769 ;
      RECT 27.4945 24.271 27.6145 24.769 ;
      RECT 24.7945 25.213 24.8745 34.3185 ;
      RECT 27.9945 25.213 28.0745 34.3185 ;
      RECT 31.1945 25.213 31.2745 34.3185 ;
      RECT 34.3945 25.213 34.4745 34.311 ;
      RECT 31.4425 25.236 31.5225 34.311 ;
      RECT 13.2545 25.2465 13.3745 44.769 ;
      RECT 13.4945 25.2465 13.6145 26.511 ;
      RECT 13.7345 25.2465 13.8545 44.769 ;
      RECT 14.4545 25.2465 14.5745 44.769 ;
      RECT 14.9345 25.2465 15.0545 44.769 ;
      RECT 16.4545 25.2465 16.5745 44.769 ;
      RECT 16.9345 25.2465 17.0545 44.769 ;
      RECT 17.6345 25.2465 17.7545 44.769 ;
      RECT 18.1145 25.2465 18.2345 44.769 ;
      RECT 34.6425 25.249 34.7225 34.311 ;
      RECT 37.8425 25.249 37.9225 34.311 ;
      RECT 26.0145 25.2535 26.2145 44.7775 ;
      RECT 2.5945 25.266 2.6745 34.3185 ;
      RECT 5.5945 25.266 5.6745 34.3185 ;
      RECT 5.7945 25.266 5.8745 34.3185 ;
      RECT 8.7945 25.266 8.8745 34.3185 ;
      RECT 8.9945 25.266 9.0745 34.3185 ;
      RECT 11.9945 25.266 12.0745 34.3185 ;
      RECT 12.1945 25.266 12.2745 34.3185 ;
      RECT 15.203 25.266 15.283 34.3185 ;
      RECT 18.3945 25.266 18.4745 34.3185 ;
      RECT 18.5945 25.266 18.6745 34.3185 ;
      RECT 21.5945 25.266 21.6745 34.3185 ;
      RECT 21.7945 25.266 21.8745 34.3185 ;
      RECT 29.8445 25.266 29.9245 34.311 ;
      RECT 30.6445 25.266 30.7245 34.311 ;
      RECT 1.6945 25.271 1.8945 34.8275 ;
      RECT 2.0545 25.271 2.2545 44.769 ;
      RECT 2.8545 25.271 3.0545 44.3625 ;
      RECT 3.2545 25.271 3.4545 33.9275 ;
      RECT 3.6545 25.271 3.8545 44.769 ;
      RECT 4.0835 25.271 4.2835 44.769 ;
      RECT 4.4545 25.271 4.6545 44.3625 ;
      RECT 4.8495 25.271 5.0495 44.769 ;
      RECT 5.2545 25.271 5.4545 44.769 ;
      RECT 6.0545 25.271 6.2545 44.3625 ;
      RECT 6.4545 25.271 6.6545 33.9275 ;
      RECT 6.8545 25.271 7.0545 44.769 ;
      RECT 7.2545 25.271 7.4545 44.769 ;
      RECT 7.6545 25.271 7.8545 44.363 ;
      RECT 8.0545 25.271 8.2545 44.769 ;
      RECT 8.4545 25.271 8.6545 44.769 ;
      RECT 9.2545 25.271 9.4545 44.363 ;
      RECT 9.6545 25.271 9.8545 33.9275 ;
      RECT 10.0545 25.271 10.2545 44.769 ;
      RECT 10.4385 25.271 10.6385 44.769 ;
      RECT 10.8545 25.271 11.0545 44.363 ;
      RECT 11.259 25.271 11.459 44.769 ;
      RECT 11.6545 25.271 11.8545 44.769 ;
      RECT 12.4545 25.271 12.6545 44.363 ;
      RECT 12.8545 25.271 13.0545 44.769 ;
      RECT 14.0545 25.271 14.2545 44.363 ;
      RECT 15.6545 25.271 15.8545 44.363 ;
      RECT 16.0345 25.271 16.2745 44.769 ;
      RECT 17.2545 25.271 17.4545 44.363 ;
      RECT 18.8545 25.271 19.0545 44.363 ;
      RECT 19.2545 25.271 19.4545 44.769 ;
      RECT 19.6545 25.271 19.8545 44.769 ;
      RECT 20.0545 25.271 20.2545 44.769 ;
      RECT 20.4545 25.271 20.6545 44.363 ;
      RECT 20.8545 25.271 21.0545 44.769 ;
      RECT 21.2545 25.271 21.4545 44.769 ;
      RECT 22.0545 25.271 22.2545 44.363 ;
      RECT 22.4545 25.271 22.6545 44.769 ;
      RECT 22.8545 25.271 23.0545 44.769 ;
      RECT 23.6545 25.271 23.8545 44.363 ;
      RECT 24.312 25.271 24.432 44.769 ;
      RECT 24.552 25.271 24.672 44.769 ;
      RECT 25.0145 25.271 25.1345 34.3005 ;
      RECT 25.2545 25.271 25.4545 44.363 ;
      POLYGON 26.6745 25.271 26.6745 44.3625 26.6545 44.3625 26.6545 44.769 26.4545 44.769 26.4545 44.3625 26.4345 44.3625 26.4345 25.271 ;
      RECT 26.8545 25.271 27.0545 44.3625 ;
      RECT 27.2545 25.271 27.3745 44.769 ;
      RECT 27.7345 25.271 27.8545 44.769 ;
      RECT 28.4545 25.271 28.6545 44.3625 ;
      RECT 28.8545 25.271 29.0545 44.769 ;
      RECT 29.2545 25.271 29.4545 44.769 ;
      RECT 30.0545 25.271 30.2545 44.3625 ;
      RECT 30.8545 25.271 31.0545 44.769 ;
      RECT 31.6545 25.271 31.8545 44.3625 ;
      RECT 32.0545 25.271 32.2545 33.9275 ;
      RECT 32.4545 25.271 32.6545 44.769 ;
      RECT 32.8545 25.271 33.0545 44.769 ;
      RECT 33.2545 25.271 33.4545 44.3625 ;
      RECT 33.6545 25.271 33.8545 44.769 ;
      RECT 34.0545 25.271 34.2545 44.769 ;
      RECT 34.8545 25.271 35.0545 44.3625 ;
      RECT 35.2545 25.271 35.4545 33.9275 ;
      RECT 35.6545 25.271 35.8545 44.769 ;
      RECT 36.4545 25.271 36.6545 44.3625 ;
      RECT 36.8545 25.271 37.0545 44.769 ;
      RECT 37.2545 25.271 37.4545 44.769 ;
      RECT 38.0545 25.271 38.2545 44.3625 ;
      RECT 38.4545 25.271 38.6545 33.945 ;
      RECT 38.8545 25.271 39.0545 44.769 ;
      RECT 25.6545 26.0215 25.8545 44.769 ;
      RECT 36.0545 26.0215 36.2545 44.769 ;
      RECT 13.4945 27.771 13.6145 28.269 ;
      RECT 39.5745 33.7605 39.7745 46.7705 ;
      RECT 39.9745 33.7605 40.1745 46.7705 ;
      RECT 32.0545 34.7555 32.2545 44.769 ;
      RECT 35.2545 34.7575 35.4545 44.769 ;
      RECT 6.4545 34.7635 6.6545 44.769 ;
      RECT 18.3945 34.7665 18.4745 44.77 ;
      RECT 27.9945 34.7665 28.0745 44.77 ;
      RECT 8.7945 34.7675 8.8745 44.77 ;
      RECT 5.5945 34.7695 5.6745 44.77 ;
      RECT 11.9945 34.7695 12.0745 44.77 ;
      RECT 34.3945 34.7695 34.4745 44.77 ;
      RECT 2.3945 34.77 2.4745 44.77 ;
      RECT 37.5945 34.77 37.6745 44.77 ;
      RECT 3.2545 34.771 3.4545 44.769 ;
      RECT 9.6545 34.771 9.8545 44.769 ;
      RECT 13.4945 34.771 13.6145 35.269 ;
      RECT 15.1745 34.771 15.2945 44.769 ;
      RECT 38.4545 34.771 38.6545 44.769 ;
      RECT 24.792 34.783 24.912 44.757 ;
      RECT 2.5945 34.8695 2.6745 44.363 ;
      RECT 5.7945 34.8695 5.8745 44.363 ;
      RECT 8.9945 34.8695 9.0745 44.363 ;
      RECT 12.1945 34.8695 12.2745 44.363 ;
      RECT 15.443 34.8695 15.523 44.363 ;
      RECT 18.5945 34.8695 18.6745 44.363 ;
      RECT 21.7945 34.8695 21.8745 44.363 ;
      RECT 25.032 34.8695 25.112 44.363 ;
      RECT 28.2445 34.8695 28.3245 44.363 ;
      RECT 31.3945 34.8695 31.4745 44.363 ;
      RECT 34.5945 34.8695 34.6745 44.363 ;
      RECT 37.7945 34.8695 37.8745 44.363 ;
      RECT 21.5945 35.1935 21.6745 44.77 ;
      RECT 31.1945 35.1935 31.2745 44.77 ;
      RECT 29.6545 35.6155 29.8545 44.769 ;
      RECT 30.4545 35.6155 30.6545 44.769 ;
      RECT 13.4945 36.271 13.6145 36.769 ;
      RECT 13.4945 38.271 13.6145 38.769 ;
      RECT 13.4945 40.271 13.6145 40.769 ;
      RECT 13.4945 42.271 13.6145 42.769 ;
      RECT 13.4945 44.271 13.6145 44.769 ;
      RECT 9.2545 44.719 9.4545 64.866 ;
      RECT 10.8545 45.27 11.0545 55.5655 ;
      RECT 14.0545 45.27 14.2545 55.5655 ;
      RECT 17.2545 45.27 17.4545 55.5655 ;
      RECT 20.4545 45.27 20.6545 55.5655 ;
      RECT 23.6545 45.27 23.8545 55.5655 ;
      RECT 26.8545 45.27 27.0545 55.5655 ;
      RECT 30.0545 45.27 30.2545 55.5655 ;
      RECT 33.2545 45.27 33.4545 55.5655 ;
      RECT 36.4545 45.27 36.6545 55.5655 ;
      RECT 12.4545 46.27 12.6545 64.866 ;
      RECT 15.6545 46.27 15.8545 64.866 ;
      RECT 18.8545 46.27 19.0545 64.866 ;
      RECT 22.0545 46.27 22.2545 64.866 ;
      RECT 25.2545 46.27 25.4545 64.866 ;
      RECT 28.4545 46.27 28.6545 64.866 ;
      RECT 31.6545 46.27 31.8545 64.866 ;
      RECT 34.8545 46.27 35.0545 64.866 ;
      RECT 38.0545 46.27 38.2545 64.866 ;
      RECT 9.6345 46.2915 9.7145 64.2505 ;
      RECT 9.7945 46.2915 9.8745 63.855 ;
      RECT 12.8345 46.2915 12.9145 64.2505 ;
      RECT 12.9945 46.2915 13.0745 63.855 ;
      RECT 16.0345 46.2915 16.1145 64.2505 ;
      RECT 16.1945 46.2915 16.2745 63.855 ;
      RECT 19.2345 46.2915 19.3145 64.2505 ;
      RECT 19.3945 46.2915 19.4745 63.855 ;
      RECT 22.4345 46.2915 22.5145 64.2505 ;
      RECT 22.5945 46.2915 22.6745 63.855 ;
      RECT 25.6345 46.2915 25.7145 64.2505 ;
      RECT 25.7945 46.2915 25.8745 63.855 ;
      RECT 28.8345 46.2915 28.9145 64.2505 ;
      RECT 28.9945 46.2915 29.0745 63.855 ;
      RECT 32.0345 46.2915 32.1145 64.2505 ;
      RECT 32.1945 46.2915 32.2745 63.855 ;
      RECT 35.2345 46.2915 35.3145 64.2505 ;
      RECT 35.3945 46.2915 35.4745 63.855 ;
      RECT 38.4345 46.2915 38.5145 64.2505 ;
      RECT 38.5945 46.2915 38.6745 63.855 ;
      RECT 20.0345 46.9555 20.1145 54.606 ;
      RECT 39.2345 46.9555 39.3145 54.606 ;
      RECT 39.6545 47.127 39.8545 55.592 ;
      RECT 1.1965 52.2245 1.5965 56.86 ;
      RECT 1.9425 52.2245 2.3425 56.86 ;
      RECT 2.6885 52.2245 3.0885 56.86 ;
      RECT 3.4345 52.2245 3.8345 56.86 ;
      RECT 4.1805 52.2245 4.5805 56.86 ;
      RECT 4.9265 52.2245 5.3265 56.86 ;
      RECT 5.6725 52.2245 6.0725 56.86 ;
      RECT 6.4185 52.2245 6.8185 56.86 ;
      RECT 7.164 52.95 7.364 56.165 ;
      RECT 10.8545 56.271 11.0545 56.769 ;
      RECT 14.0545 56.271 14.2545 56.769 ;
      RECT 17.2545 56.271 17.4545 56.769 ;
      RECT 20.4545 56.271 20.6545 56.769 ;
      RECT 23.6545 56.271 23.8545 56.769 ;
      RECT 26.8545 56.271 27.0545 56.769 ;
      RECT 30.0545 56.271 30.2545 56.769 ;
      RECT 33.2545 56.271 33.4545 56.769 ;
      RECT 36.4545 56.271 36.6545 56.769 ;
      RECT 39.6545 56.271 39.8545 56.769 ;
      RECT 39.3945 57.165 39.4745 63.9145 ;
      RECT 10.5945 57.185 10.6745 63.8555 ;
      RECT 13.7945 57.185 13.8745 63.8555 ;
      RECT 16.9945 57.185 17.0745 63.8555 ;
      RECT 20.1945 57.185 20.2745 63.8555 ;
      RECT 4.8325 59.391 5.2325 61.244 ;
      RECT 9.2545 65.271 9.4545 65.769 ;
      RECT 12.4545 65.271 12.6545 65.769 ;
      RECT 15.6545 65.271 15.8545 65.769 ;
      RECT 18.8545 65.271 19.0545 65.769 ;
      RECT 22.0545 65.271 22.2545 65.769 ;
      RECT 25.2545 65.271 25.4545 65.769 ;
      RECT 28.4545 65.271 28.6545 65.769 ;
      RECT 31.6545 65.271 31.8545 65.769 ;
      RECT 34.8545 65.271 35.0545 65.769 ;
      RECT 38.0545 65.271 38.2545 65.769 ;
      RECT 0.3 66.375 20.28 66.825 ;
      RECT 20.76 66.375 40.74 66.825 ;
      RECT 5.6 68.175 20.28 68.625 ;
      RECT 20.76 68.175 35.44 68.625 ;
      RECT 0.3 69.075 20.28 69.525 ;
      RECT 20.76 69.075 40.74 69.525 ;
      RECT 5.6 69.975 20.28 70.425 ;
      RECT 20.76 69.975 35.44 70.425 ;
      RECT 0.3 70.875 20.28 71.325 ;
      RECT 20.76 70.875 40.74 71.325 ;
      RECT 5.6 71.775 20.28 72.225 ;
      RECT 20.76 71.775 35.44 72.225 ;
      RECT 0.3 72.675 20.28 73.125 ;
      RECT 20.76 72.675 40.74 73.125 ;
      RECT 5.6 73.575 20.28 74.025 ;
      RECT 20.76 73.575 35.44 74.025 ;
      RECT 0.3 74.475 20.28 74.925 ;
      RECT 20.76 74.475 40.74 74.925 ;
      RECT 5.6 75.375 20.28 75.825 ;
      RECT 20.76 75.375 35.44 75.825 ;
      RECT 0.3 76.275 20.28 76.725 ;
      RECT 20.76 76.275 40.74 76.725 ;
      RECT 0.3 77.175 20.28 77.625 ;
      RECT 20.76 77.175 40.74 77.625 ;
      RECT 0.3 78.075 20.28 78.525 ;
      RECT 20.76 78.075 40.74 78.525 ;
      RECT 0.3 78.975 20.28 79.425 ;
      RECT 20.76 78.975 40.74 79.425 ;
      RECT 5.601 79.875 20.28 80.325 ;
      RECT 20.76 79.875 35.439 80.325 ;
      RECT 0.3 80.775 20.28 81.225 ;
      RECT 20.76 80.775 40.74 81.225 ;
      RECT 5.601 81.675 20.28 82.125 ;
      RECT 20.76 81.675 35.439 82.125 ;
      RECT 0.3 82.575 20.28 83.025 ;
      RECT 20.76 82.575 40.74 83.025 ;
      RECT 5.601 83.475 20.28 83.925 ;
      RECT 20.76 83.475 35.439 83.925 ;
      RECT 0.3 84.375 20.28 84.825 ;
      RECT 20.76 84.375 40.74 84.825 ;
      RECT 5.601 85.275 20.28 85.725 ;
      RECT 20.76 85.275 35.439 85.725 ;
      RECT 0.3 86.175 20.28 86.625 ;
      RECT 20.76 86.175 40.74 86.625 ;
      RECT 5.601 87.075 20.28 87.525 ;
      RECT 20.76 87.075 35.439 87.525 ;
    LAYER M6 ;
      RECT 0.3 19.27 40.74 19.77 ;
      RECT 0.3 20.27 40.74 20.77 ;
      RECT 0.3 21.27 40.74 21.77 ;
    LAYER M0 ;
      RECT MASK 1 0 0 41.04 90 ;
      RECT MASK 2 0 0 41.04 90 ;
    LAYER LUP_015U ;
      RECT 3.944 66.33 37.096 89.49 ;
  END
END dwc_ddrphy_vrefdacref

END LIBRARY
