# LEF OUT API 
# Creation Date : Thu Apr 11 19:56:15 IST 2019
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_zcalana
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_zcalana 0 0 ;
  SYMMETRY X Y ;
  SIZE 82.08 BY 90 ;
  PIN ZCalPDLoad
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.7736 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M4 ;
      ANTENNAMAXAREACAR 0 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 81.68 47.428 82.08 47.828 ;
    END
  END ZCalPDLoad
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M6 ;
        RECT 0.3 0.27 81.78 0.77 ;
        RECT 0.3 2.27 81.78 2.77 ;
        RECT 0.3 6.27 81.78 6.77 ;
        RECT 0.3 8.27 81.78 8.77 ;
        RECT 0.3 10.27 81.78 10.77 ;
        RECT 0.3 12.27 81.78 12.77 ;
        RECT 0.3 14.27 81.78 14.77 ;
        RECT 0.3 16.27 81.78 16.77 ;
        RECT 0.3 18.27 81.78 18.77 ;
        RECT 0.3 19.269 81.78 19.769 ;
        RECT 0.3 22.27 81.78 22.77 ;
        RECT 0.3 24.27 81.78 24.77 ;
        RECT 0.3 26.27 81.78 26.77 ;
        RECT 0.3 28.77 81.78 29.27 ;
        RECT 32.589 40.395 81.78 40.845 ;
        RECT 0.3 44.895 81.78 45.345 ;
        RECT 0.3 46.695 81.78 47.145 ;
        RECT 0.3 48.54 81.78 48.99 ;
        RECT 0.3 51.637 81.78 52.087 ;
        RECT 0.3 53.437 81.78 53.887 ;
        RECT 0.3 55.237 81.78 55.687 ;
        RECT 0.3 57.037 81.78 57.487 ;
        RECT 0.3 58.837 81.78 59.287 ;
        RECT 0.3 59.895 81.78 60.345 ;
        RECT 0.3 61.695 81.78 62.145 ;
        RECT 0.3 63.495 81.78 63.945 ;
        RECT 0.3 65.317 81.78 65.767 ;
        RECT 0.3 67.117 81.78 67.567 ;
        RECT 0.3 68.917 81.78 69.367 ;
        RECT 0.3 69.975 81.78 70.425 ;
        RECT 0.3 71.775 81.78 72.225 ;
        RECT 0.3 73.575 81.78 74.025 ;
        RECT 0.3 75.375 81.78 75.825 ;
        RECT 0.3 77.175 81.78 77.625 ;
        RECT 0.3 78.975 81.78 79.425 ;
        RECT 0.3 80.775 81.78 81.225 ;
        RECT 0.3 82.575 81.78 83.025 ;
        RECT 0.3 84.375 81.78 84.825 ;
        RECT 0.3 86.175 81.78 86.625 ;
        RECT 0.3 87.975 81.78 88.425 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 33.77 11.389 34.27 ;
        RECT 0.3 36.27 11.389 36.77 ;
        RECT 0.3 40.395 11.389 40.845 ;
        RECT 0.3 42.195 11.389 42.645 ;
        RECT 0.3 43.995 11.389 44.445 ;
    END
    PORT
      LAYER M6 ;
        RECT 32.589 33.77 81.78 34.27 ;
        RECT 32.589 36.27 81.78 36.77 ;
        RECT 0.3 38.153 81.78 38.603 ;
        RECT 32.589 42.195 81.78 42.645 ;
        RECT 32.589 43.995 81.78 44.445 ;
        RECT 10.542 49.57 81.78 50.02 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.3 60.795 81.78 61.245 ;
        RECT 0.3 64.395 81.78 64.845 ;
        RECT 0.3 66.217 81.78 66.667 ;
        RECT 0.3 68.017 81.78 68.467 ;
    END
    PORT
      LAYER M6 ;
        RECT 32.589 35.27 42.589 35.77 ;
        RECT 32.589 39.32 42.589 39.77 ;
        RECT 32.589 41.295 42.589 41.745 ;
        RECT 32.589 43.095 42.589 43.545 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 62.595 81.78 63.045 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 1.27 81.78 1.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 7.27 81.78 7.77 ;
        RECT 0.3 9.27 81.78 9.77 ;
        RECT 0.3 11.27 81.78 11.77 ;
        RECT 0.3 13.27 42.589 13.77 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 35.27 11.389 35.77 ;
        RECT 0.3 39.32 11.389 39.77 ;
        RECT 0.3 41.295 11.389 41.745 ;
        RECT 0.3 43.095 11.389 43.545 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 45.795 81.78 46.245 ;
        RECT 0.3 47.64 81.78 48.09 ;
        RECT 0.3 50.737 81.78 51.187 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 15.27 42.589 15.77 ;
        RECT 0.3 17.27 42.589 17.77 ;
        RECT 0.3 23.27 42.589 23.77 ;
        RECT 0.3 25.27 42.589 25.77 ;
        RECT 0.3 27.27 42.589 27.77 ;
        RECT 0.3 37.253 42.589 37.703 ;
        RECT 0.3 52.537 81.78 52.987 ;
        RECT 0.3 54.337 81.78 54.787 ;
        RECT 0.3 56.137 81.78 56.587 ;
        RECT 0.3 57.937 81.78 58.387 ;
    END
  END VDD
  PIN ZCalPULoad
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.34452 LAYER M6 ;
    ANTENNADIFFAREA 0 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 0 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0.3 49.57 9.9545 50.02 ;
    END
  END ZCalPULoad
  PIN csrZCalCompGainCurrAdj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.076 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 652.35 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 34.618 0 34.694 0.114 ;
    END
  END csrZCalCompGainCurrAdj[0]
  PIN csrZCalCompGainCurrAdj{1}
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06688 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 670.133 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 34.77 0 34.846 0.114 ;
    END
  END csrZCalCompGainCurrAdj[1]
  PIN csrZCalCompGainCurrAdj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05776 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 711.659 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 35.074 0 35.15 0.114 ;
    END
  END csrZCalCompGainCurrAdj[2]
  PIN csrZCalCompGainCurrAdj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.04864 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 727.248 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 35.226 0 35.302 0.114 ;
    END
  END csrZCalCompGainCurrAdj[3]
  PIN ZCalAnaEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.08512 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 639.936 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 34.466 0 34.542 0.114 ;
    END
  END ZCalAnaEn
  PIN ZCalPUEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21052 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 235.699 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 45.258 0 45.334 0.114 ;
    END
  END ZCalPUEn
  PIN ZCalPDEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21052 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 234.169 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 45.41 0 45.486 0.114 ;
    END
  END ZCalPDEn
  PIN ZCalCompEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21052 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 226.883 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 45.562 0 45.638 0.114 ;
    END
  END ZCalCompEn
  PIN ZCalCompVOHDAC[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1672 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 182.452 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 69.426 0 69.502 0.114 ;
    END
  END ZCalCompVOHDAC[0]
  PIN ZCalCompVOHDAC[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18544 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 196.393 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 69.882 0 69.958 0.114 ;
    END
  END ZCalCompVOHDAC[1]
  PIN ZCalCompVOHDAC[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1684539375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 185.646 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 70.186 0 70.262 0.114 ;
    END
  END ZCalCompVOHDAC[2]
  PIN ZCalCompVOHDAC[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18544 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 208.046 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 70.642 0 70.718 0.114 ;
    END
  END ZCalCompVOHDAC[3]
  PIN ZCalCompVOHDAC[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1672 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 186.794 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 71.098 0 71.174 0.114 ;
    END
  END ZCalCompVOHDAC[4]
  PIN ZCalCompVOHDAC[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18544 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 197.331 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 71.402 0 71.478 0.114 ;
    END
  END ZCalCompVOHDAC[5]
  PIN ZCalCompVOHDAC[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1672 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 181.809 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 72.01 0 72.086 0.114 ;
    END
  END ZCalCompVOHDAC[6]
  PIN csrZCalCompVrefDAC[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20368 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 217.66 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 69.274 0 69.35 0.114 ;
    END
  END csrZCalCompVrefDAC[0]
  PIN csrZCalCompVrefDAC[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.22192 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 228.892 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 69.578 0 69.654 0.114 ;
    END
  END csrZCalCompVrefDAC[1]
  PIN csrZCalCompVrefDAC[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20368 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 212.569 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 70.034 0 70.11 0.114 ;
    END
  END csrZCalCompVrefDAC[2]
  PIN csrZCalCompVrefDAC[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.22192 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 230.158 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 70.49 0 70.566 0.114 ;
    END
  END csrZCalCompVrefDAC[3]
  PIN csrZCalCompVrefDAC[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20368 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 231.516 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 70.794 0 70.87 0.114 ;
    END
  END csrZCalCompVrefDAC[4]
  PIN csrZCalCompVrefDAC[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.22192 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 227.757 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 71.25 0 71.326 0.114 ;
    END
  END csrZCalCompVrefDAC[5]
  PIN csrZCalCompVrefDAC[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20368 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 212.574 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 71.858 0 71.934 0.114 ;
    END
  END csrZCalCompVrefDAC[6]
  PIN PwrOkVDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3155 LAYER M6 ;
    ANTENNADIFFAREA 0.02048 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.010112 LAYER M6 ;
      ANTENNAMAXAREACAR 2300.39 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 43.149 20.27 81.78 20.77 ;
    END
  END PwrOkVDD
  PIN VrefDacRef
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 243.375 LAYER M6 ;
    ANTENNADIFFAREA 11.2202 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 0 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 43.149 13.27 81.78 13.77 ;
        RECT 43.149 15.27 81.78 15.77 ;
        RECT 43.149 17.27 81.78 17.77 ;
        RECT 43.149 23.27 81.78 23.77 ;
        RECT 43.149 25.27 81.78 25.77 ;
        RECT 43.149 27.27 81.78 27.77 ;
        RECT 43.149 31.27 81.78 31.77 ;
        RECT 43.149 35.27 81.78 35.77 ;
        RECT 43.149 37.253 81.78 37.703 ;
        RECT 43.149 39.32 81.78 39.77 ;
        RECT 43.149 41.295 81.78 41.745 ;
        RECT 43.149 43.095 81.78 43.545 ;
    END
  END VrefDacRef
  PIN ZCalAnaClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1862 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 618.466 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 6.65 0 6.726 0.114 ;
    END
  END ZCalAnaClk
  PIN ZCalCompOut
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7083199375 LAYER M5 ;
    ANTENNADIFFAREA 0.030968 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 5.282 0 5.358 0.114 ;
    END
  END ZCalCompOut
  PIN csrZCalCompGainResAdj
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.14972 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 33.402 0 33.478 0.114 ;
    END
  END csrZCalCompGainResAdj
  PIN csrZCalCompBiasBypassEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.14972 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 33.25 0 33.326 0.114 ;
    END
  END csrZCalCompBiasBypassEn
  PIN csrZCalCompBiasPowerUp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.14972 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 33.098 0 33.174 0.114 ;
    END
  END csrZCalCompBiasPowerUp
  PIN csrZCalCompGainCurrAdj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0679059375 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 748.27 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 35.378 0 35.454 0.114 ;
    END
  END csrZCalCompGainCurrAdj[4]
  PIN csrZCalCompGainCurrAdj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07372 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001216 LAYER M5 ;
      ANTENNAMAXAREACAR 725.387 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 35.682 0 35.758 0.114 ;
    END
  END csrZCalCompGainCurrAdj[5]
  PIN csrZCalCompGainCurrAdj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07372 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 35.834 0 35.91 0.114 ;
    END
  END csrZCalCompGainCurrAdj[6]
  PIN csrZCalCompGainCurrAdj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07372 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 35.986 0 36.062 0.114 ;
    END
  END csrZCalCompGainCurrAdj[7]
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.3 70.875 81.78 71.325 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 72.675 81.78 73.125 ;
        RECT 0.3 74.475 81.78 74.925 ;
        RECT 0.3 76.275 81.78 76.725 ;
        RECT 0.3 78.075 81.78 78.525 ;
        RECT 0.3 79.875 81.78 80.325 ;
        RECT 0.3 81.675 81.78 82.125 ;
        RECT 0.3 83.475 81.78 83.925 ;
        RECT 0.3 85.275 81.78 85.725 ;
        RECT 0.3 87.075 81.78 87.525 ;
        RECT 0.3 88.875 81.78 89.325 ;
    END
  END VDDQ
  PIN ZCalDACRangeSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18544 LAYER M5 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M5 ;
      ANTENNAMAXAREACAR 495.368 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 73.226 0 73.302 0.114 ;
    END
  END ZCalDACRangeSel
  OBS
    LAYER M1 ;
      
      RECT MASK 1 0 0 82.08 90 ;
    
  
      RECT MASK 2 0 0 82.08 90 ;
    LAYER M2 ;
      RECT MASK 1 0 0 82.08 90 ;
   
      RECT MASK 2 0 0 82.08 90 ;
    LAYER M3 ;
      RECT MASK 1 0 0 82.08 90 ;
    LAYER M4 ;
      POLYGON 82.08 0 82.08 47.228 81.48 47.228 81.48 48.028 82.08 48.028 82.08 90 0 90 0 0 ;
    LAYER M3 ;
      RECT MASK 2 0 0 82.08 90 ;
    LAYER M4 ;
      RECT 80.406 47.428 81.48 47.828 ;
      RECT 35.446 50.276 80.706 50.676 ;
      RECT 5.5705 50.283 8.9545 50.669 ;
      RECT 31.58 52.76 37.902 53.151 ;
      RECT 6.0345 52.76 12.343 53.151 ;
      RECT 34.3935 53.517 38.9535 53.942 ;
      RECT 4.982 53.517 9.542 53.942 ;
      RECT 34.906 55.857 38.442 56.282 ;
      RECT 5.4945 55.857 9.0305 56.282 ;
      RECT 34.3935 58.227 38.9535 58.652 ;
      RECT 4.982 58.227 9.542 58.652 ;
      RECT 34.3935 52.078 38.9535 52.503 ;
      RECT 4.982 52.078 9.542 52.503 ;
      RECT 34.906 54.418 38.442 54.843 ;
      RECT 5.4945 54.418 9.0305 54.843 ;
      RECT 34.3935 56.788 38.9535 57.213 ;
      RECT 4.982 56.788 9.542 57.213 ;
    LAYER M5 ;
      POLYGON 82.08 0 82.08 90 0 90 0 0 5.206 0 5.206 0.19 5.434 0.19 5.434 0 6.574 0 6.574 0.19 6.802 0.19 6.802 0 33.022 0 33.022 0.19 33.554 0.19 33.554 0 34.39 0 34.39 0.19 34.922 0.19 34.922 0 34.998 0 34.998 0.19 35.53 0.19 35.53 0 35.606 0 35.606 0.19 36.138 0.19 36.138 0 45.182 0 45.182 0.19 45.714 0.19 45.714 0 69.198 0 69.198 0.19 69.73 0.19 69.73 0 69.806 0 69.806 0.19 70.338 0.19 70.338 0 70.414 0 70.414 0.19 70.946 0.19 70.946 0 71.022 0 71.022 0.19 71.554 0.19 71.554 0 71.782 0 71.782 0.19 72.162 0.19 72.162 0 73.15 0 73.15 0.19 73.378 0.19 73.378 0 ;
      RECT 5.869 2.99 5.949 14.36 ;
      RECT 22.989 17 23.069 28.6 ;
      RECT 37.2735 49.57 37.5135 58.652 ;
      RECT 36.3135 49.57 36.5535 58.652 ;
      RECT 35.3535 49.57 35.5935 58.652 ;
      RECT 37.7535 49.5775 37.9935 58.652 ;
      RECT 36.7935 49.5775 37.0335 58.652 ;
      RECT 35.8335 49.5775 36.0735 58.652 ;
      RECT 34.8735 49.5775 35.1135 58.652 ;
    LAYER M6 ;
      RECT 0.3 3.27 81.78 3.77 ;
      RECT 0.3 4.27 81.78 4.77 ;
      RECT 0.3 5.27 81.78 5.77 ;
      RECT 0.3 20.269 42.589 20.77 ;
      RECT 43.149 21.27 81.78 21.77 ;
      RECT 0.3 21.27 42.589 21.77 ;
      RECT 27.4915 31.95 32.1175 32.13 ;
      RECT 22.6055 31.95 27.2315 32.13 ;
      RECT 16.8075 31.95 21.4335 32.13 ;
      RECT 11.9215 31.95 16.5475 32.13 ;
      RECT 27.7065 32.26 32.1275 32.3 ;
      RECT 22.8205 32.26 27.2415 32.3 ;
      RECT 16.7975 32.26 21.2185 32.3 ;
      RECT 11.9115 32.26 16.3325 32.3 ;
      RECT 27.4815 32.34 31.9025 32.38 ;
      RECT 22.5955 32.34 27.0165 32.38 ;
      RECT 17.0225 32.34 21.4435 32.38 ;
      RECT 12.1365 32.34 16.5575 32.38 ;
      RECT 27.7065 32.42 32.1275 32.46 ;
      RECT 22.8205 32.42 27.2415 32.46 ;
      RECT 16.7975 32.42 21.2185 32.46 ;
      RECT 11.9115 32.42 16.3325 32.46 ;
      RECT 27.4815 32.5 31.9025 32.54 ;
      RECT 22.5955 32.5 27.0165 32.54 ;
      RECT 17.0225 32.5 21.4435 32.54 ;
      RECT 12.1365 32.5 16.5575 32.54 ;
      RECT 27.7065 32.58 32.1275 32.62 ;
      RECT 22.8205 32.58 27.2415 32.62 ;
      RECT 16.7975 32.58 21.2185 32.62 ;
      RECT 11.9115 32.58 16.3325 32.62 ;
      RECT 27.4815 32.66 31.9025 32.7 ;
      RECT 22.5955 32.66 27.0165 32.7 ;
      RECT 17.0225 32.66 21.4435 32.7 ;
      RECT 12.1365 32.66 16.5575 32.7 ;
      RECT 27.7065 32.74 32.1275 32.78 ;
      RECT 22.8205 32.74 27.2415 32.78 ;
      RECT 16.7975 32.74 21.2185 32.78 ;
      RECT 11.9115 32.74 16.3325 32.78 ;
      RECT 27.4815 32.82 31.9025 32.86 ;
      RECT 22.5955 32.82 27.0165 32.86 ;
      RECT 17.0225 32.82 21.4435 32.86 ;
      RECT 12.1365 32.82 16.5575 32.86 ;
      RECT 27.7065 32.9 32.1275 32.94 ;
      RECT 22.8205 32.9 27.2415 32.94 ;
      RECT 16.7975 32.9 21.2185 32.94 ;
      RECT 11.9115 32.9 16.3325 32.94 ;
      RECT 27.4815 32.98 31.9025 33.02 ;
      RECT 22.5955 32.98 27.0165 33.02 ;
      RECT 17.0225 32.98 21.4435 33.02 ;
      RECT 12.1365 32.98 16.5575 33.02 ;
      RECT 27.7065 33.06 32.1275 33.1 ;
      RECT 22.8205 33.06 27.2415 33.1 ;
      RECT 16.7975 33.06 21.2185 33.1 ;
      RECT 11.9115 33.06 16.3325 33.1 ;
      RECT 27.4815 33.14 31.9025 33.18 ;
      RECT 22.5955 33.14 27.0165 33.18 ;
      RECT 17.0225 33.14 21.4435 33.18 ;
      RECT 12.1365 33.14 16.5575 33.18 ;
      RECT 27.7065 33.22 32.1275 33.26 ;
      RECT 22.8205 33.22 27.2415 33.26 ;
      RECT 16.7975 33.22 21.2185 33.26 ;
      RECT 11.9115 33.22 16.3325 33.26 ;
      RECT 27.4815 33.3 31.9025 33.34 ;
      RECT 22.5955 33.3 27.0165 33.34 ;
      RECT 17.0225 33.3 21.4435 33.34 ;
      RECT 12.1365 33.3 16.5575 33.34 ;
      RECT 27.7065 33.38 32.1275 33.42 ;
      RECT 22.8205 33.38 27.2415 33.42 ;
      RECT 16.7975 33.38 21.2185 33.42 ;
      RECT 11.9115 33.38 16.3325 33.42 ;
      RECT 27.4815 33.46 31.9025 33.5 ;
      RECT 22.5955 33.46 27.0165 33.5 ;
      RECT 17.0225 33.46 21.4435 33.5 ;
      RECT 12.1365 33.46 16.5575 33.5 ;
      RECT 27.7065 33.54 32.1275 33.58 ;
      RECT 22.8205 33.54 27.2415 33.58 ;
      RECT 16.7975 33.54 21.2185 33.58 ;
      RECT 11.9115 33.54 16.3325 33.58 ;
      RECT 27.4815 33.62 31.9025 33.66 ;
      RECT 22.5955 33.62 27.0165 33.66 ;
      RECT 17.0225 33.62 21.4435 33.66 ;
      RECT 12.1365 33.62 16.5575 33.66 ;
      RECT 27.7065 33.7 32.1275 33.74 ;
      RECT 22.8205 33.7 27.2415 33.74 ;
      RECT 16.7975 33.7 21.2185 33.74 ;
      RECT 11.9115 33.7 16.3325 33.74 ;
      RECT 27.4815 33.78 31.9025 33.82 ;
      RECT 22.5955 33.78 27.0165 33.82 ;
      RECT 17.0225 33.78 21.4435 33.82 ;
      RECT 12.1365 33.78 16.5575 33.82 ;
      RECT 27.7065 33.86 32.1275 33.9 ;
      RECT 22.8205 33.86 27.2415 33.9 ;
      RECT 16.7975 33.86 21.2185 33.9 ;
      RECT 11.9115 33.86 16.3325 33.9 ;
      RECT 27.4815 33.94 31.9025 33.98 ;
      RECT 22.5955 33.94 27.0165 33.98 ;
      RECT 17.0225 33.94 21.4435 33.98 ;
      RECT 12.1365 33.94 16.5575 33.98 ;
      RECT 27.7065 34.02 32.1275 34.06 ;
      RECT 22.8205 34.02 27.2415 34.06 ;
      RECT 16.7975 34.02 21.2185 34.06 ;
      RECT 11.9115 34.02 16.3325 34.06 ;
      RECT 27.4815 34.1 31.9025 34.14 ;
      RECT 22.5955 34.1 27.0165 34.14 ;
      RECT 17.0225 34.1 21.4435 34.14 ;
      RECT 12.1365 34.1 16.5575 34.14 ;
      RECT 27.7065 34.18 32.1275 34.22 ;
      RECT 22.8205 34.18 27.2415 34.22 ;
      RECT 16.7975 34.18 21.2185 34.22 ;
      RECT 11.9115 34.18 16.3325 34.22 ;
      RECT 27.4815 34.26 31.9025 34.3 ;
      RECT 22.5955 34.26 27.0165 34.3 ;
      RECT 17.0225 34.26 21.4435 34.3 ;
      RECT 12.1365 34.26 16.5575 34.3 ;
      RECT 27.7065 34.34 32.1275 34.38 ;
      RECT 22.8205 34.34 27.2415 34.38 ;
      RECT 16.7975 34.34 21.2185 34.38 ;
      RECT 11.9115 34.34 16.3325 34.38 ;
      RECT 27.4815 34.42 31.9025 34.46 ;
      RECT 22.5955 34.42 27.0165 34.46 ;
      RECT 17.0225 34.42 21.4435 34.46 ;
      RECT 12.1365 34.42 16.5575 34.46 ;
      RECT 27.7065 34.5 32.1275 34.54 ;
      RECT 22.8205 34.5 27.2415 34.54 ;
      RECT 16.7975 34.5 21.2185 34.54 ;
      RECT 11.9115 34.5 16.3325 34.54 ;
      RECT 27.4815 34.58 31.9025 34.62 ;
      RECT 22.5955 34.58 27.0165 34.62 ;
      RECT 17.0225 34.58 21.4435 34.62 ;
      RECT 12.1365 34.58 16.5575 34.62 ;
      RECT 27.7065 34.66 32.1275 34.7 ;
      RECT 22.8205 34.66 27.2415 34.7 ;
      RECT 16.7975 34.66 21.2185 34.7 ;
      RECT 11.9115 34.66 16.3325 34.7 ;
      RECT 27.4815 34.74 31.9025 34.78 ;
      RECT 22.5955 34.74 27.0165 34.78 ;
      RECT 17.0225 34.74 21.4435 34.78 ;
      RECT 12.1365 34.74 16.5575 34.78 ;
      RECT 27.7065 34.82 32.1275 34.86 ;
      RECT 22.8205 34.82 27.2415 34.86 ;
      RECT 16.7975 34.82 21.2185 34.86 ;
      RECT 11.9115 34.82 16.3325 34.86 ;
      RECT 27.4815 34.9 31.9025 34.94 ;
      RECT 22.5955 34.9 27.0165 34.94 ;
      RECT 17.0225 34.9 21.4435 34.94 ;
      RECT 12.1365 34.9 16.5575 34.94 ;
      RECT 27.7065 34.98 32.1275 35.02 ;
      RECT 22.8205 34.98 27.2415 35.02 ;
      RECT 16.7975 34.98 21.2185 35.02 ;
      RECT 11.9115 34.98 16.3325 35.02 ;
      RECT 27.4815 35.06 31.9025 35.1 ;
      RECT 22.5955 35.06 27.0165 35.1 ;
      RECT 17.0225 35.06 21.4435 35.1 ;
      RECT 12.1365 35.06 16.5575 35.1 ;
      RECT 27.7065 35.14 32.1275 35.18 ;
      RECT 22.8205 35.14 27.2415 35.18 ;
      RECT 16.7975 35.14 21.2185 35.18 ;
      RECT 11.9115 35.14 16.3325 35.18 ;
      RECT 27.4815 35.22 31.9025 35.26 ;
      RECT 22.5955 35.22 27.0165 35.26 ;
      RECT 17.0225 35.22 21.4435 35.26 ;
      RECT 12.1365 35.22 16.5575 35.26 ;
      RECT 27.7065 35.3 32.1275 35.34 ;
      RECT 22.8205 35.3 27.2415 35.34 ;
      RECT 16.7975 35.3 21.2185 35.34 ;
      RECT 11.9115 35.3 16.3325 35.34 ;
      RECT 27.4815 35.38 31.9025 35.42 ;
      RECT 22.5955 35.38 27.0165 35.42 ;
      RECT 17.0225 35.38 21.4435 35.42 ;
      RECT 12.1365 35.38 16.5575 35.42 ;
      RECT 27.7065 35.46 32.1275 35.5 ;
      RECT 22.8205 35.46 27.2415 35.5 ;
      RECT 16.7975 35.46 21.2185 35.5 ;
      RECT 11.9115 35.46 16.3325 35.5 ;
      RECT 27.4815 35.54 31.9025 35.58 ;
      RECT 22.5955 35.54 27.0165 35.58 ;
      RECT 17.0225 35.54 21.4435 35.58 ;
      RECT 12.1365 35.54 16.5575 35.58 ;
      RECT 27.7065 35.62 32.1275 35.66 ;
      RECT 22.8205 35.62 27.2415 35.66 ;
      RECT 16.7975 35.62 21.2185 35.66 ;
      RECT 11.9115 35.62 16.3325 35.66 ;
      RECT 27.4815 35.7 31.9025 35.74 ;
      RECT 22.5955 35.7 27.0165 35.74 ;
      RECT 17.0225 35.7 21.4435 35.74 ;
      RECT 12.1365 35.7 16.5575 35.74 ;
      RECT 27.7065 35.78 32.1275 35.82 ;
      RECT 22.8205 35.78 27.2415 35.82 ;
      RECT 16.7975 35.78 21.2185 35.82 ;
      RECT 11.9115 35.78 16.3325 35.82 ;
      RECT 27.4815 35.86 31.9025 35.9 ;
      RECT 22.5955 35.86 27.0165 35.9 ;
      RECT 17.0225 35.86 21.4435 35.9 ;
      RECT 12.1365 35.86 16.5575 35.9 ;
      RECT 27.7065 35.94 32.1275 35.98 ;
      RECT 22.8205 35.94 27.2415 35.98 ;
      RECT 16.7975 35.94 21.2185 35.98 ;
      RECT 11.9115 35.94 16.3325 35.98 ;
      RECT 27.4815 36.02 31.9025 36.06 ;
      RECT 22.5955 36.02 27.0165 36.06 ;
      RECT 17.0225 36.02 21.4435 36.06 ;
      RECT 12.1365 36.02 16.5575 36.06 ;
      RECT 27.7065 36.1 32.1275 36.14 ;
      RECT 22.8205 36.1 27.2415 36.14 ;
      RECT 16.7975 36.1 21.2185 36.14 ;
      RECT 11.9115 36.1 16.3325 36.14 ;
      RECT 27.4915 36.27 32.1175 36.45 ;
      RECT 22.6055 36.27 27.2315 36.45 ;
      RECT 16.8075 36.27 21.4335 36.45 ;
      RECT 11.9215 36.27 16.5475 36.45 ;
      RECT 27.4915 39.39 32.1175 39.57 ;
      RECT 22.6055 39.39 27.2315 39.57 ;
      RECT 16.8075 39.39 21.4335 39.57 ;
      RECT 11.9215 39.39 16.5475 39.57 ;
      RECT 27.7065 39.7 32.1275 39.74 ;
      RECT 22.8205 39.7 27.2415 39.74 ;
      RECT 16.7975 39.7 21.2185 39.74 ;
      RECT 11.9115 39.7 16.3325 39.74 ;
      RECT 27.4815 39.78 31.9025 39.82 ;
      RECT 22.5955 39.78 27.0165 39.82 ;
      RECT 17.0225 39.78 21.4435 39.82 ;
      RECT 12.1365 39.78 16.5575 39.82 ;
      RECT 27.7065 39.86 32.1275 39.9 ;
      RECT 22.8205 39.86 27.2415 39.9 ;
      RECT 16.7975 39.86 21.2185 39.9 ;
      RECT 11.9115 39.86 16.3325 39.9 ;
      RECT 27.4815 39.94 31.9025 39.98 ;
      RECT 22.5955 39.94 27.0165 39.98 ;
      RECT 17.0225 39.94 21.4435 39.98 ;
      RECT 12.1365 39.94 16.5575 39.98 ;
      RECT 27.7065 40.02 32.1275 40.06 ;
      RECT 22.8205 40.02 27.2415 40.06 ;
      RECT 16.7975 40.02 21.2185 40.06 ;
      RECT 11.9115 40.02 16.3325 40.06 ;
      RECT 27.4815 40.1 31.9025 40.14 ;
      RECT 22.5955 40.1 27.0165 40.14 ;
      RECT 17.0225 40.1 21.4435 40.14 ;
      RECT 12.1365 40.1 16.5575 40.14 ;
      RECT 27.7065 40.18 32.1275 40.22 ;
      RECT 22.8205 40.18 27.2415 40.22 ;
      RECT 16.7975 40.18 21.2185 40.22 ;
      RECT 11.9115 40.18 16.3325 40.22 ;
      RECT 27.4815 40.26 31.9025 40.3 ;
      RECT 22.5955 40.26 27.0165 40.3 ;
      RECT 17.0225 40.26 21.4435 40.3 ;
      RECT 12.1365 40.26 16.5575 40.3 ;
      RECT 27.7065 40.34 32.1275 40.38 ;
      RECT 22.8205 40.34 27.2415 40.38 ;
      RECT 16.7975 40.34 21.2185 40.38 ;
      RECT 11.9115 40.34 16.3325 40.38 ;
      RECT 27.4815 40.42 31.9025 40.46 ;
      RECT 22.5955 40.42 27.0165 40.46 ;
      RECT 17.0225 40.42 21.4435 40.46 ;
      RECT 12.1365 40.42 16.5575 40.46 ;
      RECT 27.7065 40.5 32.1275 40.54 ;
      RECT 22.8205 40.5 27.2415 40.54 ;
      RECT 16.7975 40.5 21.2185 40.54 ;
      RECT 11.9115 40.5 16.3325 40.54 ;
      RECT 27.4815 40.58 31.9025 40.62 ;
      RECT 22.5955 40.58 27.0165 40.62 ;
      RECT 17.0225 40.58 21.4435 40.62 ;
      RECT 12.1365 40.58 16.5575 40.62 ;
      RECT 27.7065 40.66 32.1275 40.7 ;
      RECT 22.8205 40.66 27.2415 40.7 ;
      RECT 16.7975 40.66 21.2185 40.7 ;
      RECT 11.9115 40.66 16.3325 40.7 ;
      RECT 27.4815 40.74 31.9025 40.78 ;
      RECT 22.5955 40.74 27.0165 40.78 ;
      RECT 17.0225 40.74 21.4435 40.78 ;
      RECT 12.1365 40.74 16.5575 40.78 ;
      RECT 27.7065 40.82 32.1275 40.86 ;
      RECT 22.8205 40.82 27.2415 40.86 ;
      RECT 16.7975 40.82 21.2185 40.86 ;
      RECT 11.9115 40.82 16.3325 40.86 ;
      RECT 27.4815 40.9 31.9025 40.94 ;
      RECT 22.5955 40.9 27.0165 40.94 ;
      RECT 17.0225 40.9 21.4435 40.94 ;
      RECT 12.1365 40.9 16.5575 40.94 ;
      RECT 27.7065 40.98 32.1275 41.02 ;
      RECT 22.8205 40.98 27.2415 41.02 ;
      RECT 16.7975 40.98 21.2185 41.02 ;
      RECT 11.9115 40.98 16.3325 41.02 ;
      RECT 27.4815 41.06 31.9025 41.1 ;
      RECT 22.5955 41.06 27.0165 41.1 ;
      RECT 17.0225 41.06 21.4435 41.1 ;
      RECT 12.1365 41.06 16.5575 41.1 ;
      RECT 27.7065 41.14 32.1275 41.18 ;
      RECT 22.8205 41.14 27.2415 41.18 ;
      RECT 16.7975 41.14 21.2185 41.18 ;
      RECT 11.9115 41.14 16.3325 41.18 ;
      RECT 27.4815 41.22 31.9025 41.26 ;
      RECT 22.5955 41.22 27.0165 41.26 ;
      RECT 17.0225 41.22 21.4435 41.26 ;
      RECT 12.1365 41.22 16.5575 41.26 ;
      RECT 27.7065 41.3 32.1275 41.34 ;
      RECT 22.8205 41.3 27.2415 41.34 ;
      RECT 16.7975 41.3 21.2185 41.34 ;
      RECT 11.9115 41.3 16.3325 41.34 ;
      RECT 27.4815 41.38 31.9025 41.42 ;
      RECT 22.5955 41.38 27.0165 41.42 ;
      RECT 17.0225 41.38 21.4435 41.42 ;
      RECT 12.1365 41.38 16.5575 41.42 ;
      RECT 27.7065 41.46 32.1275 41.5 ;
      RECT 22.8205 41.46 27.2415 41.5 ;
      RECT 16.7975 41.46 21.2185 41.5 ;
      RECT 11.9115 41.46 16.3325 41.5 ;
      RECT 27.4815 41.54 31.9025 41.58 ;
      RECT 22.5955 41.54 27.0165 41.58 ;
      RECT 17.0225 41.54 21.4435 41.58 ;
      RECT 12.1365 41.54 16.5575 41.58 ;
      RECT 27.7065 41.62 32.1275 41.66 ;
      RECT 22.8205 41.62 27.2415 41.66 ;
      RECT 16.7975 41.62 21.2185 41.66 ;
      RECT 11.9115 41.62 16.3325 41.66 ;
      RECT 27.4815 41.7 31.9025 41.74 ;
      RECT 22.5955 41.7 27.0165 41.74 ;
      RECT 17.0225 41.7 21.4435 41.74 ;
      RECT 12.1365 41.7 16.5575 41.74 ;
      RECT 27.7065 41.78 32.1275 41.82 ;
      RECT 22.8205 41.78 27.2415 41.82 ;
      RECT 16.7975 41.78 21.2185 41.82 ;
      RECT 11.9115 41.78 16.3325 41.82 ;
      RECT 27.4815 41.86 31.9025 41.9 ;
      RECT 22.5955 41.86 27.0165 41.9 ;
      RECT 17.0225 41.86 21.4435 41.9 ;
      RECT 12.1365 41.86 16.5575 41.9 ;
      RECT 27.7065 41.94 32.1275 41.98 ;
      RECT 22.8205 41.94 27.2415 41.98 ;
      RECT 16.7975 41.94 21.2185 41.98 ;
      RECT 11.9115 41.94 16.3325 41.98 ;
      RECT 27.4815 42.02 31.9025 42.06 ;
      RECT 22.5955 42.02 27.0165 42.06 ;
      RECT 17.0225 42.02 21.4435 42.06 ;
      RECT 12.1365 42.02 16.5575 42.06 ;
      RECT 27.7065 42.1 32.1275 42.14 ;
      RECT 22.8205 42.1 27.2415 42.14 ;
      RECT 16.7975 42.1 21.2185 42.14 ;
      RECT 11.9115 42.1 16.3325 42.14 ;
      RECT 27.4815 42.18 31.9025 42.22 ;
      RECT 22.5955 42.18 27.0165 42.22 ;
      RECT 17.0225 42.18 21.4435 42.22 ;
      RECT 12.1365 42.18 16.5575 42.22 ;
      RECT 27.7065 42.26 32.1275 42.3 ;
      RECT 22.8205 42.26 27.2415 42.3 ;
      RECT 16.7975 42.26 21.2185 42.3 ;
      RECT 11.9115 42.26 16.3325 42.3 ;
      RECT 27.4815 42.34 31.9025 42.38 ;
      RECT 22.5955 42.34 27.0165 42.38 ;
      RECT 17.0225 42.34 21.4435 42.38 ;
      RECT 12.1365 42.34 16.5575 42.38 ;
      RECT 27.7065 42.42 32.1275 42.46 ;
      RECT 22.8205 42.42 27.2415 42.46 ;
      RECT 16.7975 42.42 21.2185 42.46 ;
      RECT 11.9115 42.42 16.3325 42.46 ;
      RECT 27.4815 42.5 31.9025 42.54 ;
      RECT 22.5955 42.5 27.0165 42.54 ;
      RECT 17.0225 42.5 21.4435 42.54 ;
      RECT 12.1365 42.5 16.5575 42.54 ;
      RECT 27.7065 42.58 32.1275 42.62 ;
      RECT 22.8205 42.58 27.2415 42.62 ;
      RECT 16.7975 42.58 21.2185 42.62 ;
      RECT 11.9115 42.58 16.3325 42.62 ;
      RECT 27.4815 42.66 31.9025 42.7 ;
      RECT 22.5955 42.66 27.0165 42.7 ;
      RECT 17.0225 42.66 21.4435 42.7 ;
      RECT 12.1365 42.66 16.5575 42.7 ;
      RECT 27.7065 42.74 32.1275 42.78 ;
      RECT 22.8205 42.74 27.2415 42.78 ;
      RECT 16.7975 42.74 21.2185 42.78 ;
      RECT 11.9115 42.74 16.3325 42.78 ;
      RECT 27.4815 42.82 31.9025 42.86 ;
      RECT 22.5955 42.82 27.0165 42.86 ;
      RECT 17.0225 42.82 21.4435 42.86 ;
      RECT 12.1365 42.82 16.5575 42.86 ;
      RECT 27.7065 42.9 32.1275 42.94 ;
      RECT 22.8205 42.9 27.2415 42.94 ;
      RECT 16.7975 42.9 21.2185 42.94 ;
      RECT 11.9115 42.9 16.3325 42.94 ;
      RECT 27.4815 42.98 31.9025 43.02 ;
      RECT 22.5955 42.98 27.0165 43.02 ;
      RECT 17.0225 42.98 21.4435 43.02 ;
      RECT 12.1365 42.98 16.5575 43.02 ;
      RECT 27.7065 43.06 32.1275 43.1 ;
      RECT 22.8205 43.06 27.2415 43.1 ;
      RECT 16.7975 43.06 21.2185 43.1 ;
      RECT 11.9115 43.06 16.3325 43.1 ;
      RECT 27.4815 43.14 31.9025 43.18 ;
      RECT 22.5955 43.14 27.0165 43.18 ;
      RECT 17.0225 43.14 21.4435 43.18 ;
      RECT 12.1365 43.14 16.5575 43.18 ;
      RECT 27.7065 43.22 32.1275 43.26 ;
      RECT 22.8205 43.22 27.2415 43.26 ;
      RECT 16.7975 43.22 21.2185 43.26 ;
      RECT 11.9115 43.22 16.3325 43.26 ;
      RECT 27.4815 43.3 31.9025 43.34 ;
      RECT 22.5955 43.3 27.0165 43.34 ;
      RECT 17.0225 43.3 21.4435 43.34 ;
      RECT 12.1365 43.3 16.5575 43.34 ;
      RECT 27.7065 43.38 32.1275 43.42 ;
      RECT 22.8205 43.38 27.2415 43.42 ;
      RECT 16.7975 43.38 21.2185 43.42 ;
      RECT 11.9115 43.38 16.3325 43.42 ;
      RECT 27.4815 43.46 31.9025 43.5 ;
      RECT 22.5955 43.46 27.0165 43.5 ;
      RECT 17.0225 43.46 21.4435 43.5 ;
      RECT 12.1365 43.46 16.5575 43.5 ;
      RECT 27.7065 43.54 32.1275 43.58 ;
      RECT 22.8205 43.54 27.2415 43.58 ;
      RECT 16.7975 43.54 21.2185 43.58 ;
      RECT 11.9115 43.54 16.3325 43.58 ;
      RECT 27.4915 43.71 32.1175 43.89 ;
      RECT 22.6055 43.71 27.2315 43.89 ;
      RECT 16.8075 43.71 21.4335 43.89 ;
      RECT 11.9215 43.71 16.5475 43.89 ;
    LAYER M0 ;
      
      RECT MASK 1 0 0 82.08 90 ;
      RECT MASK 2 0 0 82.08 90 ;
  END
END dwc_ddrphy_zcalana

END LIBRARY
