# LEF OUT API 
# Creation Date : Thu Feb 24 23:22:12 IST 2022
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_lpddr5xphy_txrxdq_ew
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_lpddr5xphy_txrxdq_ew 0 0 ;
  SYMMETRY X Y ;
  SIZE 97.971 BY 37.38 ;
  PIN csrRxCurrAdj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.285665 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 194.55 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.641 0.038 2.679 ;
    END
  END csrRxCurrAdj[4]
  PIN csrRxCurrAdj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.288971 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 217.735 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.249 0.038 3.287 ;
    END
  END csrRxCurrAdj[3]
  PIN csrRxCurrAdj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.282226 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 439.065 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.033 0.038 2.071 ;
    END
  END csrRxCurrAdj[2]
  PIN csrRxCurrAdj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38873975 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 450.814 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.553 0.038 3.591 ;
    END
  END csrRxCurrAdj[1]
  PIN csrRxCurrAdj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.320188 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 399.763 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.705 0.038 3.743 ;
    END
  END csrRxCurrAdj[0]
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M10 ;
        RECT 50.637 17.831 78.672 18.431 ;
        RECT 50.637 16.031 78.672 16.631 ;
        RECT 50.637 14.231 78.672 14.831 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 26.1795 48.919 26.7795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 22.1795 48.919 22.7795 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 11.3465 78.672 11.9465 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 29.255 78.672 29.855 ;
        RECT 50.637 27.455 78.672 28.055 ;
        RECT 50.637 25.655 78.672 26.255 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 22.7705 78.672 23.3705 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 25.5895 87.277 26.1475 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 29.6215 87.277 30.1795 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 34.1945 78.672 34.7945 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 33.6535 87.277 34.2115 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 27.6055 88.673 28.1635 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 31.6375 88.673 32.1955 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 2.9765 48.919 3.5765 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 11.4775 88.673 12.0355 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 7.4455 88.673 8.0035 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 3.4135 88.673 3.9715 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 9.4615 87.277 10.0195 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 5.4295 87.277 5.9875 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 15.5095 88.673 16.0675 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 23.5735 88.673 24.1315 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 19.5415 88.673 20.0995 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 21.5575 87.277 22.1155 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 17.5255 87.277 18.0835 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 13.4935 87.277 14.0515 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 6.5365 48.919 7.1365 ;
    END
    PORT
      LAYER M10 ;
        RECT 79.335 2.4055 97.065 2.9635 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 29.7795 48.919 30.3795 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 6.407 78.672 7.007 ;
        RECT 50.637 4.607 78.672 5.207 ;
        RECT 50.637 2.807 78.672 3.407 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 1.1965 48.919 1.7965 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 4.7565 48.919 5.3565 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 20.3795 48.919 20.9795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 13.4165 48.919 14.0165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 11.3165 48.919 11.9165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 10.4165 48.919 11.0165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 27.9795 48.919 28.5795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 23.9795 48.919 24.5795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 17.099 26.941 17.699 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 8.6365 48.919 9.2365 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 35.6185 48.919 36.2185 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 33.8185 48.919 34.4185 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 31.5795 48.919 32.1795 ;
    END
  END VSS
  PIN VIO_PwrOk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4546 LAYER M10 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.21816 LAYER M10 ;
      ANTENNAMAXAREACAR 40.6162 LAYER M10 ;
    PORT
      LAYER M10 ;
        RECT 47.393 7.4365 51.484 8.0365 ;
    END
  END VIO_PwrOk
  PIN VIO_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.298 LAYER M10 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAMAXAREACAR 6.51602 LAYER M10 ;
    PORT
      LAYER M10 ;
        RECT 64.3825 30.9755 76.436 31.4255 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 26.6515 95.823 27.1015 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 28.6675 95.823 29.1175 ;
    END
    PORT
      LAYER M10 ;
        RECT 27.823 17.099 31.653 17.699 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 10.5235 95.823 10.9735 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 6.4915 95.823 6.9415 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 4.4755 95.823 4.9255 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 8.5075 95.823 8.9575 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 20.6035 95.823 21.0535 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 14.5555 95.823 15.0055 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 12.5395 95.823 12.9895 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 16.5715 95.823 17.0215 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 22.6195 95.823 23.0695 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 24.6355 95.823 25.0855 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 18.5875 95.823 19.0375 ;
    END
    PORT
      LAYER M10 ;
        RECT 64.3825 19.5515 76.436 20.0015 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 32.6995 95.823 33.1495 ;
    END
    PORT
      LAYER M10 ;
        RECT 80.577 30.6835 95.823 31.1335 ;
    END
    PORT
      LAYER M10 ;
        RECT 64.3825 8.1275 76.436 8.5775 ;
    END
  END VIO_PAD
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M10 ;
        RECT 79.335 34.6615 97.065 35.2195 ;
    END
    PORT
      LAYER M10 ;
        RECT 63.6785 35.0945 78.672 35.6945 ;
        RECT 63.6785 33.2945 78.672 33.8945 ;
        RECT 63.6785 23.6705 78.672 24.2705 ;
        RECT 63.6785 21.8705 78.672 22.4705 ;
        RECT 63.6785 12.2465 78.672 12.8465 ;
        RECT 63.6785 10.4465 78.672 11.0465 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.6375 28.355 78.6725 28.955 ;
        RECT 63.6785 26.555 78.672 27.155 ;
        RECT 63.6785 24.755 78.672 25.355 ;
    END
    PORT
      LAYER M10 ;
        RECT 89.123 31.6375 97.065 32.1955 ;
    END
    PORT
      LAYER M10 ;
        RECT 89.123 27.6055 97.065 28.1635 ;
    END
    PORT
      LAYER M10 ;
        RECT 87.727 25.5895 97.065 26.1475 ;
    END
    PORT
      LAYER M10 ;
        RECT 87.727 33.6535 97.065 34.2115 ;
    END
    PORT
      LAYER M10 ;
        RECT 33.928 34.7185 48.919 35.3185 ;
    END
    PORT
      LAYER M10 ;
        RECT 87.727 9.4615 97.065 10.0195 ;
    END
    PORT
      LAYER M10 ;
        RECT 87.727 5.4295 97.065 5.9875 ;
    END
    PORT
      LAYER M10 ;
        RECT 89.123 11.4775 97.065 12.0355 ;
    END
    PORT
      LAYER M10 ;
        RECT 89.123 7.4455 97.065 8.0035 ;
    END
    PORT
      LAYER M10 ;
        RECT 89.123 3.4135 97.065 3.9715 ;
    END
    PORT
      LAYER M10 ;
        RECT 87.727 17.5255 97.065 18.0835 ;
    END
    PORT
      LAYER M10 ;
        RECT 87.727 13.4935 97.065 14.0515 ;
    END
    PORT
      LAYER M10 ;
        RECT 87.727 21.5575 97.065 22.1155 ;
    END
    PORT
      LAYER M10 ;
        RECT 89.123 19.5415 97.065 20.0995 ;
    END
    PORT
      LAYER M10 ;
        RECT 89.123 23.5735 97.065 24.1315 ;
    END
    PORT
      LAYER M10 ;
        RECT 89.123 15.5095 97.065 16.0675 ;
    END
    PORT
      LAYER M10 ;
        RECT 87.727 29.6215 97.065 30.1795 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.6375 5.507 78.6725 6.107 ;
        RECT 63.6785 3.707 78.672 4.307 ;
        RECT 63.6785 1.907 78.672 2.507 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.6375 16.931 78.6725 17.531 ;
        RECT 63.6785 15.131 78.672 15.731 ;
        RECT 63.6785 13.331 78.672 13.931 ;
    END
    PORT
      LAYER M10 ;
        RECT 33.928 3.8765 48.919 4.4765 ;
    END
    PORT
      LAYER M10 ;
        RECT 33.928 2.1075 48.919 2.7075 ;
    END
    PORT
      LAYER M10 ;
        RECT 33.928 5.6565 48.919 6.2565 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M10 ;
        RECT 50.637 12.2465 63.1455 12.8465 ;
        RECT 50.637 10.4465 63.1455 11.0465 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 26.555 63.1455 27.155 ;
        RECT 50.637 24.755 63.1455 25.355 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 23.6705 63.1455 24.2705 ;
        RECT 50.637 21.8705 63.1455 22.4705 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 35.0945 63.1455 35.6945 ;
        RECT 50.637 33.2945 63.1455 33.8945 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 3.707 63.1455 4.307 ;
        RECT 50.637 1.907 63.1455 2.507 ;
    END
    PORT
      LAYER M10 ;
        RECT 50.637 15.131 63.1455 15.731 ;
        RECT 50.637 13.331 63.1455 13.931 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 34.7185 33.328 35.3185 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 30.6795 48.919 31.2795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 28.8795 48.919 29.4795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 25.2795 48.919 25.8795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 14.3165 48.919 14.9165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 5.6565 33.328 6.2565 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 32.7795 48.919 33.3795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 27.0795 48.919 27.6795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 23.0795 48.919 23.6795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 21.2795 48.919 21.8795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 19.1795 48.919 19.7795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 17.999 48.919 18.599 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 16.199 48.919 16.799 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 15.2165 48.919 15.8165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 12.2165 48.919 12.8165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 9.5365 48.919 10.1365 ;
        RECT 0.3 7.4365 46.793 8.0365 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 3.8765 33.328 4.4765 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 2.0965 33.328 2.6965 ;
    END
  END VDD
  PIN RxStandBy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.285931 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 386.576 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.969 0.038 1.007 ;
    END
  END RxStandBy
  PIN RxPowerDown
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.28234 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 389.245 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.665 0.038 0.703 ;
    END
  END RxPowerDown
  PIN RxFwdClkT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.351823 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 20.653 0.038 20.691 ;
    END
  END RxFwdClkT
  PIN RxFwdClkC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.352165 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 15.485 0.038 15.523 ;
    END
  END RxFwdClkC
  PIN RxDataOdd
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.347738 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 15.561 0.038 15.599 ;
    END
  END RxDataOdd
  PIN RxDataEven
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.351823 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 21.261 0.038 21.299 ;
    END
  END RxDataEven
  PIN RxDFEInit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.296001 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 361.236 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 5.529 0.038 5.567 ;
    END
  END RxDFEInit
  PIN RxClkT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.46933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03444 LAYER M6 ;
      ANTENNAMAXAREACAR 104.649 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 21.109 0.038 21.147 ;
    END
  END RxClkT
  PIN RxClkC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.46933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03444 LAYER M6 ;
      ANTENNAMAXAREACAR 113.796 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 15.713 0.038 15.751 ;
    END
  END RxClkC
  PIN RxBypassRcvEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.263739 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 127.745 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.525 0.038 18.563 ;
    END
  END RxBypassRcvEn
  PIN RxBypassPadEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.28667175 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 397.137 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 5.073 0.038 5.111 ;
    END
  END RxBypassPadEn
  PIN RxBypassDataPad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.447602 LAYER M6 ;
    ANTENNADIFFAREA 0.00918 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 11.837 0.038 11.875 ;
    END
  END RxBypassDataPad
  PIN RxBypassData[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.351823 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 20.957 0.038 20.995 ;
    END
  END RxBypassData[1]
  PIN RxBypassData[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.284943 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 15.789 0.038 15.827 ;
    END
  END RxBypassData[0]
  PIN Pclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.282169 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 189.961 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 6.593 0.038 6.631 ;
    END
  END Pclk
  PIN IDDQ_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.25957775 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06222 LAYER M6 ;
      ANTENNAMAXAREACAR 60.0531 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.829 0.038 18.867 ;
    END
  END IDDQ_mode
  PIN PwrOkVDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.44522 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0132 LAYER M7 ;
      ANTENNAMAXAREACAR 1032.5899998 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 48.507 0.05 48.545 37.33 ;
    END
  END PwrOkVDD
  PIN TxClkDcdSampleClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.303544 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 211.148 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 30.001 0.038 30.039 ;
    END
  END TxClkDcdSampleClk
  PIN TxClkDcdOut
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.309453 LAYER M6 ;
    ANTENNADIFFAREA 0.01836 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 29.697 0.038 29.735 ;
    END
  END TxClkDcdOut
  PIN csrTxClkDcdOffset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.311714 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 183.575 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 29.545 0.038 29.583 ;
    END
  END csrTxClkDcdOffset[0]
  PIN csrTxClkDcdOffset[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267368 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 180.327 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 30.153 0.038 30.191 ;
    END
  END csrTxClkDcdOffset[1]
  PIN csrTxClkDcdOffset[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.277305 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 179.135 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 29.849 0.038 29.887 ;
    END
  END csrTxClkDcdOffset[3]
  PIN csrTxClkDcdOffset[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27322 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 176.373 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 30.305 0.038 30.343 ;
    END
  END csrTxClkDcdOffset[2]
  PIN csrTxClkDcdMode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.318383 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 192.041 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 29.089 0.038 29.127 ;
    END
  END csrTxClkDcdMode[0]
  PIN csrTxClkDcdMode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.30584275 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 192.884 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 29.393 0.038 29.431 ;
    END
  END csrTxClkDcdMode[1]
  PIN csrTxClkDcdOffset[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.304114 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 173.115 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 29.241 0.038 29.279 ;
    END
  END csrTxClkDcdOffset[4]
  PIN csrRxVrefDac[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 657.527 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.917 0.038 36.955 ;
    END
  END csrRxVrefDac[3]
  PIN csrRxVrefDac[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 452.109 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.689 0.038 36.727 ;
    END
  END csrRxVrefDac[0]
  PIN csrRxVrefDac[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 684.374 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.993 0.038 37.031 ;
    END
  END csrRxVrefDac[4]
  PIN csrRxVrefDac[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 690.916 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 37.145 0.038 37.183 ;
    END
  END csrRxVrefDac[6]
  PIN csrRxVrefDac[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 446.827 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.765 0.038 36.803 ;
    END
  END csrRxVrefDac[1]
  PIN csrRxVrefDac[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 661.555 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.841 0.038 36.879 ;
    END
  END csrRxVrefDac[2]
  PIN csrRxVrefDac[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 424.218 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.613 0.038 36.651 ;
    END
  END csrRxVrefDac[8]
  PIN csrRxVrefDac[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 441.886 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 37.221 0.038 37.259 ;
    END
  END csrRxVrefDac[7]
  PIN csrRxVrefDac[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49804 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M6 ;
      ANTENNAMAXAREACAR 690.087 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 37.069 0.038 37.107 ;
    END
  END csrRxVrefDac[5]
  PIN csrLsTxCalCodePD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 483.062 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.723 0.05 49.761 37.33 ;
    END
  END csrLsTxCalCodePD[2]
  PIN csrLsTxCalCodePD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 492.014 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.647 0.05 49.685 37.33 ;
    END
  END csrLsTxCalCodePD[1]
  PIN csrLsTxCalCodePD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 503.15 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.571 0.05 49.609 37.33 ;
    END
  END csrLsTxCalCodePD[0]
  PIN csrLsTxSlewLPPU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 324.068 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 48.887 0.05 48.925 37.33 ;
    END
  END csrLsTxSlewLPPU[0]
  PIN csrLsTxSlewPD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 313.061 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.191 0.05 49.229 37.33 ;
    END
  END csrLsTxSlewPD[2]
  PIN BurnIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0.026068 LAYER M7 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAGATEAREA 0.00204 LAYER M7 ;
      ANTENNAGATEAREA 0.00102 LAYER VIA6 ;
      ANTENNAMAXAREACAR 151.921 LAYER M6 ;
      ANTENNAMAXAREACAR 407.648 LAYER M7 ;
      ANTENNAMAXCUTCAR 5.92158 LAYER VIA6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.781 0.038 3.819 ;
    END
  END BurnIn
  PIN csrLsTxCalCodePD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 475.128 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.799 0.05 49.837 37.33 ;
    END
  END csrLsTxCalCodePD[3]
  PIN csrLsTxCalCodePD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 468.695 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.875 0.05 49.913 37.33 ;
    END
  END csrLsTxCalCodePD[4]
  PIN csrLsTxCalCodePD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 461.94 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.951 0.05 49.989 37.33 ;
    END
  END csrLsTxCalCodePD[5]
  PIN csrLsTxCalCodePD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 429.749 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.027 0.05 50.065 37.33 ;
    END
  END csrLsTxCalCodePD[6]
  PIN csrLsTxCalCodePD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 450.303 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.103 0.05 50.141 37.33 ;
    END
  END csrLsTxCalCodePD[7]
  PIN csrLsTxCalCodePD[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 437.299 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.179 0.05 50.217 37.33 ;
    END
  END csrLsTxCalCodePD[8]
  PIN csrLsTxCalCodeLPPU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 485.647 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.255 0.05 50.293 37.33 ;
    END
  END csrLsTxCalCodeLPPU[0]
  PIN csrLsTxCalCodeLPPU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 468.125 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.407 0.05 50.445 37.33 ;
    END
  END csrLsTxCalCodeLPPU[2]
  PIN csrLsTxCalCodeLPPU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 465.284 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.331 0.05 50.369 37.33 ;
    END
  END csrLsTxCalCodeLPPU[1]
  PIN csrLsTxCalCodeLPPU[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 456.238 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.483 0.05 50.521 37.33 ;
    END
  END csrLsTxCalCodeLPPU[3]
  PIN csrLsTxCalCodeLPPU[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 431.632 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.559 0.05 50.597 37.33 ;
    END
  END csrLsTxCalCodeLPPU[4]
  PIN csrLsTxCalCodeLPPU[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 430.815 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.635 0.05 50.673 37.33 ;
    END
  END csrLsTxCalCodeLPPU[5]
  PIN csrLsTxCalCodeLPPU[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 401.525 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.711 0.05 50.749 37.33 ;
    END
  END csrLsTxCalCodeLPPU[6]
  PIN csrLsTxCalCodeLPPU[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 388.23 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.787 0.05 50.825 37.33 ;
    END
  END csrLsTxCalCodeLPPU[7]
  PIN csrLsTxCalCodeLPPU[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 375.148 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 50.863 0.05 50.901 37.33 ;
    END
  END csrLsTxCalCodeLPPU[8]
  PIN csrLsTxSlewPD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 310.9 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.115 0.05 49.153 37.33 ;
    END
  END csrLsTxSlewPD[1]
  PIN csrLsTxSlewLPPU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 359.473 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 48.811 0.05 48.849 37.33 ;
    END
  END csrLsTxSlewLPPU[2]
  PIN csrLsTxSlewLPPU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 317.177 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 48.963 0.05 49.001 37.33 ;
    END
  END csrLsTxSlewLPPU[1]
  PIN csrLsTxSlewPD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 314.937 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.039 0.05 49.077 37.33 ;
    END
  END csrLsTxSlewPD[0]
  PIN csrLsTxSlewPD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 334.647 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 49.267 0.05 49.305 37.33 ;
    END
  END csrLsTxSlewPD[3]
  PIN scan_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.283271 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.05201975 LAYER M6 ;
      ANTENNAMAXAREACAR 488.558 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 11.685 0.038 11.723 ;
    END
  END scan_mode
  PIN csrTxSeg120PU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 91.5509 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 4.389 0.038 4.427 ;
    END
  END csrTxSeg120PU[2]
  PIN csrTxSeg120PU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 85.5019 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 30.989 0.038 31.027 ;
    END
  END csrTxSeg120PU[1]
  PIN csrTxSeg120PU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.8774 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.877 0.038 33.915 ;
    END
  END csrTxSeg120PU[0]
  PIN csrTxSeg120PD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024529 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.1897 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 6.213 0.038 6.251 ;
    END
  END csrTxSeg120PD[2]
  PIN csrTxSeg120PD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.8632 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 32.585 0.038 32.623 ;
    END
  END csrTxSeg120PD[1]
  PIN csrTxSeg120PD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 92.5245 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.473 0.038 35.511 ;
    END
  END csrTxSeg120PD[0]
  PIN csrTxDcaMode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.159353 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 209.134 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 11.533 0.038 11.571 ;
    END
  END csrTxDcaMode
  PIN csrTxDcaFinePU[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 85.19929975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.021 0.033 3.059 ;
    END
  END csrTxDcaFinePU[3]
  PIN csrTxDcaFinePU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 137.038 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.717 0.033 2.755 ;
    END
  END csrTxDcaFinePU[2]
  PIN csrTxDcaFinePU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 113.297 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.413 0.033 2.451 ;
    END
  END csrTxDcaFinePU[1]
  PIN csrTxDcaFinePU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 85.9592 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.261 0.033 2.299 ;
    END
  END csrTxDcaFinePU[0]
  PIN csrTxDcaFinePD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 82.3451 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.197 0.034 1.235 ;
    END
  END csrTxDcaFinePD[3]
  PIN csrTxDcaFinePD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 179.17 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.501 0.034 1.539 ;
    END
  END csrTxDcaFinePD[2]
  PIN csrTxDcaFinePD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 126.295 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.653 0.034 1.691 ;
    END
  END csrTxDcaFinePD[1]
  PIN csrTxDcaFinePD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 75.8058 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.957 0.034 1.995 ;
    END
  END csrTxDcaFinePD[0]
  PIN csrTxDcaCoarse[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 116.091 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.173 0.033 3.211 ;
    END
  END csrTxDcaCoarse[1]
  PIN csrTxDcaCoarse[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 125.773 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.477 0.033 3.515 ;
    END
  END csrTxDcaCoarse[0]
  PIN csrOdtSeg120PU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 96.6108 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.933 0.038 3.971 ;
    END
  END csrOdtSeg120PU[2]
  PIN csrOdtSeg120PU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 98.2799 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 31.217 0.038 31.255 ;
    END
  END csrOdtSeg120PU[1]
  PIN csrOdtSeg120PU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 101.721 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 34.257 0.038 34.295 ;
    END
  END csrOdtSeg120PU[0]
  PIN csrOdtSeg120PD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.1059 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 6.061 0.038 6.099 ;
    END
  END csrOdtSeg120PD[2]
  PIN csrOdtSeg120PD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 97.7667 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 32.889 0.038 32.927 ;
    END
  END csrOdtSeg120PD[1]
  PIN csrOdtSeg120PD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 100.681 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.853 0.038 35.891 ;
    END
  END csrOdtSeg120PD[0]
  PIN csrCoreLoopBackMode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0051 LAYER M6 ;
      ANTENNAMAXAREACAR 127.561 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 15.941 0.038 15.979 ;
    END
  END csrCoreLoopBackMode
  PIN csrRxOffsetSelOdd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.282568 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 123.986 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 8.113 0.038 8.151 ;
    END
  END csrRxOffsetSelOdd[2]
  PIN csrRxOffsetSelOdd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.28425875 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 131.656 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 8.569 0.038 8.607 ;
    END
  END csrRxOffsetSelOdd[3]
  PIN TxOEOdd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026619 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00867 LAYER M6 ;
      ANTENNAMAXAREACAR 34.4283 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 17.081 0.038 17.119 ;
    END
  END TxOEOdd
  PIN TxOEEven
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034789 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00867 LAYER M6 ;
      ANTENNAMAXAREACAR 34.0927 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 16.777 0.038 16.815 ;
    END
  END TxOEEven
  PIN TxFwdClk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.029564 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.905 0.038 18.943 ;
    END
  END TxFwdClk
  PIN TxDataOdd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026182 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 82.7265 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 20.729 0.038 20.767 ;
    END
  END TxDataOdd
  PIN TxDataEven
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034808 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 65.25889975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 20.273 0.038 20.311 ;
    END
  END TxDataEven
  PIN csrRxOffsetSelOdd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.282853 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 133.249 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 8.265 0.038 8.303 ;
    END
  END csrRxOffsetSelOdd[4]
  PIN scan_shift
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286729 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0204 LAYER M6 ;
      ANTENNAMAXAREACAR 25.2499 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.857 0.038 3.895 ;
    END
  END scan_shift
  PIN TxClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.078014 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.01533 LAYER M6 ;
      ANTENNAMAXAREACAR 12.7818 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 22.933 0.038 22.971 ;
    END
  END TxClk
  PIN TxBypassOEInt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.027949 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 364.115 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.297 0.038 18.335 ;
    END
  END TxBypassOEInt
  PIN TxBypassOEExt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022781 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 377.175 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 19.969 0.038 20.007 ;
    END
  END TxBypassOEExt
  PIN TxBypassModeInt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026619 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 195.885 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.069 0.038 18.107 ;
    END
  END TxBypassModeInt
  PIN TxBypassModeExt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034998 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 134.881 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.981 0.038 19.019 ;
    END
  END TxBypassModeExt
  PIN TxBypassDataInt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.025156 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 324.389 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 19.741 0.038 19.779 ;
    END
  END TxBypassDataInt
  PIN TxBypassDataExt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024282 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 327.172 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 19.361 0.038 19.399 ;
    END
  END TxBypassDataExt
  PIN scan_shift_cg
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289598 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 364.145 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 5.985 0.038 6.023 ;
    END
  END scan_shift_cg
  PIN scan_si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286729 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 441.872 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 4.161 0.038 4.199 ;
    END
  END scan_si
  PIN OdtEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022952 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 105.397 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.449 0.038 18.487 ;
    END
  END OdtEn
  PIN scan_so
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.38402775 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 7.657 0.038 7.695 ;
    END
  END scan_so
  PIN csrRxOffsetSelOdd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.295526 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 133.766 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 7.353 0.038 7.391 ;
    END
  END csrRxOffsetSelOdd[1]
  PIN csrRxOffsetSelOdd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.282302 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 140.801 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 7.961 0.038 7.999 ;
    END
  END csrRxOffsetSelOdd[0]
  PIN csrRxOffsetSelEven[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.28524675 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 135.091 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 9.329 0.038 9.367 ;
    END
  END csrRxOffsetSelEven[4]
  PIN csrRxOffsetSelEven[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286596 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 129.887 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 9.481 0.038 9.519 ;
    END
  END csrRxOffsetSelEven[3]
  PIN csrRxOffsetSelEven[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.285228 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 125.012 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 9.177 0.038 9.215 ;
    END
  END csrRxOffsetSelEven[2]
  PIN csrRxOffsetSelEven[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.29953475 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 134.867 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 8.417 0.038 8.455 ;
    END
  END csrRxOffsetSelEven[1]
  PIN csrRxOffsetSelEven[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.283404 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 145.422 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 9.025 0.038 9.063 ;
    END
  END csrRxOffsetSelEven[0]
  PIN csrRxOffsetEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.282891 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 400.048 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 6.897 0.038 6.935 ;
    END
  END csrRxOffsetEn
  PIN csrRxModeCtl[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.40582075 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 476.609 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.285 0.038 0.323 ;
    END
  END csrRxModeCtl[3]
  PIN csrRxModeCtl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.408082 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 469.433 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.361 0.038 0.399 ;
    END
  END csrRxModeCtl[2]
  PIN csrRxModeCtl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.40582075 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 457.168 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.437 0.038 0.475 ;
    END
  END csrRxModeCtl[1]
  PIN csrRxModeCtl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.389671 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 228.186 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.513 0.038 0.551 ;
    END
  END csrRxModeCtl[0]
  PIN csrRxGainCtrl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.388056 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 222.198 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.185 0.038 2.223 ;
    END
  END csrRxGainCtrl[2]
  PIN csrRxGainCtrl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.441522 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 260.91699975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.881 0.038 1.919 ;
    END
  END csrRxGainCtrl[1]
  PIN csrRxGainCtrl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.281979 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 227.033 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.273 0.038 1.311 ;
    END
  END csrRxGainCtrl[0]
  PIN csrRxDFETap2Sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.302062 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 182.608 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 4.921 0.038 4.959 ;
    END
  END csrRxDFETap2Sel[4]
  PIN csrRxDFETap2Sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.284525 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 241.198 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.121 0.038 1.159 ;
    END
  END csrRxDFETap2Sel[3]
  PIN csrRxDFETap2Sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286881 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 181.877 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 5.377 0.038 5.415 ;
    END
  END csrRxDFETap2Sel[2]
  PIN csrRxDFETap2Sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.297768 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 188.724 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 4.465 0.038 4.503 ;
    END
  END csrRxDFETap2Sel[1]
  PIN csrRxDFETap2Sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286881 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 191.593 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 5.225 0.038 5.263 ;
    END
  END csrRxDFETap2Sel[0]
  PIN csrRxDFETap1Sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.28348 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 183.676 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 4.009 0.038 4.047 ;
    END
  END csrRxDFETap1Sel[4]
  PIN csrRxDFETap1Sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.282226 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 196.36 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.401 0.038 3.439 ;
    END
  END csrRxDFETap1Sel[3]
  PIN csrRxDFETap1Sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286767 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 215.547 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.793 0.038 2.831 ;
    END
  END csrRxDFETap1Sel[2]
  PIN csrRxDFETap1Sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.308218 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 227.866 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.489 0.038 2.527 ;
    END
  END csrRxDFETap1Sel[1]
  PIN csrRxDFETap1Sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.29241 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 225.445 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.337 0.038 2.375 ;
    END
  END csrRxDFETap1Sel[0]
  PIN csrRxDFECtrl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.286881 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 249.904 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 4.617 0.038 4.655 ;
    END
  END csrRxDFECtrl[2]
  PIN csrRxDFECtrl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.405194 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 231.557 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.893 0.038 0.931 ;
    END
  END csrRxDFECtrl[1]
  PIN csrRxDFECtrl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.298091 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 152.612 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.741 0.038 0.779 ;
    END
  END csrRxDFECtrl[0]
  PIN csrRxDFEBiasSel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.294481 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 376.53 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 5.681 0.038 5.719 ;
    END
  END csrRxDFEBiasSel[1]
  PIN csrRxDFEBiasSel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289104 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 352.063 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 5.833 0.038 5.871 ;
    END
  END csrRxDFEBiasSel[0]
  PIN csrRxCurrAdj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.373046 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 522.866 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 4.769 0.038 4.807 ;
    END
  END csrRxCurrAdj[7]
  PIN csrRxCurrAdj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.28270075 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 206.124 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.945 0.038 2.983 ;
    END
  END csrRxCurrAdj[6]
  PIN csrRxCurrAdj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.299763 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 197.412 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.097 0.038 3.135 ;
    END
  END csrRxCurrAdj[5]
  OBS
    LAYER M0 SPACING 0 ;
      RECT MASK 1 0 0 97.971 37.38 ;
    LAYER M0 SPACING 0 ;
      RECT MASK 2 0 0 97.971 37.38 ;
    LAYER M1 SPACING 0 ;
      RECT MASK 1 0 0 97.971 37.38 ;
    LAYER M1 SPACING 0 ;
      RECT MASK 2 0 0 97.971 37.38 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 1 0 0 97.971 37.38 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 2 0 0 97.971 37.38 ;
    LAYER M3 SPACING 0 ;
      RECT MASK 1 0 0 97.971 37.38 ;
    LAYER M4 SPACING 0 ;
      RECT MASK 1 0 0 97.971 37.38 ;
    LAYER M5 SPACING 0 ;
      RECT 0 0 97.971 37.38 ;
    LAYER M3 SPACING 0 ;
      RECT MASK 2 0 0 97.971 37.38 ;
    LAYER M4 SPACING 0 ;
      RECT MASK 2 0 0 97.971 37.38 ;
    LAYER M6 SPACING 0 ;
      POLYGON 97.971 0 97.971 37.38 0 37.38 0 37.259 0.038 37.259 0.038 37.221 0 37.221 0 37.183 0.038 37.183 0.038 37.145 0 37.145 0 37.107 0.038 37.107 0.038 37.069 0 37.069 0 37.031 0.038 37.031 0.038 36.993 0 36.993 0 36.955 0.038 36.955 0.038 36.917 0 36.917 0 36.879 0.038 36.879 0.038 36.841 0 36.841 0 36.803 0.038 36.803 0.038 36.765 0 36.765 0 36.727 0.038 36.727 0.038 36.689 0 36.689 0 36.651 0.038 36.651 0.038 36.613 0 36.613 0 35.891 0.038 35.891 0.038 35.853 0 35.853 0 35.511 0.038 35.511 0.038 35.473 0 35.473 0 34.295 0.038 34.295 0.038 34.257 0 34.257 0 33.915 0.038 33.915 0.038 33.877 0 33.877 0 32.927 0.038 32.927 0.038 32.889 0 32.889 0 32.623 0.038 32.623 0.038 32.585 0 32.585 0 31.255 0.038 31.255 0.038 31.217 0 31.217 0 31.027 0.038 31.027 0.038 30.989 0 30.989 0 30.343 0.038 30.343 0.038 30.305 0 30.305 0 30.191 0.038 30.191 0.038 30.153 0 30.153 0 30.039 0.038 30.039 0.038 30.001 0 30.001 0 29.887 0.038 29.887 0.038 29.849 0 29.849 0 29.735 0.038 29.735 0.038 29.697 0 29.697 0 29.583 0.038 29.583 0.038 29.545 0 29.545 0 29.431 0.038 29.431 0.038 29.393 0 29.393 0 29.279 0.038 29.279 0.038 29.241 0 29.241 0 29.127 0.038 29.127 0.038 29.089 0 29.089 0 22.971 0.038 22.971 0.038 22.933 0 22.933 0 21.299 0.038 21.299 0.038 21.261 0 21.261 0 21.147 0.038 21.147 0.038 21.109 0 21.109 0 20.995 0.038 20.995 0.038 20.957 0 20.957 0 20.767 0.038 20.767 0.038 20.729 0 20.729 0 20.691 0.038 20.691 0.038 20.653 0 20.653 0 20.311 0.038 20.311 0.038 20.273 0 20.273 0 20.007 0.038 20.007 0.038 19.969 0 19.969 0 19.779 0.038 19.779 0.038 19.741 0 19.741 0 19.399 0.038 19.399 0.038 19.361 0 19.361 0 19.019 0.038 19.019 0.038 18.981 0 18.981 0 18.943 0.038 18.943 0.038 18.905 0 18.905 0 18.867 0.038 18.867 0.038 18.829 0 18.829 0 18.563 0.038 18.563 0.038 18.525 0 18.525 0 18.487 0.038 18.487 0.038 18.449 0 18.449 0 18.335 0.038 18.335 0.038 18.297 0 18.297 0 18.107 0.038 18.107 0.038 18.069 0 18.069 0 17.119 0.038 17.119 0.038 17.081 0 17.081 0 16.815 0.038 16.815 0.038 16.777 0 16.777 0 15.979 0.038 15.979 0.038 15.941 0 15.941 0 15.827 0.038 15.827 0.038 15.789 0 15.789 0 15.751 0.038 15.751 0.038 15.713 0 15.713 0 15.599 0.038 15.599 0.038 15.561 0 15.561 0 15.523 0.038 15.523 0.038 15.485 0 15.485 0 11.875 0.038 11.875 0.038 11.837 0 11.837 0 11.723 0.038 11.723 0.038 11.685 0 11.685 0 11.571 0.038 11.571 0.038 11.533 0 11.533 0 9.519 0.038 9.519 0.038 9.481 0 9.481 0 9.367 0.038 9.367 0.038 9.329 0 9.329 0 9.215 0.038 9.215 0.038 9.177 0 9.177 0 9.063 0.038 9.063 0.038 9.025 0 9.025 0 8.607 0.038 8.607 0.038 8.569 0 8.569 0 8.455 0.038 8.455 0.038 8.417 0 8.417 0 8.303 0.038 8.303 0.038 8.265 0 8.265 0 8.151 0.038 8.151 0.038 8.113 0 8.113 0 7.999 0.038 7.999 0.038 7.961 0 7.961 0 7.695 0.038 7.695 0.038 7.657 0 7.657 0 7.391 0.038 7.391 0.038 7.353 0 7.353 0 6.935 0.038 6.935 0.038 6.897 0 6.897 0 6.631 0.038 6.631 0.038 6.593 0 6.593 0 6.251 0.038 6.251 0.038 6.213 0 6.213 0 6.099 0.038 6.099 0.038 6.061 0 6.061 0 6.023 0.038 6.023 0.038 5.985 0 5.985 0 5.871 0.038 5.871 0.038 5.833 0 5.833 0 5.719 0.038 5.719 0.038 5.681 0 5.681 0 5.567 0.038 5.567 0.038 5.529 0 5.529 0 5.415 0.038 5.415 0.038 5.377 0 5.377 0 5.263 0.038 5.263 0.038 5.225 0 5.225 0 5.111 0.038 5.111 0.038 5.073 0 5.073 0 4.959 0.038 4.959 0.038 4.921 0 4.921 0 4.807 0.038 4.807 0.038 4.769 0 4.769 0 4.655 0.038 4.655 0.038 4.617 0 4.617 0 4.503 0.038 4.503 0.038 4.465 0 4.465 0 4.427 0.038 4.427 0.038 4.389 0 4.389 0 4.199 0.038 4.199 0.038 4.161 0 4.161 0 4.047 0.038 4.047 0.038 4.009 0 4.009 0 3.971 0.038 3.971 0.038 3.933 0 3.933 0 3.895 0.038 3.895 0.038 3.857 0 3.857 0 3.819 0.038 3.819 0.038 3.781 0 3.781 0 3.743 0.038 3.743 0.038 3.705 0 3.705 0 3.591 0.038 3.591 0.038 3.553 0 3.553 0 3.515 0.033 3.515 0.033 3.477 0 3.477 0 3.439 0.038 3.439 0.038 3.401 0 3.401 0 3.287 0.038 3.287 0.038 3.249 0 3.249 0 3.211 0.033 3.211 0.033 3.173 0 3.173 0 3.135 0.038 3.135 0.038 3.097 0 3.097 0 3.059 0.033 3.059 0.033 3.021 0 3.021 0 2.983 0.038 2.983 0.038 2.945 0 2.945 0 2.831 0.038 2.831 0.038 2.793 0 2.793 0 2.755 0.033 2.755 0.033 2.717 0 2.717 0 2.679 0.038 2.679 0.038 2.641 0 2.641 0 2.527 0.038 2.527 0.038 2.489 0 2.489 0 2.451 0.033 2.451 0.033 2.413 0 2.413 0 2.375 0.038 2.375 0.038 2.337 0 2.337 0 2.299 0.033 2.299 0.033 2.261 0 2.261 0 2.223 0.038 2.223 0.038 2.185 0 2.185 0 2.071 0.038 2.071 0.038 2.033 0 2.033 0 1.995 0.034 1.995 0.034 1.957 0 1.957 0 1.919 0.038 1.919 0.038 1.881 0 1.881 0 1.691 0.034 1.691 0.034 1.653 0 1.653 0 1.539 0.034 1.539 0.034 1.501 0 1.501 0 1.311 0.038 1.311 0.038 1.273 0 1.273 0 1.235 0.034 1.235 0.034 1.197 0 1.197 0 1.159 0.038 1.159 0.038 1.121 0 1.121 0 1.007 0.038 1.007 0.038 0.969 0 0.969 0 0.931 0.038 0.931 0.038 0.893 0 0.893 0 0.779 0.038 0.779 0.038 0.741 0 0.741 0 0.703 0.038 0.703 0.038 0.665 0 0.665 0 0.551 0.038 0.551 0.038 0.513 0 0.513 0 0.475 0.038 0.475 0.038 0.437 0 0.437 0 0.399 0.038 0.399 0.038 0.361 0 0.361 0 0.323 0.038 0.323 0.038 0.285 0 0.285 0 0 ;
    LAYER M7 SPACING 0 ;
      POLYGON 0 0 0 37.38 97.971 37.38 97.971 37.33 48.507 37.33 48.507 0.05 48.545 0.05 48.545 37.33 48.811 37.33 48.811 0.05 48.849 0.05 48.849 37.33 48.887 37.33 48.887 0.05 48.925 0.05 48.925 37.33 48.963 37.33 48.963 0.05 49.001 0.05 49.001 37.33 49.039 37.33 49.039 0.05 49.077 0.05 49.077 37.33 49.115 37.33 49.115 0.05 49.153 0.05 49.153 37.33 49.191 37.33 49.191 0.05 49.229 0.05 49.229 37.33 49.267 37.33 49.267 0.05 49.305 0.05 49.305 37.33 49.571 37.33 49.571 0.05 49.609 0.05 49.609 37.33 49.647 37.33 49.647 0.05 49.685 0.05 49.685 37.33 49.723 37.33 49.723 0.05 49.761 0.05 49.761 37.33 49.799 37.33 49.799 0.05 49.837 0.05 49.837 37.33 49.875 37.33 49.875 0.05 49.913 0.05 49.913 37.33 49.951 37.33 49.951 0.05 49.989 0.05 49.989 37.33 50.027 37.33 50.027 0.05 50.065 0.05 50.065 37.33 50.103 37.33 50.103 0.05 50.141 0.05 50.141 37.33 50.179 37.33 50.179 0.05 50.217 0.05 50.217 37.33 50.255 37.33 50.255 0.05 50.293 0.05 50.293 37.33 50.331 37.33 50.331 0.05 50.369 0.05 50.369 37.33 50.407 37.33 50.407 0.05 50.445 0.05 50.445 37.33 50.483 37.33 50.483 0.05 50.521 0.05 50.521 37.33 50.559 37.33 50.559 0.05 50.597 0.05 50.597 37.33 50.635 37.33 50.635 0.05 50.673 0.05 50.673 37.33 50.711 37.33 50.711 0.05 50.749 0.05 50.749 37.33 50.787 37.33 50.787 0.05 50.825 0.05 50.825 37.33 50.863 37.33 50.863 0.05 50.901 0.05 50.901 37.33 97.971 37.33 97.971 0 ;
    LAYER M8 SPACING 0 ;
      RECT 0 0 97.971 37.38 ;
    LAYER M9 SPACING 0 ;
      RECT 0 0 97.971 37.38 ;
    LAYER M10 SPACING 0 ;
      POLYGON 0 0 0 37.38 97.971 37.38 97.971 36.2185 0.3 36.2185 0.3 35.6185 48.919 35.6185 48.919 36.2185 97.971 36.2185 97.971 35.6945 50.637 35.6945 50.637 35.3185 0.3 35.3185 0.3 34.7185 33.328 34.7185 33.328 35.3185 33.928 35.3185 33.928 34.7185 48.919 34.7185 48.919 35.3185 50.637 35.3185 50.637 35.0945 63.1455 35.0945 63.1455 35.6945 63.6785 35.6945 63.6785 35.0945 78.672 35.0945 78.672 35.6945 97.971 35.6945 97.971 35.2195 79.335 35.2195 79.335 34.7945 50.637 34.7945 50.637 34.4185 0.3 34.4185 0.3 33.8185 48.919 33.8185 48.919 34.4185 50.637 34.4185 50.637 34.1945 78.672 34.1945 78.672 34.7945 79.335 34.7945 79.335 34.6615 97.065 34.6615 97.065 35.2195 97.971 35.2195 97.971 34.2115 79.335 34.2115 79.335 33.8945 50.637 33.8945 50.637 33.3795 0.3 33.3795 0.3 32.7795 48.919 32.7795 48.919 33.3795 50.637 33.3795 50.637 33.2945 63.1455 33.2945 63.1455 33.8945 63.6785 33.8945 63.6785 33.2945 78.672 33.2945 78.672 33.8945 79.335 33.8945 79.335 33.6535 87.277 33.6535 87.277 34.2115 87.727 34.2115 87.727 33.6535 97.065 33.6535 97.065 34.2115 97.971 34.2115 97.971 33.1495 80.577 33.1495 80.577 32.6995 95.823 32.6995 95.823 33.1495 97.971 33.1495 97.971 32.1955 79.335 32.1955 79.335 32.1795 0.3 32.1795 0.3 31.5795 48.919 31.5795 48.919 32.1795 79.335 32.1795 79.335 31.6375 88.673 31.6375 88.673 32.1955 89.123 32.1955 89.123 31.6375 97.065 31.6375 97.065 32.1955 97.971 32.1955 97.971 31.4255 64.3825 31.4255 64.3825 31.2795 0.3 31.2795 0.3 30.6795 48.919 30.6795 48.919 31.2795 64.3825 31.2795 64.3825 30.9755 76.436 30.9755 76.436 31.4255 97.971 31.4255 97.971 31.1335 80.577 31.1335 80.577 30.6835 95.823 30.6835 95.823 31.1335 97.971 31.1335 97.971 30.3795 0.3 30.3795 0.3 29.7795 48.919 29.7795 48.919 30.3795 97.971 30.3795 97.971 30.1795 79.335 30.1795 79.335 29.855 50.637 29.855 50.637 29.4795 0.3 29.4795 0.3 28.8795 48.919 28.8795 48.919 29.4795 50.637 29.4795 50.637 29.255 78.672 29.255 78.672 29.855 79.335 29.855 79.335 29.6215 87.277 29.6215 87.277 30.1795 87.727 30.1795 87.727 29.6215 97.065 29.6215 97.065 30.1795 97.971 30.1795 97.971 29.1175 80.577 29.1175 80.577 28.955 50.6375 28.955 50.6375 28.5795 0.3 28.5795 0.3 27.9795 48.919 27.9795 48.919 28.5795 50.6375 28.5795 50.6375 28.355 78.6725 28.355 78.6725 28.955 80.577 28.955 80.577 28.6675 95.823 28.6675 95.823 29.1175 97.971 29.1175 97.971 28.1635 79.335 28.1635 79.335 28.055 50.637 28.055 50.637 27.6795 0.3 27.6795 0.3 27.0795 48.919 27.0795 48.919 27.6795 50.637 27.6795 50.637 27.455 78.672 27.455 78.672 28.055 79.335 28.055 79.335 27.6055 88.673 27.6055 88.673 28.1635 89.123 28.1635 89.123 27.6055 97.065 27.6055 97.065 28.1635 97.971 28.1635 97.971 27.155 50.637 27.155 50.637 26.7795 0.3 26.7795 0.3 26.1795 48.919 26.1795 48.919 26.7795 50.637 26.7795 50.637 26.555 63.1455 26.555 63.1455 27.155 63.6785 27.155 63.6785 26.555 78.672 26.555 78.672 27.155 97.971 27.155 97.971 27.1015 80.577 27.1015 80.577 26.6515 95.823 26.6515 95.823 27.1015 97.971 27.1015 97.971 26.255 50.637 26.255 50.637 25.8795 0.3 25.8795 0.3 25.2795 48.919 25.2795 48.919 25.8795 50.637 25.8795 50.637 25.655 78.672 25.655 78.672 26.255 97.971 26.255 97.971 26.1475 79.335 26.1475 79.335 25.5895 87.277 25.5895 87.277 26.1475 87.727 26.1475 87.727 25.5895 97.065 25.5895 97.065 26.1475 97.971 26.1475 97.971 25.355 50.637 25.355 50.637 24.755 63.1455 24.755 63.1455 25.355 63.6785 25.355 63.6785 24.755 78.672 24.755 78.672 25.355 97.971 25.355 97.971 25.0855 80.577 25.0855 80.577 24.6355 95.823 24.6355 95.823 25.0855 97.971 25.0855 97.971 24.5795 0.3 24.5795 0.3 23.9795 48.919 23.9795 48.919 24.5795 97.971 24.5795 97.971 24.2705 50.637 24.2705 50.637 23.6795 0.3 23.6795 0.3 23.0795 48.919 23.0795 48.919 23.6795 50.637 23.6795 50.637 23.6705 63.1455 23.6705 63.1455 24.2705 63.6785 24.2705 63.6785 23.6705 78.672 23.6705 78.672 24.2705 97.971 24.2705 97.971 24.1315 79.335 24.1315 79.335 23.5735 88.673 23.5735 88.673 24.1315 89.123 24.1315 89.123 23.5735 97.065 23.5735 97.065 24.1315 97.971 24.1315 97.971 23.3705 50.637 23.3705 50.637 22.7795 0.3 22.7795 0.3 22.1795 48.919 22.1795 48.919 22.7795 50.637 22.7795 50.637 22.7705 78.672 22.7705 78.672 23.3705 97.971 23.3705 97.971 23.0695 80.577 23.0695 80.577 22.6195 95.823 22.6195 95.823 23.0695 97.971 23.0695 97.971 22.4705 50.637 22.4705 50.637 21.8795 0.3 21.8795 0.3 21.2795 48.919 21.2795 48.919 21.8795 50.637 21.8795 50.637 21.8705 63.1455 21.8705 63.1455 22.4705 63.6785 22.4705 63.6785 21.8705 78.672 21.8705 78.672 22.4705 97.971 22.4705 97.971 22.1155 79.335 22.1155 79.335 21.5575 87.277 21.5575 87.277 22.1155 87.727 22.1155 87.727 21.5575 97.065 21.5575 97.065 22.1155 97.971 22.1155 97.971 21.0535 80.577 21.0535 80.577 20.9795 0.3 20.9795 0.3 20.3795 48.919 20.3795 48.919 20.9795 80.577 20.9795 80.577 20.6035 95.823 20.6035 95.823 21.0535 97.971 21.0535 97.971 20.0995 79.335 20.0995 79.335 20.0015 64.3825 20.0015 64.3825 19.7795 0.3 19.7795 0.3 19.1795 48.919 19.1795 48.919 19.7795 64.3825 19.7795 64.3825 19.5515 76.436 19.5515 76.436 20.0015 79.335 20.0015 79.335 19.5415 88.673 19.5415 88.673 20.0995 89.123 20.0995 89.123 19.5415 97.065 19.5415 97.065 20.0995 97.971 20.0995 97.971 19.0375 80.577 19.0375 80.577 18.599 0.3 18.599 0.3 17.999 48.919 17.999 48.919 18.599 80.577 18.599 80.577 18.5875 95.823 18.5875 95.823 19.0375 97.971 19.0375 97.971 18.431 50.637 18.431 50.637 17.831 78.672 17.831 78.672 18.431 97.971 18.431 97.971 18.0835 79.335 18.0835 79.335 17.699 0.3 17.699 0.3 17.099 26.941 17.099 26.941 17.699 27.823 17.699 27.823 17.099 31.653 17.099 31.653 17.699 79.335 17.699 79.335 17.531 50.6375 17.531 50.6375 16.931 78.6725 16.931 78.6725 17.531 79.335 17.531 79.335 17.5255 87.277 17.5255 87.277 18.0835 87.727 18.0835 87.727 17.5255 97.065 17.5255 97.065 18.0835 97.971 18.0835 97.971 17.0215 80.577 17.0215 80.577 16.799 0.3 16.799 0.3 16.199 48.919 16.199 48.919 16.799 80.577 16.799 80.577 16.631 50.637 16.631 50.637 16.031 78.672 16.031 78.672 16.631 80.577 16.631 80.577 16.5715 95.823 16.5715 95.823 17.0215 97.971 17.0215 97.971 16.0675 79.335 16.0675 79.335 15.8165 0.3 15.8165 0.3 15.2165 48.919 15.2165 48.919 15.8165 79.335 15.8165 79.335 15.731 50.637 15.731 50.637 15.131 63.1455 15.131 63.1455 15.731 63.6785 15.731 63.6785 15.131 78.672 15.131 78.672 15.731 79.335 15.731 79.335 15.5095 88.673 15.5095 88.673 16.0675 89.123 16.0675 89.123 15.5095 97.065 15.5095 97.065 16.0675 97.971 16.0675 97.971 15.0055 80.577 15.0055 80.577 14.9165 0.3 14.9165 0.3 14.3165 48.919 14.3165 48.919 14.9165 80.577 14.9165 80.577 14.831 50.637 14.831 50.637 14.231 78.672 14.231 78.672 14.831 80.577 14.831 80.577 14.5555 95.823 14.5555 95.823 15.0055 97.971 15.0055 97.971 14.0515 79.335 14.0515 79.335 14.0165 0.3 14.0165 0.3 13.4165 48.919 13.4165 48.919 14.0165 79.335 14.0165 79.335 13.931 50.637 13.931 50.637 13.331 63.1455 13.331 63.1455 13.931 63.6785 13.931 63.6785 13.331 78.672 13.331 78.672 13.931 79.335 13.931 79.335 13.4935 87.277 13.4935 87.277 14.0515 87.727 14.0515 87.727 13.4935 97.065 13.4935 97.065 14.0515 97.971 14.0515 97.971 12.9895 80.577 12.9895 80.577 12.8465 50.637 12.8465 50.637 12.8165 0.3 12.8165 0.3 12.2165 48.919 12.2165 48.919 12.8165 50.637 12.8165 50.637 12.2465 63.1455 12.2465 63.1455 12.8465 63.6785 12.8465 63.6785 12.2465 78.672 12.2465 78.672 12.8465 80.577 12.8465 80.577 12.5395 95.823 12.5395 95.823 12.9895 97.971 12.9895 97.971 12.0355 79.335 12.0355 79.335 11.9465 50.637 11.9465 50.637 11.9165 0.3 11.9165 0.3 11.3165 48.919 11.3165 48.919 11.9165 50.637 11.9165 50.637 11.3465 78.672 11.3465 78.672 11.9465 79.335 11.9465 79.335 11.4775 88.673 11.4775 88.673 12.0355 89.123 12.0355 89.123 11.4775 97.065 11.4775 97.065 12.0355 97.971 12.0355 97.971 11.0465 50.637 11.0465 50.637 11.0165 0.3 11.0165 0.3 10.4165 48.919 10.4165 48.919 11.0165 50.637 11.0165 50.637 10.4465 63.1455 10.4465 63.1455 11.0465 63.6785 11.0465 63.6785 10.4465 78.672 10.4465 78.672 11.0465 97.971 11.0465 97.971 10.9735 80.577 10.9735 80.577 10.5235 95.823 10.5235 95.823 10.9735 97.971 10.9735 97.971 10.1365 0.3 10.1365 0.3 9.5365 48.919 9.5365 48.919 10.1365 97.971 10.1365 97.971 10.0195 79.335 10.0195 79.335 9.4615 87.277 9.4615 87.277 10.0195 87.727 10.0195 87.727 9.4615 97.065 9.4615 97.065 10.0195 97.971 10.0195 97.971 9.2365 0.3 9.2365 0.3 8.6365 48.919 8.6365 48.919 9.2365 97.971 9.2365 97.971 8.9575 80.577 8.9575 80.577 8.5775 64.3825 8.5775 64.3825 8.1275 76.436 8.1275 76.436 8.5775 80.577 8.5775 80.577 8.5075 95.823 8.5075 95.823 8.9575 97.971 8.9575 97.971 8.0365 0.3 8.0365 0.3 7.4365 46.793 7.4365 46.793 8.0365 47.393 8.0365 47.393 7.4365 51.484 7.4365 51.484 8.0365 97.971 8.0365 97.971 8.0035 79.335 8.0035 79.335 7.4455 88.673 7.4455 88.673 8.0035 89.123 8.0035 89.123 7.4455 97.065 7.4455 97.065 8.0035 97.971 8.0035 97.971 7.1365 0.3 7.1365 0.3 6.5365 48.919 6.5365 48.919 7.1365 97.971 7.1365 97.971 7.007 50.637 7.007 50.637 6.407 78.672 6.407 78.672 7.007 97.971 7.007 97.971 6.9415 80.577 6.9415 80.577 6.4915 95.823 6.4915 95.823 6.9415 97.971 6.9415 97.971 6.2565 0.3 6.2565 0.3 5.6565 33.328 5.6565 33.328 6.2565 33.928 6.2565 33.928 5.6565 48.919 5.6565 48.919 6.2565 97.971 6.2565 97.971 6.107 50.6375 6.107 50.6375 5.507 78.6725 5.507 78.6725 6.107 97.971 6.107 97.971 5.9875 79.335 5.9875 79.335 5.4295 87.277 5.4295 87.277 5.9875 87.727 5.9875 87.727 5.4295 97.065 5.4295 97.065 5.9875 97.971 5.9875 97.971 5.3565 0.3 5.3565 0.3 4.7565 48.919 4.7565 48.919 5.3565 97.971 5.3565 97.971 5.207 50.637 5.207 50.637 4.607 78.672 4.607 78.672 5.207 97.971 5.207 97.971 4.9255 80.577 4.9255 80.577 4.4765 0.3 4.4765 0.3 3.8765 33.328 3.8765 33.328 4.4765 33.928 4.4765 33.928 3.8765 48.919 3.8765 48.919 4.4765 80.577 4.4765 80.577 4.4755 95.823 4.4755 95.823 4.9255 97.971 4.9255 97.971 4.307 50.637 4.307 50.637 3.707 63.1455 3.707 63.1455 4.307 63.6785 4.307 63.6785 3.707 78.672 3.707 78.672 4.307 97.971 4.307 97.971 3.9715 79.335 3.9715 79.335 3.5765 0.3 3.5765 0.3 2.9765 48.919 2.9765 48.919 3.5765 79.335 3.5765 79.335 3.4135 88.673 3.4135 88.673 3.9715 89.123 3.9715 89.123 3.4135 97.065 3.4135 97.065 3.9715 97.971 3.9715 97.971 3.407 50.637 3.407 50.637 2.807 78.672 2.807 78.672 3.407 97.971 3.407 97.971 2.9635 79.335 2.9635 79.335 2.7075 33.928 2.7075 33.928 2.6965 0.3 2.6965 0.3 2.0965 33.328 2.0965 33.328 2.6965 33.928 2.6965 33.928 2.1075 48.919 2.1075 48.919 2.7075 79.335 2.7075 79.335 2.507 50.637 2.507 50.637 1.907 63.1455 1.907 63.1455 2.507 63.6785 2.507 63.6785 1.907 78.672 1.907 78.672 2.507 79.335 2.507 79.335 2.4055 97.065 2.4055 97.065 2.9635 97.971 2.9635 97.971 1.7965 0.3 1.7965 0.3 1.1965 48.919 1.1965 48.919 1.7965 97.971 1.7965 97.971 0 ;
  END
END dwc_lpddr5xphy_txrxdq_ew

END LIBRARY
