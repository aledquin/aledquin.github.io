.options scale=1
*.LENGTH_UNIT lr wr rad gdis s pj S spacing ftip dw al aw
*.AREA_UNIT a 
*.NON_UNIT nr m lay passw ctapw ppitch
*.SCALE METER
*.LDD
.subckt dwc_lpddr5xphy_techrevision_sg_tiehigh_lp5x VBN VBP VDD VSS X
*.PININFO VBN:I VBP:I VDD:I VSS:I X:O
MlxDummyGroup_1[0] VDD VDD VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_1[1] VDD VDD VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_1[2] X VDD VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MMP3 X NL VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_0[0] VSS VSS VSS VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_0[1] VSS VSS VSS VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_0[2] VSS VSS NL VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MMN2 NL NL VSS VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
.ends dwc_lpddr5xphy_techrevision_sg_tiehigh_lp5x
.subckt dwc_lpddr5xphy_techrevision_sg_tielow_lp5x VBN VBP VDD VSS X
*.PININFO VBN:I VBP:I VDD:I VSS:I X:O
MlxDummyGroup_1[0] VSS VSS VSS VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_1[1] VSS VSS VSS VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_1[2] VSS VSS X VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MMN3 X NH VSS VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_0[0] VDD VDD VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_0[1] VDD VDD VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MlxDummyGroup_0[2] VDD VDD NH VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MMP2 NH NH VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
.ends dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
.subckt dwc_lpddr5xphy_techrevision_sg_endcell_right_lp5x VBN VBP VDD VSS
*.PININFO VBN:I VBP:I VDD:I VSS:I
MMNA VSS VSS VSS VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MMPA VDD VDD VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
.ends dwc_lpddr5xphy_techrevision_sg_endcell_right_lp5x
.subckt dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x VBN VBP VDD VSS
*.PININFO VBN:I VBP:I VDD:I VSS:I
MN1 VSS VSS VSS VBN nch_lvt_mac l=3n nfin=2 m=4 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MP0 VDD VDD VDD VBP pch_lvt_mac l=3n nfin=2 m=4 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
.ends dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
.subckt dwc_lpddr5xphy_techrevision_sg_endcell_left_lp5x VBN VBP VDD VSS
*.PININFO VBN:I VBP:I VDD:I VSS:I
MMNA VSS VSS VSS VBN nch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
MMPA VDD VDD VDD VBP pch_lvt_mac l=3n nfin=2 m=2 ppitch=0  mosdmy=0 fbound=1 fboundt=1 fboundb=1
.ends dwc_lpddr5xphy_techrevision_sg_endcell_left_lp5x
.subckt dwc_lpddr5xphy_techrevision VDD VSS tech_revision[15] tech_revision[14] tech_revision[13] tech_revision[12] tech_revision[11] tech_revision[10] tech_revision[9] tech_revision[8] tech_revision[7] tech_revision[6] tech_revision[5] tech_revision[4]
+ tech_revision[3] tech_revision[2] tech_revision[1] tech_revision[0]
*.PININFO VDD:I VSS:I tech_revision[15]:O tech_revision[14]:O tech_revision[13]:O tech_revision[12]:O tech_revision[11]:O tech_revision[10]:O tech_revision[9]:O tech_revision[8]:O tech_revision[7]:O tech_revision[6]:O tech_revision[5]:O tech_revision[4]:O
*.PININFO tech_revision[3]:O tech_revision[2]:O tech_revision[1]:O tech_revision[0]:O
XXREV5 VSS VDD VDD VSS tech_revision[5] dwc_lpddr5xphy_techrevision_sg_tiehigh_lp5x
XXREV7 VSS VDD VDD VSS tech_revision[7] dwc_lpddr5xphy_techrevision_sg_tiehigh_lp5x
XXREV11 VSS VDD VDD VSS tech_revision[11] dwc_lpddr5xphy_techrevision_sg_tiehigh_lp5x
XXREV14 VSS VDD VDD VSS tech_revision[14] dwc_lpddr5xphy_techrevision_sg_tiehigh_lp5x
XI0 VSS VDD VDD VSS tech_revision[0] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV1 VSS VDD VDD VSS tech_revision[1] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV2 VSS VDD VDD VSS tech_revision[2] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV3 VSS VDD VDD VSS tech_revision[3] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV4 VSS VDD VDD VSS tech_revision[4] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV6 VSS VDD VDD VSS tech_revision[6] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV8 VSS VDD VDD VSS tech_revision[8] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV9 VSS VDD VDD VSS tech_revision[9] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV10 VSS VDD VDD VSS tech_revision[10] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV12 VSS VDD VDD VSS tech_revision[12] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV13 VSS VDD VDD VSS tech_revision[13] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XXREV15 VSS VDD VDD VSS tech_revision[15] dwc_lpddr5xphy_techrevision_sg_tielow_lp5x
XI257[3] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_endcell_right_lp5x
XI257[2] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_endcell_right_lp5x
XI257[1] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_endcell_right_lp5x
XI257[0] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_endcell_right_lp5x
XXFILLER[0] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[1] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[2] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[3] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[4] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[5] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[6] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[7] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[8] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[9] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[10] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[11] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[12] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[13] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[14] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[15] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[16] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[17] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[18] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[19] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[20] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[21] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[22] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[23] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[24] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[25] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[26] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[27] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[28] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[29] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[30] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[31] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[32] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[33] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[34] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[35] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[36] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[37] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[38] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[39] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[40] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[41] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[42] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[43] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[44] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[45] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[46] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[47] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[48] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[49] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[50] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[51] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[52] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[53] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[54] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[55] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[56] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[57] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[58] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[59] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[60] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[61] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[62] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[63] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[64] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[65] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[66] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[67] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[68] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[69] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[70] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[71] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[72] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[73] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[74] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[75] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[76] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[77] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[78] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[79] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[80] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[81] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[82] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[83] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[84] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[85] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[86] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[87] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[88] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[89] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[90] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[91] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[92] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[93] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[94] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[95] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[96] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[97] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[98] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[99] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[100] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[101] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[102] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[103] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[104] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[105] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[106] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[107] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[108] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[109] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[110] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[111] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[112] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[113] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[114] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[115] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[116] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[117] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[118] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[119] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[120] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[121] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[122] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[123] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[124] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[125] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[126] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[127] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[128] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[129] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[130] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[131] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[132] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[133] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[134] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[135] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[136] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[137] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[138] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[139] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[140] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[141] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[142] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[143] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[144] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[145] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[146] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[147] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[148] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[149] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[150] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[151] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[152] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[153] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[154] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[155] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[156] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[157] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[158] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[159] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[160] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[161] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[162] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[163] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[164] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[165] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[166] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[167] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[168] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[169] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[170] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[171] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[172] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[173] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[174] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[175] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[176] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[177] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[178] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[179] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[180] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[181] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[182] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[183] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[184] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[185] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[186] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[187] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[188] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[189] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[190] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[191] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[192] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[193] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[194] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[195] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[196] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[197] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[198] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[199] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[200] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[201] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[202] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[203] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[204] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[205] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[206] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XXFILLER[207] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_fillerx2r_lp5x
XI258[3] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_endcell_left_lp5x
XI258[2] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_endcell_left_lp5x
XI258[1] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_endcell_left_lp5x
XI258[0] VSS VDD VDD VSS dwc_lpddr5xphy_techrevision_sg_endcell_left_lp5x
.ends dwc_lpddr5xphy_techrevision
