# LEF OUT API 
# Creation Date : Wed Jun 22 09:27:00 IST 2022
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_lpddr5xphy_zcalio_ew
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_lpddr5xphy_zcalio_ew 0 0 ;
  SYMMETRY X Y ;
  SIZE 194.055 BY 74.76 ;
  PIN csrTxDcaFinePU0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 137.038 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.717 0.038 2.755 ;
    END
  END csrTxDcaFinePU0[2]
  PIN csrTxDcaFinePU0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 113.297 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.413 0.033 2.451 ;
    END
  END csrTxDcaFinePU0[1]
  PIN csrTxDcaFinePD0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 126.295 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.653 0.034 1.691 ;
    END
  END csrTxDcaFinePD0[1]
  PIN csrLsTxCalCodePD1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 489.454 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.731 37.43 145.769 74.71 ;
    END
  END csrLsTxCalCodePD1[1]
  PIN csrLsTxCalCodePD1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 481.928 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.807 37.43 145.845 74.71 ;
    END
  END csrLsTxCalCodePD1[2]
  PIN csrLsTxCalCodePD1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 473.961 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.883 37.43 145.921 74.71 ;
    END
  END csrLsTxCalCodePD1[3]
  PIN csrLsTxCalCodePD1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 467.395 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.959 37.43 145.997 74.71 ;
    END
  END csrLsTxCalCodePD1[4]
  PIN csrLsTxCalCodePD1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 460.751 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.035 37.43 146.073 74.71 ;
    END
  END csrLsTxCalCodePD1[5]
  PIN csrLsTxCalCodePD1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 429.749 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.111 37.43 146.149 74.71 ;
    END
  END csrLsTxCalCodePD1[6]
  PIN csrLsTxCalCodePD0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 473.961 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.883 0.05 145.921 37.33 ;
    END
  END csrLsTxCalCodePD0[3]
  PIN csrLsTxCalCodePD1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 440.839 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.263 37.43 146.301 74.71 ;
    END
  END csrLsTxCalCodePD1[8]
  PIN csrLsTxCalCodeLPPU0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 482.52 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.339 0.05 146.377 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[0]
  PIN csrLsTxCalCodeLPPU0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 466.08 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.491 0.05 146.529 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[2]
  PIN csrLsTxCalCodeLPPU0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 378.076 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.947 0.05 146.985 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[8]
  PIN csrLsTxCalCodeLPPU0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 399.026 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.795 0.05 146.833 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[6]
  PIN csrLsTxCalCodeLPPU0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 428.826 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.719 0.05 146.757 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[5]
  PIN csrLsTxCalCodeLPPU0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 429.877 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.643 0.05 146.681 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[4]
  PIN csrLsTxCalCodeLPPU0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 453.838 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.567 0.05 146.605 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[3]
  PIN csrLsTxCalCodeLPPU0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 462.54 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.415 0.05 146.453 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[1]
  PIN csrLsTxCalCodeLPPU1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 482.52 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.339 37.43 146.377 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[0]
  PIN csrLsTxCalCodeLPPU1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 462.54 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.415 37.43 146.453 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[1]
  PIN csrLsTxSlewLPPU0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 321.322 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 144.971 0.05 145.009 37.33 ;
    END
  END csrLsTxSlewLPPU0[0]
  PIN csrLsTxSlewLPPU0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 319.472 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.047 0.05 145.085 37.33 ;
    END
  END csrLsTxSlewLPPU0[1]
  PIN csrLsTxSlewLPPU0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 347.754 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 144.895 0.05 144.933 37.33 ;
    END
  END csrLsTxSlewLPPU0[2]
  PIN csrLsTxSlewPD0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 314.013 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.123 0.05 145.161 37.33 ;
    END
  END csrLsTxSlewPD0[0]
  PIN csrLsTxSlewPD0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 308.815 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.199 0.05 145.237 37.33 ;
    END
  END csrLsTxSlewPD0[1]
  PIN VIO_TXBE0_PAD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8607 LAYER M10 ;
    ANTENNADIFFAREA 3.9769 LAYER M10 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 6.5367 LAYER M10 ;
      ANTENNAMAXAREACAR 6.51602 LAYER M10 ;
    PORT
      LAYER M10 ;
        RECT 160.4665 30.9755 172.52 31.4255 ;
        RECT 160.4665 19.5515 172.52 20.0015 ;
        RECT 160.4665 8.1275 172.52 8.5775 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 6.4915 191.907 6.9415 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 4.4755 191.907 4.9255 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 8.5075 191.907 8.9575 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 18.5875 191.907 19.0375 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 10.5235 191.907 10.9735 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 12.5395 191.907 12.9895 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 16.5715 191.907 17.0215 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 22.6195 191.907 23.0695 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 24.6355 191.907 25.0855 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 20.6035 191.907 21.0535 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 14.5555 191.907 15.0055 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 26.6515 191.907 27.1015 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 30.6835 191.907 31.1335 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 32.6995 191.907 33.1495 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 28.6675 191.907 29.1175 ;
    END
  END VIO_TXBE0_PAD
  PIN TIEHI0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.46024 LAYER M6 ;
    ANTENNADIFFAREA 0.00459 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.354 0.038 0.392 ;
    END
  END TIEHI0
  PIN VIO_TXBE1_PAD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8607 LAYER M10 ;
    ANTENNADIFFAREA 3.9769 LAYER M10 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 6.5367 LAYER M10 ;
      ANTENNAMAXAREACAR 6.51602 LAYER M10 ;
    PORT
      LAYER M10 ;
        RECT 160.4665 45.5075 172.52 45.9575 ;
    END
    PORT
      LAYER M10 ;
        RECT 160.4665 56.9315 172.52 57.3815 ;
    END
    PORT
      LAYER M10 ;
        RECT 160.4665 68.3555 172.52 68.8055 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 43.8715 191.907 44.3215 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 41.8555 191.907 42.3055 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 45.8875 191.907 46.3375 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 55.9675 191.907 56.4175 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 47.9035 191.907 48.3535 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 49.9195 191.907 50.3695 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 53.9515 191.907 54.4015 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 59.9995 191.907 60.4495 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 62.0155 191.907 62.4655 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 57.9835 191.907 58.4335 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 51.9355 191.907 52.3855 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 64.0315 191.907 64.4815 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 68.0635 191.907 68.5135 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 70.0795 191.907 70.5295 ;
    END
    PORT
      LAYER M10 ;
        RECT 176.661 66.0475 191.907 66.4975 ;
    END
  END VIO_TXBE1_PAD
  PIN csrLsTxSlewPD0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 305.882 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.275 0.05 145.313 37.33 ;
    END
  END csrLsTxSlewPD0[2]
  PIN csrLsTxCalCodeLPPU1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 466.08 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.491 37.43 146.529 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[2]
  PIN TIELO0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.45342 LAYER M6 ;
    ANTENNADIFFAREA 0.00918 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 0.278 0.038 0.316 ;
    END
  END TIELO0
  PIN csrLsTxSlewPD0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 331.005 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.351 0.05 145.389 37.33 ;
    END
  END csrLsTxSlewPD0[3]
  PIN csrLsTxSlewPD1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 331.005 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.351 37.43 145.389 74.71 ;
    END
  END csrLsTxSlewPD1[3]
  PIN csrTxSeg120PU1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 91.5509 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 41.629 0.038 41.667 ;
    END
  END csrTxSeg120PU1[2]
  PIN csrOdtSeg120PU1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 96.6108 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 41.173 0.038 41.211 ;
    END
  END csrOdtSeg120PU1[2]
  PIN csrOdtSeg120PD1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.1059 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 43.301 0.038 43.339 ;
    END
  END csrOdtSeg120PD1[2]
  PIN csrTxSeg120PD1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024529 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.1897 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 43.453 0.038 43.491 ;
    END
  END csrTxSeg120PD1[2]
  PIN csrTxDcaFinePD0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 75.8058 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.957 0.034 1.995 ;
    END
  END csrTxDcaFinePD0[0]
  PIN scan_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.080959 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.09384 LAYER M6 ;
      ANTENNAMAXAREACAR 90.30759975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 48.925 0.038 48.963 ;
    END
  END scan_mode
  PIN csrTxDcaMode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.02964 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0.465234 LAYER M7 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00816 LAYER M7 ;
      ANTENNAMAXAREACAR 384.2 LAYER M7 ;
    PORT
      LAYER M6 ;
        RECT 0 37.373 0.038 37.411 ;
    END
  END csrTxDcaMode
  PIN csrTxDcaFinePU1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 85.19929975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 40.261 0.033 40.299 ;
    END
  END csrTxDcaFinePU1[3]
  PIN csrTxSeg120PD1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.8632 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 69.825 0.038 69.863 ;
    END
  END csrTxSeg120PD1[1]
  PIN csrTxSeg120PD1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 92.5245 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 72.713 0.038 72.751 ;
    END
  END csrTxSeg120PD1[0]
  PIN csrTxSeg120PU1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.8774 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 71.117 0.038 71.155 ;
    END
  END csrTxSeg120PU1[0]
  PIN csrOdtSeg120PD1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 97.7667 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 70.129 0.038 70.167 ;
    END
  END csrOdtSeg120PD1[1]
  PIN csrOdtSeg120PD1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 100.681 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 73.093 0.038 73.131 ;
    END
  END csrOdtSeg120PD1[0]
  PIN csrTxSeg120PU1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 85.5019 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 68.229 0.038 68.267 ;
    END
  END csrTxSeg120PU1[1]
  PIN csrOdtSeg120PU1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 101.721 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 71.497 0.038 71.535 ;
    END
  END csrOdtSeg120PU1[0]
  PIN csrCoreLoopBackMode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.084721 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00816 LAYER M6 ;
      ANTENNAMAXAREACAR 138.722 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 15.941 0.038 15.979 ;
    END
  END csrCoreLoopBackMode
  PIN TxFwdClk1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.029564 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 56.145 0.038 56.183 ;
    END
  END TxFwdClk1
  PIN TxClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028633 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 1.42671 LAYER M7 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03066 LAYER M7 ;
      ANTENNAMAXAREACAR 58.1773 LAYER M7 ;
    PORT
      LAYER M6 ;
        RECT 0 37.601 0.038 37.639 ;
    END
  END TxClk
  PIN TxDataEven1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034808 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 65.25889975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 57.513 0.038 57.551 ;
    END
  END TxDataEven1
  PIN TxOEOdd1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026619 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00867 LAYER M6 ;
      ANTENNAMAXAREACAR 34.4283 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 54.321 0.038 54.359 ;
    END
  END TxOEOdd1
  PIN TxOEEven1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034789 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00867 LAYER M6 ;
      ANTENNAMAXAREACAR 34.0927 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 54.017 0.038 54.055 ;
    END
  END TxOEEven1
  PIN OdtEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.04339 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 0.00758 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 0.16908 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 0.028025 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 1.42263975 LAYER M7 ;
    ANTENNAPARTIALCUTAREA 0.000256 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.001 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M2 ;
      ANTENNAGATEAREA 0.00305975 LAYER M3 ;
      ANTENNAGATEAREA 0.00305975 LAYER M4 ;
      ANTENNAGATEAREA 0.00611975 LAYER M7 ;
      ANTENNAGATEAREA 0.00305975 LAYER VIA2 ;
      ANTENNAGATEAREA 0.00305975 LAYER VIA3 ;
      ANTENNAGATEAREA 0.00305975 LAYER VIA4 ;
      ANTENNAMAXAREACAR 31.9385 LAYER M2 ;
      ANTENNAMAXAREACAR 34.4156 LAYER M3 ;
      ANTENNAMAXAREACAR 89.6705 LAYER M4 ;
      ANTENNAMAXAREACAR 337.886 LAYER M7 ;
      ANTENNAMAXCUTCAR 0.52679675 LAYER VIA2 ;
      ANTENNAMAXCUTCAR 0.85359375 LAYER VIA3 ;
      ANTENNAMAXCUTCAR 1.32549 LAYER VIA4 ;
    PORT
      LAYER M6 ;
        RECT 0 37.525 0.038 37.563 ;
    END
  END OdtEn
  PIN csrLsTxCalCodePD0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 500.006 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.655 0.05 145.693 37.33 ;
    END
  END csrLsTxCalCodePD0[0]
  PIN csrTxDcaFinePU1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 137.038 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 39.957 0.038 39.995 ;
    END
  END csrTxDcaFinePU1[2]
  PIN csrTxDcaFinePU1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 113.297 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 39.653 0.033 39.691 ;
    END
  END csrTxDcaFinePU1[1]
  PIN csrTxDcaFinePD1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 126.295 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.893 0.034 38.931 ;
    END
  END csrTxDcaFinePD1[1]
  PIN csrTxDcaFinePD1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 75.8058 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 39.197 0.034 39.235 ;
    END
  END csrTxDcaFinePD1[0]
  PIN csrTxDcaFinePD1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 82.3451 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.437 0.034 38.475 ;
    END
  END csrTxDcaFinePD1[3]
  PIN csrTxDcaFinePU1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 85.9592 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 39.501 0.033 39.539 ;
    END
  END csrTxDcaFinePU1[0]
  PIN csrTxDcaFinePD1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 179.17 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.741 0.034 38.779 ;
    END
  END csrTxDcaFinePD1[2]
  PIN csrTxDcaCoarse1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 116.091 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 40.413 0.033 40.451 ;
    END
  END csrTxDcaCoarse1[1]
  PIN csrLsTxCalCodePD1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 500.006 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.655 37.43 145.693 74.71 ;
    END
  END csrLsTxCalCodePD1[0]
  PIN csrTxDcaCoarse1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 125.773 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 40.717 0.033 40.755 ;
    END
  END csrTxDcaCoarse1[0]
  PIN csrTxDcaFinePD0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 82.3451 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.197 0.034 1.235 ;
    END
  END csrTxDcaFinePD0[3]
  PIN csrTxDcaFinePU0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 85.9592 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 2.261 0.033 2.299 ;
    END
  END csrTxDcaFinePU0[0]
  PIN csrTxDcaFinePD0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 179.17 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 1.501 0.034 1.539 ;
    END
  END csrTxDcaFinePD0[2]
  PIN csrTxDcaCoarse0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 116.091 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.173 0.033 3.211 ;
    END
  END csrTxDcaCoarse0[1]
  PIN TxDataOdd1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026182 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 82.7265 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 57.969 0.038 58.007 ;
    END
  END TxDataOdd1
  PIN csrLsTxCalCodePD0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 467.395 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.959 0.05 145.997 37.33 ;
    END
  END csrLsTxCalCodePD0[4]
  PIN TxBypassModeInt1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026619 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 195.885 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 55.309 0.038 55.347 ;
    END
  END TxBypassModeInt1
  PIN TxBypassDataInt1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.025156 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 324.389 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 56.981 0.038 57.019 ;
    END
  END TxBypassDataInt1
  PIN TxBypassModeExt1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034998 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 134.881 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 56.221 0.038 56.259 ;
    END
  END TxBypassModeExt1
  PIN TxBypassOEExt1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022781 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 377.175 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 57.209 0.038 57.247 ;
    END
  END TxBypassOEExt1
  PIN TxBypassOEInt1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.027949 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 364.115 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 55.537 0.038 55.575 ;
    END
  END TxBypassOEInt1
  PIN csrTxDcaCoarse0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 125.773 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.477 0.033 3.515 ;
    END
  END csrTxDcaCoarse0[0]
  PIN csrLsTxCalCodePD0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 460.751 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.035 0.05 146.073 37.33 ;
    END
  END csrLsTxCalCodePD0[5]
  PIN TxOEEven0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034789 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00867 LAYER M6 ;
      ANTENNAMAXAREACAR 34.0927 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 16.777 0.038 16.815 ;
    END
  END TxOEEven0
  PIN csrLsTxCalCodePD0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 429.749 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.111 0.05 146.149 37.33 ;
    END
  END csrLsTxCalCodePD0[6]
  PIN csrLsTxCalCodePD0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 440.839 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.263 0.05 146.301 37.33 ;
    END
  END csrLsTxCalCodePD0[8]
  PIN csrLsTxCalCodePD0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 448.87 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.187 0.05 146.225 37.33 ;
    END
  END csrLsTxCalCodePD0[7]
  PIN csrLsTxCalCodePD0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 489.454 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.731 0.05 145.769 37.33 ;
    END
  END csrLsTxCalCodePD0[1]
  PIN csrOdtSeg120PU1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 98.2799 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 68.457 0.038 68.495 ;
    END
  END csrOdtSeg120PU1[1]
  PIN csrTxSeg120PU0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 91.5509 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 4.389 0.038 4.427 ;
    END
  END csrTxSeg120PU0[2]
  PIN csrOdtSeg120PU0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 96.6108 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.933 0.038 3.971 ;
    END
  END csrOdtSeg120PU0[2]
  PIN csrOdtSeg120PD0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.1059 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 6.061 0.038 6.099 ;
    END
  END csrOdtSeg120PD0[2]
  PIN TxBypassDataExt1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024282 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 327.172 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 56.601 0.038 56.639 ;
    END
  END TxBypassDataExt1
  PIN csrTxSeg120PD0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024529 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.1897 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 6.213 0.038 6.251 ;
    END
  END csrTxSeg120PD0[2]
  PIN csrOdtSeg120PU0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 98.2799 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 31.217 0.038 31.255 ;
    END
  END csrOdtSeg120PU0[1]
  PIN csrTxSeg120PD0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022933 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.8632 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 32.585 0.038 32.623 ;
    END
  END csrTxSeg120PD0[1]
  PIN csrTxSeg120PD0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 92.5245 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.473 0.038 35.511 ;
    END
  END csrTxSeg120PD0[0]
  PIN csrTxSeg120PU0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 87.8774 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.877 0.038 33.915 ;
    END
  END csrTxSeg120PU0[0]
  PIN csrOdtSeg120PD0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 97.7667 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 32.889 0.038 32.927 ;
    END
  END csrOdtSeg120PD0[1]
  PIN csrOdtSeg120PD0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 100.681 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.853 0.038 35.891 ;
    END
  END csrOdtSeg120PD0[0]
  PIN csrTxSeg120PU0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023636 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 85.5019 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 30.989 0.038 31.027 ;
    END
  END csrTxSeg120PU0[1]
  PIN TxDataOdd0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026182 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 82.7265 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 20.729 0.038 20.767 ;
    END
  END TxDataOdd0
  PIN csrLsTxCalCodePD0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 481.928 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.807 0.05 145.845 37.33 ;
    END
  END csrLsTxCalCodePD0[2]
  PIN TxBypassOEExt0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.022781 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 377.175 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 19.969 0.038 20.007 ;
    END
  END TxBypassOEExt0
  PIN TxBypassOEInt0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.027949 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 364.115 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.297 0.038 18.335 ;
    END
  END TxBypassOEInt0
  PIN TxBypassModeInt0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026619 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 195.885 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.069 0.038 18.107 ;
    END
  END TxBypassModeInt0
  PIN TxBypassDataInt0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.025156 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 324.389 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 19.741 0.038 19.779 ;
    END
  END TxBypassDataInt0
  PIN TxBypassModeExt0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034998 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 134.881 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.981 0.038 19.019 ;
    END
  END TxBypassModeExt0
  PIN TxBypassDataExt0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024282 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 327.172 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 19.361 0.038 19.399 ;
    END
  END TxBypassDataExt0
  PIN csrLsTxCalCodePD1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 448.87 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.187 37.43 146.225 74.71 ;
    END
  END csrLsTxCalCodePD1[7]
  PIN csrOdtSeg120PU0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.024662 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 101.721 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 34.257 0.038 34.295 ;
    END
  END csrOdtSeg120PU0[0]
  PIN TxFwdClk0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.029564 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 18.905 0.038 18.943 ;
    END
  END TxFwdClk0
  PIN TxDataEven0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.034808 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 65.25889975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 20.273 0.038 20.311 ;
    END
  END TxDataEven0
  PIN TxOEOdd0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.026619 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00867 LAYER M6 ;
      ANTENNAMAXAREACAR 34.4283 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 17.081 0.038 17.119 ;
    END
  END TxOEOdd0
  PIN csrTxDcaFinePU0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.028823 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 85.19929975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 3.021 0.033 3.059 ;
    END
  END csrTxDcaFinePU0[3]
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M10 ;
        RECT 159.7625 63.935 174.756 64.535 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 62.135 174.756 62.735 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 10.4465 174.756 11.0465 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 70.6745 174.756 71.2745 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 52.511 174.756 53.111 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.608 60.3195 122.5515 60.9195 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 23.6705 174.756 24.2705 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 41.087 174.756 41.687 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 42.887 174.7565 43.487 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 72.4745 174.756 73.0745 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6575 41.1165 122.5515 41.7165 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 47.8265 174.756 48.4265 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 24.755 174.756 25.355 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 1.907 174.756 2.507 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 21.8705 174.756 22.4705 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 5.507 174.7565 6.107 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 13.331 174.756 13.931 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 15.131 174.756 15.731 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 3.707 174.756 4.307 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 26.555 174.756 27.155 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 49.6265 174.756 50.2265 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 16.931 174.7565 17.531 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 61.0505 174.756 61.6505 ;
    END
    PORT
      LAYER M10 ;
        RECT 144.198 65.735 174.756 66.335 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 28.355 174.756 28.955 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 59.2505 174.756 59.8505 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.5945 54.311 174.7565 54.911 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 33.2945 174.756 33.8945 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6575 34.7185 122.5515 35.3185 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 50.711 174.756 51.311 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 39.287 174.756 39.887 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 12.2465 174.756 12.8465 ;
    END
    PORT
      LAYER M10 ;
        RECT 159.7625 35.0945 174.756 35.6945 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 70.0195 144.6645 70.6195 ;
    END
    PORT
      LAYER M10 ;
        RECT 106.5155 37.4775 122.5515 38.0775 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 42.8095 193.149 43.3675 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 46.8415 193.149 47.3995 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 40.7935 193.149 41.3515 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 44.8255 193.149 45.3835 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 48.8575 193.149 49.4155 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 58.9375 193.149 59.4955 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 50.8735 193.149 51.4315 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 54.9055 193.149 55.4635 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 52.8895 193.149 53.4475 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 60.9535 193.149 61.5115 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 56.9215 193.149 57.4795 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 72.0415 193.149 72.5995 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 62.9695 193.149 63.5275 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 71.0335 193.149 71.5915 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 67.0015 193.149 67.5595 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 64.9855 193.149 65.5435 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 69.0175 193.149 69.5755 ;
    END
    PORT
      LAYER M10 ;
        RECT 106.5155 44.6765 122.5515 45.2765 ;
    END
    PORT
      LAYER M10 ;
        RECT 106.5155 49.4565 122.5515 50.0565 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6155 48.5565 122.5515 49.1565 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6125 21.5375 122.5515 22.0375 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 5.4295 193.149 5.9875 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 9.4615 193.149 10.0195 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 3.4135 193.149 3.9715 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 7.4455 193.149 8.0035 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 11.4775 193.149 12.0355 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 21.5575 193.149 22.1155 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 13.4935 193.149 14.0515 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 17.5255 193.149 18.0835 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 15.5095 193.149 16.0675 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 23.5735 193.149 24.1315 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 19.5415 193.149 20.0995 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 34.6615 193.149 35.2195 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 25.5895 193.149 26.1475 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 33.6535 193.149 34.2115 ;
    END
    PORT
      LAYER M10 ;
        RECT 183.811 29.6215 193.149 30.1795 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 27.6055 193.149 28.1635 ;
    END
    PORT
      LAYER M10 ;
        RECT 185.207 31.6375 193.149 32.1955 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 67.9195 104.4075 68.5195 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 66.1195 104.4075 66.7195 ;
    END
    PORT
      LAYER M10 ;
        RECT 30.1505 71.9585 104.4075 72.5585 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 64.3195 104.4075 64.9195 ;
    END
    PORT
      LAYER M10 ;
        RECT 106.5155 51.5565 122.5515 52.1565 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.608 58.3505 122.5515 58.9505 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6575 30.6795 122.5515 31.2795 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 62.5195 144.5875 63.1195 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6575 27.0795 122.5515 27.6795 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M10 ;
        RECT 0.3 41.1165 6.225 41.7165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 52.4565 6.225 53.0565 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 58.5195 23.561 59.1195 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 34.7185 14.994 35.3185 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 28.8795 14.331 29.4795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 39.3365 6.225 39.9365 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 53.439 6.225 54.039 ;
    END
    PORT
      LAYER M10 ;
        RECT 16.3205 21.4575 36.1665 21.9575 ;
    END
    PORT
      LAYER M10 ;
        RECT 12.643 18.2795 29.657 18.8795 ;
    END
    PORT
      LAYER M10 ;
        RECT 12.643 16.4795 25.6785 17.0795 ;
    END
    PORT
      LAYER M10 ;
        RECT 6.4745 15.5795 17.2005 16.1795 ;
    END
    PORT
      LAYER M10 ;
        RECT 6.475 17.3795 12.393 17.9795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 23.0795 6.225 23.6795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 16.199 6.225 16.799 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 17.999 6.225 18.599 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 14.3165 6.225 14.9165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 55.239 6.225 55.839 ;
    END
    PORT
      LAYER M10 ;
        RECT 37.835 34.7215 104.4075 35.3215 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 0.1465 146.1975 0.5965 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 12.2165 25.6785 12.8165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 21.2795 14.8105 21.8795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 2.0965 6.225 2.6965 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 3.8765 6.225 4.4765 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 7.4365 146.1975 8.0365 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 15.2165 6.225 15.8165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 32.7795 122.5515 33.3795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 30.6795 104.4075 31.2795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 62.5195 36.164 63.1195 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 44.6765 106.3105 45.2765 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 67.9195 25.5555 68.5195 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 42.8965 122.5515 43.4965 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 64.3195 36.164 64.9195 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 46.7765 122.5515 47.3765 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 39.3365 122.5515 39.9365 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 41.1165 104.4075 41.7165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 60.3195 23.561 60.9195 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 49.4565 36.164 50.0565 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 51.5565 6.225 52.1565 ;
    END
    PORT
      LAYER M10 ;
        RECT 6.475 13.2095 146.1975 13.7895 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 66.1195 25.5555 66.7195 ;
    END
    PORT
      LAYER M10 ;
        RECT 120.928 17.7315 146.1975 18.1815 ;
    END
    PORT
      LAYER M10 ;
        RECT 125.927 11.3165 146.1975 11.9165 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6125 22.7375 122.5515 23.3375 ;
    END
    PORT
      LAYER M10 ;
        RECT 124.627 21.5375 141.574 22.1375 ;
    END
    PORT
      LAYER M10 ;
        RECT 146.721 62.135 159.2295 62.735 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 5.6565 146.1975 6.2565 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 15.8095 146.198 16.3895 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 21.4575 104.4075 22.0375 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 13.331 159.2295 13.931 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 58.3705 104.4075 58.9505 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 56.4195 36.164 57.0195 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 35.0945 159.2295 35.6945 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 3.707 159.2295 4.307 ;
        RECT 36.414 2.0965 146.1975 2.6965 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 24.0575 104.4075 24.6375 ;
    END
    PORT
      LAYER M10 ;
        RECT 29.1195 22.7375 36.1665 23.3375 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 41.087 159.2295 41.687 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 9.5365 146.1975 10.1365 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 3.8765 146.1975 4.4765 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 70.0195 36.164 70.6195 ;
    END
    PORT
      LAYER M10 ;
        RECT 146.721 70.6745 159.2295 71.2745 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 21.8705 159.2295 22.4705 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 39.287 159.2295 39.887 ;
    END
    PORT
      LAYER M10 ;
        RECT 146.721 72.4745 159.2295 73.0745 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 50.711 159.2295 51.311 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 26.555 159.2295 27.155 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 47.8265 159.2295 48.4265 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 10.4465 159.2295 11.0465 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 33.2945 159.2295 33.8945 ;
    END
    PORT
      LAYER M10 ;
        RECT 146.721 63.935 159.2295 64.535 ;
    END
    PORT
      LAYER M10 ;
        RECT 146.721 61.0505 159.2295 61.6505 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 60.9705 104.4075 61.5505 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 49.6265 159.2295 50.2265 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 52.511 159.2295 53.111 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 12.2465 159.2295 12.8465 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 19.1795 104.4075 19.7795 ;
    END
    PORT
      LAYER M10 ;
        RECT 6.427 52.7225 106.3105 53.3025 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 50.1225 106.3105 50.7025 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 1.907 159.2295 2.507 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 15.131 159.2295 15.731 ;
    END
    PORT
      LAYER M10 ;
        RECT 146.721 59.2505 159.2295 59.8505 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 23.6705 159.2295 24.2705 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 42.8965 6.225 43.4965 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 46.7765 6.225 47.3765 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 27.0795 104.4075 27.6795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 71.9585 25.5555 72.5585 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6565 28.8795 122.5515 29.4795 ;
    END
    PORT
      LAYER M10 ;
        RECT 142.55 24.755 159.2295 25.355 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 25.2795 104.4075 25.8795 ;
    END
  END VDD
  PIN PwrOkVDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.22458 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 3.94872 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0038 LAYER VIA7 ;
    ANTENNADIFFAREA 0.081528 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER M7 ;
      ANTENNAGATEAREA 0.09294 LAYER M8 ;
      ANTENNAGATEAREA 0.0162 LAYER VIA7 ;
      ANTENNAMAXAREACAR 459.694 LAYER M7 ;
      ANTENNAMAXAREACAR 502.181 LAYER M8 ;
      ANTENNAMAXCUTCAR 1.19062 LAYER VIA7 ;
    PORT
      LAYER M7 ;
        RECT 144.591 0.05 144.629 37.33 ;
    END
  END PwrOkVDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M10 ;
        RECT 0.3 59.4195 23.561 60.0195 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 43.7765 6.225 44.3765 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 38.4365 6.225 39.0365 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 35.6185 14.994 36.2185 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 41.9965 6.225 42.5965 ;
    END
    PORT
      LAYER M10 ;
        RECT 106.5155 52.4565 122.5515 53.0565 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.608 59.4195 122.5515 60.0195 ;
    END
    PORT
      LAYER M10 ;
        RECT 12.643 17.3795 25.6785 17.9795 ;
    END
    PORT
      LAYER M10 ;
        RECT 106.5155 36.5775 122.5515 37.1775 ;
    END
    PORT
      LAYER M10 ;
        RECT 17.47 15.5795 25.6785 16.1795 ;
    END
    PORT
      LAYER M10 ;
        RECT 146.721 63.035 174.756 63.635 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 48.7265 174.756 49.3265 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 41.987 174.756 42.587 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 34.1945 174.756 34.7945 ;
    END
    PORT
      LAYER M10 ;
        RECT 6.475 16.4795 12.393 17.0795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 61.2195 34.1535 61.8195 ;
    END
    PORT
      LAYER M10 ;
        RECT 6.475 18.2795 12.393 18.8795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 22.1795 6.225 22.7795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 17.099 6.225 17.699 ;
    END
    PORT
      LAYER M10 ;
        RECT 144.198 64.835 174.756 65.435 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 16.031 174.756 16.631 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 14.231 174.756 14.831 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 22.7705 174.756 23.3705 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 40.187 174.756 40.787 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 20.3795 146.198 20.9795 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 43.787 174.756 44.387 ;
        RECT 125.8405 10.4165 146.1975 11.0165 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 29.255 174.756 29.855 ;
    END
    PORT
      LAYER M10 ;
        RECT 144.198 71.5745 174.756 72.1745 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 6.5365 146.1975 7.1365 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 8.6365 146.1975 9.2365 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 51.611 174.756 52.211 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 23.9795 36.1665 24.5795 ;
    END
    PORT
      LAYER M10 ;
        RECT 146.721 60.1505 174.756 60.7505 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 2.9765 6.225 3.5765 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 2.807 174.756 3.407 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 4.7565 6.225 5.3565 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 55.211 174.756 55.811 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 10.4165 6.225 11.0165 ;
    END
    PORT
      LAYER M10 ;
        RECT 144.198 66.635 174.756 67.235 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 31.5795 122.5515 32.1795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 45.8765 122.5515 46.4765 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 33.8185 122.5515 34.4185 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 41.9965 122.5515 42.5965 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 43.7765 122.5515 44.3765 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 40.2165 122.5515 40.8165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 50.6565 6.225 51.2565 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 38.4365 122.5515 39.0365 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 53.411 174.756 54.011 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 48.829 104.4075 49.279 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 33.8185 25.842 34.4185 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 39.7855 193.149 40.3435 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 40.7935 184.757 41.3515 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 44.8255 184.757 45.3835 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 48.8575 184.757 49.4155 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 42.8095 183.361 43.3675 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 46.8415 183.361 47.3995 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 56.9215 184.757 57.4795 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 60.9535 184.757 61.5115 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 52.8895 184.757 53.4475 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 50.8735 183.361 51.4315 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 54.9055 183.361 55.4635 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 58.9375 183.361 59.4955 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 64.9855 184.757 65.5435 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 69.0175 184.757 69.5755 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 71.0335 183.361 71.5915 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 67.0015 183.361 67.5595 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 62.9695 183.361 63.5275 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 57.058 104.4075 57.638 ;
    END
    PORT
      LAYER M10 ;
        RECT 120.928 17.046 146.1975 17.496 ;
    END
    PORT
      LAYER M10 ;
        RECT 142.42 25.655 174.756 26.255 ;
    END
    PORT
      LAYER M10 ;
        RECT 122.232 12.2165 146.1975 12.8165 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 17.831 174.756 18.431 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 63.4195 104.4075 64.0195 ;
    END
    PORT
      LAYER M10 ;
        RECT 106.574 50.6565 122.5515 51.2565 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.6125 24.0375 122.5515 24.6375 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 4.607 174.756 5.207 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 6.407 174.756 7.007 ;
    END
    PORT
      LAYER M10 ;
        RECT 147.594 11.3465 174.756 11.9465 ;
    END
    PORT
      LAYER M10 ;
        RECT 141.8235 27.455 174.756 28.055 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 2.9765 146.1975 3.5765 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 5.0065 146.1975 5.4565 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 18.3795 104.4075 18.9795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 67.0195 25.5555 67.6195 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 22.7575 104.4075 23.3375 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 2.4055 193.149 2.9635 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 3.4135 184.757 3.9715 ;
    END
    PORT
      LAYER M10 ;
        RECT 6.475 14.5095 146.1975 15.0895 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 11.3165 6.225 11.9165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 1.1965 146.1975 1.7965 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 13.4165 6.225 14.0165 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 7.4455 184.757 8.0035 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 11.4775 184.757 12.0355 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 5.4295 183.361 5.9875 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 9.4615 183.361 10.0195 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 19.5415 184.757 20.0995 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 23.5735 184.757 24.1315 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 15.5095 184.757 16.0675 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 13.4935 183.361 14.0515 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 17.5255 183.361 18.0835 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 21.5575 183.361 22.1155 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 27.6055 184.757 28.1635 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 31.6375 184.757 32.1955 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 33.6535 183.361 34.2115 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 29.6215 183.361 30.1795 ;
    END
    PORT
      LAYER M10 ;
        RECT 175.419 25.5895 183.361 26.1475 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 57.6195 34.1535 58.2195 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.608 61.3575 144.5875 61.9575 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 54.339 104.4075 54.939 ;
    END
    PORT
      LAYER M10 ;
        RECT 6.427 51.4225 106.3105 52.0025 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 67.0195 104.4075 67.6195 ;
    END
    PORT
      LAYER M10 ;
        RECT 30.1505 71.0585 104.4075 71.6585 ;
    END
    PORT
      LAYER M10 ;
        RECT 36.414 59.6705 104.4075 60.2505 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 68.8195 144.6645 69.4195 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 72.8585 144.6645 73.4585 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 65.2195 143.9645 65.8195 ;
    END
    PORT
      LAYER M10 ;
        RECT 104.407 47.6565 122.5515 48.2565 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 40.2165 6.225 40.8165 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 47.6565 6.225 48.2565 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 48.5565 6.225 49.1565 ;
    END
    PORT
      LAYER M10 ;
        RECT 105.842 35.6185 122.5515 36.2185 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 29.7795 122.5515 30.3795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 71.0585 25.5555 71.6585 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 27.9795 122.5515 28.5795 ;
    END
    PORT
      LAYER M10 ;
        RECT 0.3 26.1795 122.5515 26.7795 ;
    END
  END VSS
  PIN VIO_PwrOk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.43948 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.31535975 LAYER M8 ;
      ANTENNAMAXAREACAR 24.9057 LAYER M8 ;
    PORT
      LAYER M8 ;
        RECT 36.414 37.992 36.494 38.072 ;
    END
  END VIO_PwrOk
  PIN LsScan_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3379 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 125.263 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 28.48 36.657 28.52 ;
    END
  END LsScan_mode
  PIN csrLsZCalAttDisable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.00987975 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M8 ;
      ANTENNAMAXAREACAR 2111.65 LAYER M8 ;
    PORT
      LAYER M8 ;
        RECT 36.414 37.892 36.454 37.932 ;
    END
  END csrLsZCalAttDisable
  PIN VIO_ZCalPULoad
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.93455 LAYER M10 ;
    PORT
      LAYER M10 ;
        RECT 100.0285 56.398 104.3275 56.848 ;
    END
  END VIO_ZCalPULoad
  PIN VIO_ZCalPDLoad
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9132 LAYER M10 ;
    PORT
      LAYER M10 ;
        RECT 82.5375 56.398 91.2335 56.848 ;
    END
  END VIO_ZCalPDLoad
  PIN LsZCalAnaClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23237 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0.40017 LAYER M7 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M7 ;
      ANTENNAMAXAREACAR 513.318 LAYER M7 ;
    PORT
      LAYER M6 ;
        RECT 36.614 28.88 36.654 28.918 ;
    END
  END LsZCalAnaClk
  PIN LsZCalAnaEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23096 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 168.886 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.18 36.654 25.22 ;
    END
  END LsZCalAnaEn
  PIN LsZCalCompEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16592 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 134.249 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 24.94 36.654 24.98 ;
    END
  END LsZCalCompEn
  PIN LsZCalCompVOHDAC[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.30006 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 180.617 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 26.78 36.654 26.82 ;
    END
  END LsZCalCompVOHDAC[0]
  PIN LsZCalCompVOHDAC[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23518 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 154.715 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 27.66 36.654 27.7 ;
    END
  END LsZCalCompVOHDAC[1]
  PIN LsZCalCompVOHDAC[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26958 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 163.18 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 27.74 36.654 27.78 ;
    END
  END LsZCalCompVOHDAC[2]
  PIN LsZCalCompVOHDAC[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2338 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 150.318 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 26.46 36.654 26.5 ;
    END
  END LsZCalCompVOHDAC[3]
  PIN LsZCalCompVOHDAC[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16258 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 119.793 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 27.58 36.654 27.62 ;
    END
  END LsZCalCompVOHDAC[4]
  PIN LsZCalCompVOHDAC[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16832 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 118.166 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 27.82 36.654 27.86 ;
    END
  END LsZCalCompVOHDAC[5]
  PIN LsZCalCompVOHDAC[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20421 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 144.661 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.6145 28.18 36.6745 28.24 ;
    END
  END LsZCalCompVOHDAC[6]
  PIN LsZCalDACRangeSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2878 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M8 ;
      ANTENNAMAXAREACAR 532.093 LAYER M8 ;
    PORT
      LAYER M8 ;
        RECT 36.414 37.332 36.454 37.372 ;
    END
  END LsZCalDACRangeSel
  PIN LsZCalPDEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.14174 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 100.553 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.74 36.654 25.78 ;
    END
  END LsZCalPDEn
  PIN LsZCalPUEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.14606 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 104.318 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.34 36.654 25.38 ;
    END
  END LsZCalPUEn
  PIN csrLsZCalCompGainCurrAdj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.30864 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 180.891 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.26 36.654 25.3 ;
    END
  END csrLsZCalCompGainCurrAdj[0]
  PIN csrLsZCalCompGainCurrAdj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27194 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 166.979 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.1 36.654 25.14 ;
    END
  END csrLsZCalCompGainCurrAdj[1]
  PIN csrLsZCalCompGainCurrAdj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23398 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 143.259 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.66 36.654 25.7 ;
    END
  END csrLsZCalCompGainCurrAdj[2]
  PIN csrLsZCalCompGainCurrAdj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.17204 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 123.303 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.58 36.654 25.62 ;
    END
  END csrLsZCalCompGainCurrAdj[3]
  PIN csrLsZCalCompGainCurrAdj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.31353975 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 184.332 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 26.38 36.654 26.42 ;
    END
  END csrLsZCalCompGainCurrAdj[4]
  PIN csrLsZCalCompGainCurrAdj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23834 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 156.798 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.02 36.654 25.06 ;
    END
  END csrLsZCalCompGainCurrAdj[5]
  PIN csrLsZCalCompGainCurrAdj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.24468 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.5 36.654 25.54 ;
    END
  END csrLsZCalCompGainCurrAdj[6]
  PIN csrLsZCalCompGainCurrAdj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16104 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.42 36.654 25.46 ;
    END
  END csrLsZCalCompGainCurrAdj[7]
  PIN csrLsZCalCompVrefDAC[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34138 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 201.573 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 27.34 36.654 27.38 ;
    END
  END csrLsZCalCompVrefDAC[0]
  PIN csrLsZCalCompVrefDAC[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.30328 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 184.455 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 27.42 36.654 27.46 ;
    END
  END csrLsZCalCompVrefDAC[1]
  PIN csrLsZCalCompVrefDAC[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26485975 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 180.788 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 27.9 36.654 27.94 ;
    END
  END csrLsZCalCompVrefDAC[2]
  PIN csrLsZCalCompVrefDAC[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.26166 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 167.528 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 25.82 36.654 25.86 ;
    END
  END csrLsZCalCompVrefDAC[3]
  PIN csrLsZCalCompVrefDAC[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.20566 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 136.465 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 27.5 36.654 27.54 ;
    END
  END csrLsZCalCompVrefDAC[4]
  PIN csrLsZCalCompVrefDAC[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16786 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 125.396 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 26.54 36.654 26.58 ;
    END
  END csrLsZCalCompVrefDAC[5]
  PIN csrLsZCalCompVrefDAC[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.15766 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 114.264 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 36.614 26.7 36.654 26.74 ;
    END
  END csrLsZCalCompVrefDAC[6]
  PIN ZCalCompOut
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.499719 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.041 0.031 33.079 ;
    END
  END ZCalCompOut
  PIN IDDQ_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.654322 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0.023522 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 1.06016 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA6 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.11628 LAYER M6 ;
      ANTENNAGATEAREA 0.11628 LAYER M7 ;
      ANTENNAGATEAREA 0.12239975 LAYER M8 ;
      ANTENNAGATEAREA 0.11628 LAYER VIA6 ;
      ANTENNAGATEAREA 0.11628 LAYER VIA7 ;
      ANTENNAMAXAREACAR 57.6302 LAYER M6 ;
      ANTENNAMAXAREACAR 57.8325 LAYER M7 ;
      ANTENNAMAXAREACAR 147.929 LAYER M8 ;
      ANTENNAMAXCUTCAR 0.567491 LAYER VIA6 ;
      ANTENNAMAXCUTCAR 0.579909 LAYER VIA7 ;
    PORT
      LAYER M6 ;
        RECT 0 36.917 0.038 36.955 ;
    END
  END IDDQ_mode
  PIN BurnIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.39335 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 1.92025 LAYER M7 ;
    ANTENNAPARTIALCUTAREA 0.002888 LAYER VIA6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M7 ;
      ANTENNAMAXAREACAR 1004.15 LAYER M7 ;
    PORT
      LAYER M6 ;
        RECT 0 37.221 0.038 37.259 ;
    END
  END BurnIn
  PIN csrLsTxSlewLPPU1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 319.472 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.047 37.43 145.085 74.71 ;
    END
  END csrLsTxSlewLPPU1[1]
  PIN csrLsTxSlewPD1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 308.815 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.199 37.43 145.237 74.71 ;
    END
  END csrLsTxSlewPD1[1]
  PIN csrLsTxSlewPD1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 314.013 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.123 37.43 145.161 74.71 ;
    END
  END csrLsTxSlewPD1[0]
  PIN csrLsTxSlewLPPU1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 347.754 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 144.895 37.43 144.933 74.71 ;
    END
  END csrLsTxSlewLPPU1[2]
  PIN csrLsTxCalCodeLPPU1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 453.838 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.567 37.43 146.605 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[3]
  PIN csrLsTxCalCodeLPPU1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 429.877 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.643 37.43 146.681 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[4]
  PIN csrLsTxCalCodeLPPU1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 428.826 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.719 37.43 146.757 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[5]
  PIN csrLsTxCalCodeLPPU1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 399.026 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.795 37.43 146.833 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[6]
  PIN csrLsTxCalCodeLPPU1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 378.076 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.947 37.43 146.985 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[8]
  PIN csrLsTxSlewLPPU1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 321.322 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 144.971 37.43 145.009 74.71 ;
    END
  END csrLsTxSlewLPPU1[0]
  PIN TIEHI1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37786 LAYER M6 ;
    ANTENNADIFFAREA 0.00459 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 65.721 0.038 65.759 ;
    END
  END TIEHI1
  PIN TIELO1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37511 LAYER M6 ;
    ANTENNADIFFAREA 0.00918 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 65.873 0.038 65.911 ;
    END
  END TIELO1
  PIN csrLsTxCalCodeLPPU1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 385.675 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.871 37.43 146.909 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[7]
  PIN csrLsTxCalCodeLPPU0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0081 LAYER M7 ;
      ANTENNAMAXAREACAR 385.675 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 146.871 0.05 146.909 37.33 ;
    END
  END csrLsTxCalCodeLPPU0[7]
  PIN csrLsTxSlewPD1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41663975 LAYER M7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0054 LAYER M7 ;
      ANTENNAMAXAREACAR 305.882 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 145.275 37.43 145.313 74.71 ;
    END
  END csrLsTxSlewPD1[2]
  OBS
    LAYER M0 SPACING 0 ;
      RECT MASK 1 0 0 194.055 74.76 ;
    LAYER M0 SPACING 0 ;
      RECT MASK 2 0 0 194.055 74.76 ;
    LAYER M1 SPACING 0 ;
      RECT MASK 1 0 0 194.055 74.76 ;
    LAYER M1 SPACING 0 ;
      RECT MASK 2 0 0 194.055 74.76 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 1 0 0 194.055 74.76 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 2 0 0 194.055 74.76 ;
    LAYER M3 SPACING 0 ;
      RECT MASK 1 0 0 194.055 74.76 ;
      RECT MASK 2 0 0 194.055 74.76 ;
    LAYER M5 SPACING 0 ;
      RECT 0 0 194.055 74.76 ;
    LAYER M4 SPACING 0 ;
      RECT MASK 1 0 0 194.055 74.76 ;
      RECT MASK 2 0 0 194.055 74.76 ;
    LAYER M6 SPACING 0 ;
      POLYGON 0 0 0 0.278 0.038 0.278 0.038 0.316 0 0.316 0 0.354 0.038 0.354 0.038 0.392 0 0.392 0 1.197 0.034 1.197 0.034 1.235 0 1.235 0 1.501 0.034 1.501 0.034 1.539 0 1.539 0 1.653 0.034 1.653 0.034 1.691 0 1.691 0 1.957 0.034 1.957 0.034 1.995 0 1.995 0 2.261 0.033 2.261 0.033 2.299 0 2.299 0 2.413 0.033 2.413 0.033 2.451 0 2.451 0 2.717 0.038 2.717 0.038 2.755 0 2.755 0 3.021 0.033 3.021 0.033 3.059 0 3.059 0 3.173 0.033 3.173 0.033 3.211 0 3.211 0 3.477 0.033 3.477 0.033 3.515 0 3.515 0 3.933 0.038 3.933 0.038 3.971 0 3.971 0 4.389 0.038 4.389 0.038 4.427 0 4.427 0 6.061 0.038 6.061 0.038 6.099 0 6.099 0 6.213 0.038 6.213 0.038 6.251 0 6.251 0 15.941 0.038 15.941 0.038 15.979 0 15.979 0 16.777 0.038 16.777 0.038 16.815 0 16.815 0 17.081 0.038 17.081 0.038 17.119 0 17.119 0 18.069 0.038 18.069 0.038 18.107 0 18.107 0 18.297 0.038 18.297 0.038 18.335 0 18.335 0 18.905 0.038 18.905 0.038 18.943 0 18.943 0 18.981 0.038 18.981 0.038 19.019 0 19.019 0 19.361 0.038 19.361 0.038 19.399 0 19.399 0 19.741 0.038 19.741 0.038 19.779 0 19.779 0 19.969 0.038 19.969 0.038 20.007 0 20.007 0 20.273 0.038 20.273 0.038 20.311 0 20.311 0 20.729 0.038 20.729 0.038 20.767 0 20.767 0 30.989 0.038 30.989 0.038 31.027 0 31.027 0 31.217 0.038 31.217 0.038 31.255 0 31.255 0 32.585 0.038 32.585 0.038 32.623 0 32.623 0 32.889 0.038 32.889 0.038 32.927 0 32.927 0 33.041 0.031 33.041 0.031 33.079 0 33.079 0 33.877 0.038 33.877 0.038 33.915 0 33.915 0 34.257 0.038 34.257 0.038 34.295 0 34.295 0 35.473 0.038 35.473 0.038 35.511 0 35.511 0 35.853 0.038 35.853 0.038 35.891 0 35.891 0 36.917 0.038 36.917 0.038 36.955 0 36.955 0 37.221 0.038 37.221 0.038 37.259 0 37.259 0 37.373 0.038 37.373 0.038 37.411 0 37.411 0 37.525 0.038 37.525 0.038 37.563 0 37.563 0 37.601 0.038 37.601 0.038 37.639 0 37.639 0 38.437 0.034 38.437 0.034 38.475 0 38.475 0 38.741 0.034 38.741 0.034 38.779 0 38.779 0 38.893 0.034 38.893 0.034 38.931 0 38.931 0 39.197 0.034 39.197 0.034 39.235 0 39.235 0 39.501 0.033 39.501 0.033 39.539 0 39.539 0 39.653 0.033 39.653 0.033 39.691 0 39.691 0 39.957 0.038 39.957 0.038 39.995 0 39.995 0 40.261 0.033 40.261 0.033 40.299 0 40.299 0 40.413 0.033 40.413 0.033 40.451 0 40.451 0 40.717 0.033 40.717 0.033 40.755 0 40.755 0 41.173 0.038 41.173 0.038 41.211 0 41.211 0 41.629 0.038 41.629 0.038 41.667 0 41.667 0 43.301 0.038 43.301 0.038 43.339 0 43.339 0 43.453 0.038 43.453 0.038 43.491 0 43.491 0 48.925 0.038 48.925 0.038 48.963 0 48.963 0 54.017 0.038 54.017 0.038 54.055 0 54.055 0 54.321 0.038 54.321 0.038 54.359 0 54.359 0 55.309 0.038 55.309 0.038 55.347 0 55.347 0 55.537 0.038 55.537 0.038 55.575 0 55.575 0 56.145 0.038 56.145 0.038 56.183 0 56.183 0 56.221 0.038 56.221 0.038 56.259 0 56.259 0 56.601 0.038 56.601 0.038 56.639 0 56.639 0 56.981 0.038 56.981 0.038 57.019 0 57.019 0 57.209 0.038 57.209 0.038 57.247 0 57.247 0 57.513 0.038 57.513 0.038 57.551 0 57.551 0 57.969 0.038 57.969 0.038 58.007 0 58.007 0 65.721 0.038 65.721 0.038 65.759 0 65.759 0 65.873 0.038 65.873 0.038 65.911 0 65.911 0 68.229 0.038 68.229 0.038 68.267 0 68.267 0 68.457 0.038 68.457 0.038 68.495 0 68.495 0 69.825 0.038 69.825 0.038 69.863 0 69.863 0 70.129 0.038 70.129 0.038 70.167 0 70.167 0 71.117 0.038 71.117 0.038 71.155 0 71.155 0 71.497 0.038 71.497 0.038 71.535 0 71.535 0 72.713 0.038 72.713 0.038 72.751 0 72.751 0 73.093 0.038 73.093 0.038 73.131 0 73.131 0 74.76 194.055 74.76 194.055 28.918 36.614 28.918 36.614 28.88 36.654 28.88 36.654 28.918 194.055 28.918 194.055 28.52 36.614 28.52 36.614 28.48 36.657 28.48 36.657 28.52 194.055 28.52 194.055 28.24 36.6145 28.24 36.6145 28.18 36.6745 28.18 36.6745 28.24 194.055 28.24 194.055 27.94 36.614 27.94 36.614 27.9 36.654 27.9 36.654 27.94 194.055 27.94 194.055 27.86 36.614 27.86 36.614 27.82 36.654 27.82 36.654 27.86 194.055 27.86 194.055 27.78 36.614 27.78 36.614 27.74 36.654 27.74 36.654 27.78 194.055 27.78 194.055 27.7 36.614 27.7 36.614 27.66 36.654 27.66 36.654 27.7 194.055 27.7 194.055 27.62 36.614 27.62 36.614 27.58 36.654 27.58 36.654 27.62 194.055 27.62 194.055 27.54 36.614 27.54 36.614 27.5 36.654 27.5 36.654 27.54 194.055 27.54 194.055 27.46 36.614 27.46 36.614 27.42 36.654 27.42 36.654 27.46 194.055 27.46 194.055 27.38 36.614 27.38 36.614 27.34 36.654 27.34 36.654 27.38 194.055 27.38 194.055 26.82 36.614 26.82 36.614 26.78 36.654 26.78 36.654 26.82 194.055 26.82 194.055 26.74 36.614 26.74 36.614 26.7 36.654 26.7 36.654 26.74 194.055 26.74 194.055 26.58 36.614 26.58 36.614 26.54 36.654 26.54 36.654 26.58 194.055 26.58 194.055 26.5 36.614 26.5 36.614 26.46 36.654 26.46 36.654 26.5 194.055 26.5 194.055 26.42 36.614 26.42 36.614 26.38 36.654 26.38 36.654 26.42 194.055 26.42 194.055 25.86 36.614 25.86 36.614 25.82 36.654 25.82 36.654 25.86 194.055 25.86 194.055 25.78 36.614 25.78 36.614 25.74 36.654 25.74 36.654 25.78 194.055 25.78 194.055 25.7 36.614 25.7 36.614 25.66 36.654 25.66 36.654 25.7 194.055 25.7 194.055 25.62 36.614 25.62 36.614 25.58 36.654 25.58 36.654 25.62 194.055 25.62 194.055 25.54 36.614 25.54 36.614 25.5 36.654 25.5 36.654 25.54 194.055 25.54 194.055 25.46 36.614 25.46 36.614 25.42 36.654 25.42 36.654 25.46 194.055 25.46 194.055 25.38 36.614 25.38 36.614 25.34 36.654 25.34 36.654 25.38 194.055 25.38 194.055 25.3 36.614 25.3 36.614 25.26 36.654 25.26 36.654 25.3 194.055 25.3 194.055 25.22 36.614 25.22 36.614 25.18 36.654 25.18 36.654 25.22 194.055 25.22 194.055 25.14 36.614 25.14 36.614 25.1 36.654 25.1 36.654 25.14 194.055 25.14 194.055 25.06 36.614 25.06 36.614 25.02 36.654 25.02 36.654 25.06 194.055 25.06 194.055 24.98 36.614 24.98 36.614 24.94 36.654 24.94 36.654 24.98 194.055 24.98 194.055 0 ;
    LAYER M7 SPACING 0 ;
      POLYGON 0 0 0 74.76 194.055 74.76 194.055 74.71 144.895 74.71 144.895 37.43 144.933 37.43 144.933 74.71 144.971 74.71 144.971 37.43 145.009 37.43 145.009 74.71 145.047 74.71 145.047 37.43 145.085 37.43 145.085 74.71 145.123 74.71 145.123 37.43 145.161 37.43 145.161 74.71 145.199 74.71 145.199 37.43 145.237 37.43 145.237 74.71 145.275 74.71 145.275 37.43 145.313 37.43 145.313 74.71 145.351 74.71 145.351 37.43 145.389 37.43 145.389 74.71 145.655 74.71 145.655 37.43 145.693 37.43 145.693 74.71 145.731 74.71 145.731 37.43 145.769 37.43 145.769 74.71 145.807 74.71 145.807 37.43 145.845 37.43 145.845 74.71 145.883 74.71 145.883 37.43 145.921 37.43 145.921 74.71 145.959 74.71 145.959 37.43 145.997 37.43 145.997 74.71 146.035 74.71 146.035 37.43 146.073 37.43 146.073 74.71 146.111 74.71 146.111 37.43 146.149 37.43 146.149 74.71 146.187 74.71 146.187 37.43 146.225 37.43 146.225 74.71 146.263 74.71 146.263 37.43 146.301 37.43 146.301 74.71 146.339 74.71 146.339 37.43 146.377 37.43 146.377 74.71 146.415 74.71 146.415 37.43 146.453 37.43 146.453 74.71 146.491 74.71 146.491 37.43 146.529 37.43 146.529 74.71 146.567 74.71 146.567 37.43 146.605 37.43 146.605 74.71 146.643 74.71 146.643 37.43 146.681 37.43 146.681 74.71 146.719 74.71 146.719 37.43 146.757 37.43 146.757 74.71 146.795 74.71 146.795 37.43 146.833 37.43 146.833 74.71 146.871 74.71 146.871 37.43 146.909 37.43 146.909 74.71 146.947 74.71 146.947 37.43 146.985 37.43 146.985 74.71 194.055 74.71 194.055 37.33 144.591 37.33 144.591 0.05 144.629 0.05 144.629 37.33 144.895 37.33 144.895 0.05 144.933 0.05 144.933 37.33 144.971 37.33 144.971 0.05 145.009 0.05 145.009 37.33 145.047 37.33 145.047 0.05 145.085 0.05 145.085 37.33 145.123 37.33 145.123 0.05 145.161 0.05 145.161 37.33 145.199 37.33 145.199 0.05 145.237 0.05 145.237 37.33 145.275 37.33 145.275 0.05 145.313 0.05 145.313 37.33 145.351 37.33 145.351 0.05 145.389 0.05 145.389 37.33 145.655 37.33 145.655 0.05 145.693 0.05 145.693 37.33 145.731 37.33 145.731 0.05 145.769 0.05 145.769 37.33 145.807 37.33 145.807 0.05 145.845 0.05 145.845 37.33 145.883 37.33 145.883 0.05 145.921 0.05 145.921 37.33 145.959 37.33 145.959 0.05 145.997 0.05 145.997 37.33 146.035 37.33 146.035 0.05 146.073 0.05 146.073 37.33 146.111 37.33 146.111 0.05 146.149 0.05 146.149 37.33 146.187 37.33 146.187 0.05 146.225 0.05 146.225 37.33 146.263 37.33 146.263 0.05 146.301 0.05 146.301 37.33 146.339 37.33 146.339 0.05 146.377 0.05 146.377 37.33 146.415 37.33 146.415 0.05 146.453 0.05 146.453 37.33 146.491 37.33 146.491 0.05 146.529 0.05 146.529 37.33 146.567 37.33 146.567 0.05 146.605 0.05 146.605 37.33 146.643 37.33 146.643 0.05 146.681 0.05 146.681 37.33 146.719 37.33 146.719 0.05 146.757 0.05 146.757 37.33 146.795 37.33 146.795 0.05 146.833 0.05 146.833 37.33 146.871 37.33 146.871 0.05 146.909 0.05 146.909 37.33 146.947 37.33 146.947 0.05 146.985 0.05 146.985 37.33 194.055 37.33 194.055 0 ;
    LAYER M8 SPACING 0 ;
      POLYGON 0 0 0 74.76 194.055 74.76 194.055 38.072 36.414 38.072 36.414 37.992 36.494 37.992 36.494 38.072 194.055 38.072 194.055 37.932 36.414 37.932 36.414 37.892 36.454 37.892 36.454 37.932 194.055 37.932 194.055 37.372 36.414 37.372 36.414 37.332 36.454 37.332 36.454 37.372 194.055 37.372 194.055 0 ;
    LAYER M9 SPACING 0 ;
      RECT 0 0 194.055 74.76 ;
    LAYER M10 SPACING 0 ;
      POLYGON 0 0 0 74.76 194.055 74.76 194.055 73.4585 0.3 73.4585 0.3 72.8585 144.6645 72.8585 144.6645 73.4585 194.055 73.4585 194.055 73.0745 146.721 73.0745 146.721 72.5585 0.3 72.5585 0.3 71.9585 25.5555 71.9585 25.5555 72.5585 30.1505 72.5585 30.1505 71.9585 104.4075 71.9585 104.4075 72.5585 146.721 72.5585 146.721 72.4745 159.2295 72.4745 159.2295 73.0745 159.7625 73.0745 159.7625 72.4745 174.756 72.4745 174.756 73.0745 194.055 73.0745 194.055 72.5995 175.419 72.5995 175.419 72.1745 144.198 72.1745 144.198 71.6585 0.3 71.6585 0.3 71.0585 25.5555 71.0585 25.5555 71.6585 30.1505 71.6585 30.1505 71.0585 104.4075 71.0585 104.4075 71.6585 144.198 71.6585 144.198 71.5745 174.756 71.5745 174.756 72.1745 175.419 72.1745 175.419 72.0415 193.149 72.0415 193.149 72.5995 194.055 72.5995 194.055 71.5915 175.419 71.5915 175.419 71.2745 146.721 71.2745 146.721 70.6745 159.2295 70.6745 159.2295 71.2745 159.7625 71.2745 159.7625 70.6745 174.756 70.6745 174.756 71.2745 175.419 71.2745 175.419 71.0335 183.361 71.0335 183.361 71.5915 183.811 71.5915 183.811 71.0335 193.149 71.0335 193.149 71.5915 194.055 71.5915 194.055 70.6195 0.3 70.6195 0.3 70.0195 36.164 70.0195 36.164 70.6195 36.414 70.6195 36.414 70.0195 144.6645 70.0195 144.6645 70.6195 194.055 70.6195 194.055 70.5295 176.661 70.5295 176.661 70.0795 191.907 70.0795 191.907 70.5295 194.055 70.5295 194.055 69.5755 175.419 69.5755 175.419 69.4195 0.3 69.4195 0.3 68.8195 144.6645 68.8195 144.6645 69.4195 175.419 69.4195 175.419 69.0175 184.757 69.0175 184.757 69.5755 185.207 69.5755 185.207 69.0175 193.149 69.0175 193.149 69.5755 194.055 69.5755 194.055 68.8055 160.4665 68.8055 160.4665 68.5195 0.3 68.5195 0.3 67.9195 25.5555 67.9195 25.5555 68.5195 36.414 68.5195 36.414 67.9195 104.4075 67.9195 104.4075 68.5195 160.4665 68.5195 160.4665 68.3555 172.52 68.3555 172.52 68.8055 194.055 68.8055 194.055 68.5135 176.661 68.5135 176.661 68.0635 191.907 68.0635 191.907 68.5135 194.055 68.5135 194.055 67.6195 0.3 67.6195 0.3 67.0195 25.5555 67.0195 25.5555 67.6195 36.414 67.6195 36.414 67.0195 104.4075 67.0195 104.4075 67.6195 194.055 67.6195 194.055 67.5595 175.419 67.5595 175.419 67.235 144.198 67.235 144.198 66.7195 0.3 66.7195 0.3 66.1195 25.5555 66.1195 25.5555 66.7195 36.414 66.7195 36.414 66.1195 104.4075 66.1195 104.4075 66.7195 144.198 66.7195 144.198 66.635 174.756 66.635 174.756 67.235 175.419 67.235 175.419 67.0015 183.361 67.0015 183.361 67.5595 183.811 67.5595 183.811 67.0015 193.149 67.0015 193.149 67.5595 194.055 67.5595 194.055 66.4975 176.661 66.4975 176.661 66.335 144.198 66.335 144.198 65.8195 0.3 65.8195 0.3 65.2195 143.9645 65.2195 143.9645 65.8195 144.198 65.8195 144.198 65.735 174.756 65.735 174.756 66.335 176.661 66.335 176.661 66.0475 191.907 66.0475 191.907 66.4975 194.055 66.4975 194.055 65.5435 175.419 65.5435 175.419 65.435 144.198 65.435 144.198 64.9195 0.3 64.9195 0.3 64.3195 36.164 64.3195 36.164 64.9195 36.414 64.9195 36.414 64.3195 104.4075 64.3195 104.4075 64.9195 144.198 64.9195 144.198 64.835 174.756 64.835 174.756 65.435 175.419 65.435 175.419 64.9855 184.757 64.9855 184.757 65.5435 185.207 65.5435 185.207 64.9855 193.149 64.9855 193.149 65.5435 194.055 65.5435 194.055 64.535 146.721 64.535 146.721 64.0195 0.3 64.0195 0.3 63.4195 104.4075 63.4195 104.4075 64.0195 146.721 64.0195 146.721 63.935 159.2295 63.935 159.2295 64.535 159.7625 64.535 159.7625 63.935 174.756 63.935 174.756 64.535 194.055 64.535 194.055 64.4815 176.661 64.4815 176.661 64.0315 191.907 64.0315 191.907 64.4815 194.055 64.4815 194.055 63.635 146.721 63.635 146.721 63.1195 0.3 63.1195 0.3 62.5195 36.164 62.5195 36.164 63.1195 36.414 63.1195 36.414 62.5195 144.5875 62.5195 144.5875 63.1195 146.721 63.1195 146.721 63.035 174.756 63.035 174.756 63.635 194.055 63.635 194.055 63.5275 175.419 63.5275 175.419 62.9695 183.361 62.9695 183.361 63.5275 183.811 63.5275 183.811 62.9695 193.149 62.9695 193.149 63.5275 194.055 63.5275 194.055 62.735 146.721 62.735 146.721 62.135 159.2295 62.135 159.2295 62.735 159.7625 62.735 159.7625 62.135 174.756 62.135 174.756 62.735 194.055 62.735 194.055 62.4655 176.661 62.4655 176.661 62.0155 191.907 62.0155 191.907 62.4655 194.055 62.4655 194.055 61.9575 104.608 61.9575 104.608 61.8195 0.3 61.8195 0.3 61.2195 34.1535 61.2195 34.1535 61.8195 104.608 61.8195 104.608 61.5505 36.414 61.5505 36.414 60.9705 104.4075 60.9705 104.4075 61.5505 104.608 61.5505 104.608 61.3575 144.5875 61.3575 144.5875 61.9575 194.055 61.9575 194.055 61.6505 146.721 61.6505 146.721 61.0505 159.2295 61.0505 159.2295 61.6505 159.7625 61.6505 159.7625 61.0505 174.756 61.0505 174.756 61.6505 194.055 61.6505 194.055 61.5115 175.419 61.5115 175.419 60.9535 184.757 60.9535 184.757 61.5115 185.207 61.5115 185.207 60.9535 193.149 60.9535 193.149 61.5115 194.055 61.5115 194.055 60.9195 0.3 60.9195 0.3 60.3195 23.561 60.3195 23.561 60.9195 104.608 60.9195 104.608 60.3195 122.5515 60.3195 122.5515 60.9195 194.055 60.9195 194.055 60.7505 146.721 60.7505 146.721 60.2505 36.414 60.2505 36.414 60.0195 0.3 60.0195 0.3 59.4195 23.561 59.4195 23.561 60.0195 36.414 60.0195 36.414 59.6705 104.4075 59.6705 104.4075 60.2505 146.721 60.2505 146.721 60.1505 174.756 60.1505 174.756 60.7505 194.055 60.7505 194.055 60.4495 176.661 60.4495 176.661 60.0195 104.608 60.0195 104.608 59.4195 122.5515 59.4195 122.5515 60.0195 176.661 60.0195 176.661 59.9995 191.907 59.9995 191.907 60.4495 194.055 60.4495 194.055 59.8505 146.721 59.8505 146.721 59.2505 159.2295 59.2505 159.2295 59.8505 159.7625 59.8505 159.7625 59.2505 174.756 59.2505 174.756 59.8505 194.055 59.8505 194.055 59.4955 175.419 59.4955 175.419 59.1195 0.3 59.1195 0.3 58.5195 23.561 58.5195 23.561 59.1195 175.419 59.1195 175.419 58.9505 36.414 58.9505 36.414 58.3705 104.4075 58.3705 104.4075 58.9505 104.608 58.9505 104.608 58.3505 122.5515 58.3505 122.5515 58.9505 175.419 58.9505 175.419 58.9375 183.361 58.9375 183.361 59.4955 183.811 59.4955 183.811 58.9375 193.149 58.9375 193.149 59.4955 194.055 59.4955 194.055 58.4335 176.661 58.4335 176.661 58.2195 0.3 58.2195 0.3 57.6195 34.1535 57.6195 34.1535 58.2195 176.661 58.2195 176.661 57.9835 191.907 57.9835 191.907 58.4335 194.055 58.4335 194.055 57.638 36.414 57.638 36.414 57.058 104.4075 57.058 104.4075 57.638 194.055 57.638 194.055 57.4795 175.419 57.4795 175.419 57.3815 160.4665 57.3815 160.4665 57.0195 0.3 57.0195 0.3 56.4195 36.164 56.4195 36.164 57.0195 160.4665 57.0195 160.4665 56.9315 172.52 56.9315 172.52 57.3815 175.419 57.3815 175.419 56.9215 184.757 56.9215 184.757 57.4795 185.207 57.4795 185.207 56.9215 193.149 56.9215 193.149 57.4795 194.055 57.4795 194.055 56.848 82.5375 56.848 82.5375 56.398 91.2335 56.398 91.2335 56.848 100.0285 56.848 100.0285 56.398 104.3275 56.398 104.3275 56.848 194.055 56.848 194.055 56.4175 176.661 56.4175 176.661 55.9675 191.907 55.9675 191.907 56.4175 194.055 56.4175 194.055 55.839 0.3 55.839 0.3 55.239 6.225 55.239 6.225 55.839 194.055 55.839 194.055 55.811 147.594 55.811 147.594 55.211 174.756 55.211 174.756 55.811 194.055 55.811 194.055 55.4635 175.419 55.4635 175.419 54.939 0.3 54.939 0.3 54.339 104.4075 54.339 104.4075 54.939 175.419 54.939 175.419 54.911 147.5945 54.911 147.5945 54.311 174.7565 54.311 174.7565 54.911 175.419 54.911 175.419 54.9055 183.361 54.9055 183.361 55.4635 183.811 55.4635 183.811 54.9055 193.149 54.9055 193.149 55.4635 194.055 55.4635 194.055 54.4015 176.661 54.4015 176.661 54.039 0.3 54.039 0.3 53.439 6.225 53.439 6.225 54.039 176.661 54.039 176.661 54.011 147.594 54.011 147.594 53.411 174.756 53.411 174.756 54.011 176.661 54.011 176.661 53.9515 191.907 53.9515 191.907 54.4015 194.055 54.4015 194.055 53.4475 175.419 53.4475 175.419 53.3025 6.427 53.3025 6.427 53.0565 0.3 53.0565 0.3 52.4565 6.225 52.4565 6.225 53.0565 6.427 53.0565 6.427 52.7225 106.3105 52.7225 106.3105 53.3025 175.419 53.3025 175.419 53.111 141.8235 53.111 141.8235 53.0565 106.5155 53.0565 106.5155 52.4565 122.5515 52.4565 122.5515 53.0565 141.8235 53.0565 141.8235 52.511 159.2295 52.511 159.2295 53.111 159.7625 53.111 159.7625 52.511 174.756 52.511 174.756 53.111 175.419 53.111 175.419 52.8895 184.757 52.8895 184.757 53.4475 185.207 53.4475 185.207 52.8895 193.149 52.8895 193.149 53.4475 194.055 53.4475 194.055 52.3855 176.661 52.3855 176.661 52.211 141.8235 52.211 141.8235 52.1565 0.3 52.1565 0.3 51.5565 6.225 51.5565 6.225 52.1565 106.5155 52.1565 106.5155 52.0025 6.427 52.0025 6.427 51.4225 106.3105 51.4225 106.3105 52.0025 106.5155 52.0025 106.5155 51.5565 122.5515 51.5565 122.5515 52.1565 141.8235 52.1565 141.8235 51.611 174.756 51.611 174.756 52.211 176.661 52.211 176.661 51.9355 191.907 51.9355 191.907 52.3855 194.055 52.3855 194.055 51.4315 175.419 51.4315 175.419 51.311 141.8235 51.311 141.8235 51.2565 0.3 51.2565 0.3 50.6565 6.225 50.6565 6.225 51.2565 106.574 51.2565 106.574 50.7025 36.414 50.7025 36.414 50.1225 106.3105 50.1225 106.3105 50.7025 106.574 50.7025 106.574 50.6565 122.5515 50.6565 122.5515 51.2565 141.8235 51.2565 141.8235 50.711 159.2295 50.711 159.2295 51.311 159.7625 51.311 159.7625 50.711 174.756 50.711 174.756 51.311 175.419 51.311 175.419 50.8735 183.361 50.8735 183.361 51.4315 183.811 51.4315 183.811 50.8735 193.149 50.8735 193.149 51.4315 194.055 51.4315 194.055 50.3695 176.661 50.3695 176.661 50.2265 141.8235 50.2265 141.8235 50.0565 0.3 50.0565 0.3 49.4565 36.164 49.4565 36.164 50.0565 106.5155 50.0565 106.5155 49.4565 122.5515 49.4565 122.5515 50.0565 141.8235 50.0565 141.8235 49.6265 159.2295 49.6265 159.2295 50.2265 159.7625 50.2265 159.7625 49.6265 174.756 49.6265 174.756 50.2265 176.661 50.2265 176.661 49.9195 191.907 49.9195 191.907 50.3695 194.055 50.3695 194.055 49.4155 175.419 49.4155 175.419 49.3265 141.8235 49.3265 141.8235 49.279 36.414 49.279 36.414 49.1565 0.3 49.1565 0.3 48.5565 6.225 48.5565 6.225 49.1565 36.414 49.1565 36.414 48.829 104.4075 48.829 104.4075 49.279 141.8235 49.279 141.8235 49.1565 104.6155 49.1565 104.6155 48.5565 122.5515 48.5565 122.5515 49.1565 141.8235 49.1565 141.8235 48.7265 174.756 48.7265 174.756 49.3265 175.419 49.3265 175.419 48.8575 184.757 48.8575 184.757 49.4155 185.207 49.4155 185.207 48.8575 193.149 48.8575 193.149 49.4155 194.055 49.4155 194.055 48.4265 141.8235 48.4265 141.8235 48.2565 0.3 48.2565 0.3 47.6565 6.225 47.6565 6.225 48.2565 104.407 48.2565 104.407 47.6565 122.5515 47.6565 122.5515 48.2565 141.8235 48.2565 141.8235 47.8265 159.2295 47.8265 159.2295 48.4265 159.7625 48.4265 159.7625 47.8265 174.756 47.8265 174.756 48.4265 194.055 48.4265 194.055 48.3535 176.661 48.3535 176.661 47.9035 191.907 47.9035 191.907 48.3535 194.055 48.3535 194.055 47.3995 175.419 47.3995 175.419 47.3765 0.3 47.3765 0.3 46.7765 6.225 46.7765 6.225 47.3765 36.414 47.3765 36.414 46.7765 122.5515 46.7765 122.5515 47.3765 175.419 47.3765 175.419 46.8415 183.361 46.8415 183.361 47.3995 183.811 47.3995 183.811 46.8415 193.149 46.8415 193.149 47.3995 194.055 47.3995 194.055 46.4765 0.3 46.4765 0.3 45.8765 122.5515 45.8765 122.5515 46.4765 194.055 46.4765 194.055 46.3375 176.661 46.3375 176.661 45.9575 160.4665 45.9575 160.4665 45.5075 172.52 45.5075 172.52 45.9575 176.661 45.9575 176.661 45.8875 191.907 45.8875 191.907 46.3375 194.055 46.3375 194.055 45.3835 175.419 45.3835 175.419 45.2765 0.3 45.2765 0.3 44.6765 106.3105 44.6765 106.3105 45.2765 106.5155 45.2765 106.5155 44.6765 122.5515 44.6765 122.5515 45.2765 175.419 45.2765 175.419 44.8255 184.757 44.8255 184.757 45.3835 185.207 45.3835 185.207 44.8255 193.149 44.8255 193.149 45.3835 194.055 45.3835 194.055 44.387 141.8235 44.387 141.8235 44.3765 0.3 44.3765 0.3 43.7765 6.225 43.7765 6.225 44.3765 36.414 44.3765 36.414 43.7765 122.5515 43.7765 122.5515 44.3765 141.8235 44.3765 141.8235 43.787 174.756 43.787 174.756 44.387 194.055 44.387 194.055 44.3215 176.661 44.3215 176.661 43.8715 191.907 43.8715 191.907 44.3215 194.055 44.3215 194.055 43.4965 0.3 43.4965 0.3 42.8965 6.225 42.8965 6.225 43.4965 36.414 43.4965 36.414 42.8965 122.5515 42.8965 122.5515 43.4965 194.055 43.4965 194.055 43.487 141.8235 43.487 141.8235 42.887 174.7565 42.887 174.7565 43.487 194.055 43.487 194.055 43.3675 175.419 43.3675 175.419 42.8095 183.361 42.8095 183.361 43.3675 183.811 43.3675 183.811 42.8095 193.149 42.8095 193.149 43.3675 194.055 43.3675 194.055 42.5965 0.3 42.5965 0.3 41.9965 6.225 41.9965 6.225 42.5965 36.414 42.5965 36.414 41.9965 122.5515 41.9965 122.5515 42.5965 194.055 42.5965 194.055 42.587 141.8235 42.587 141.8235 41.987 174.756 41.987 174.756 42.587 194.055 42.587 194.055 42.3055 176.661 42.3055 176.661 41.8555 191.907 41.8555 191.907 42.3055 194.055 42.3055 194.055 41.7165 0.3 41.7165 0.3 41.1165 6.225 41.1165 6.225 41.7165 36.414 41.7165 36.414 41.1165 104.4075 41.1165 104.4075 41.7165 104.6575 41.7165 104.6575 41.1165 122.5515 41.1165 122.5515 41.7165 194.055 41.7165 194.055 41.687 141.8235 41.687 141.8235 41.087 159.2295 41.087 159.2295 41.687 159.7625 41.687 159.7625 41.087 174.756 41.087 174.756 41.687 194.055 41.687 194.055 41.3515 175.419 41.3515 175.419 40.8165 0.3 40.8165 0.3 40.2165 6.225 40.2165 6.225 40.8165 36.414 40.8165 36.414 40.2165 122.5515 40.2165 122.5515 40.8165 175.419 40.8165 175.419 40.7935 184.757 40.7935 184.757 41.3515 185.207 41.3515 185.207 40.7935 193.149 40.7935 193.149 41.3515 194.055 41.3515 194.055 40.787 141.8235 40.787 141.8235 40.187 174.756 40.187 174.756 40.787 194.055 40.787 194.055 40.3435 175.419 40.3435 175.419 39.9365 0.3 39.9365 0.3 39.3365 6.225 39.3365 6.225 39.9365 36.414 39.9365 36.414 39.3365 122.5515 39.3365 122.5515 39.9365 175.419 39.9365 175.419 39.887 141.8235 39.887 141.8235 39.287 159.2295 39.287 159.2295 39.887 159.7625 39.887 159.7625 39.287 174.756 39.287 174.756 39.887 175.419 39.887 175.419 39.7855 193.149 39.7855 193.149 40.3435 194.055 40.3435 194.055 39.0365 0.3 39.0365 0.3 38.4365 6.225 38.4365 6.225 39.0365 36.414 39.0365 36.414 38.4365 122.5515 38.4365 122.5515 39.0365 194.055 39.0365 194.055 38.0775 106.5155 38.0775 106.5155 37.4775 122.5515 37.4775 122.5515 38.0775 194.055 38.0775 194.055 37.1775 106.5155 37.1775 106.5155 36.5775 122.5515 36.5775 122.5515 37.1775 194.055 37.1775 194.055 36.2185 0.3 36.2185 0.3 35.6185 14.994 35.6185 14.994 36.2185 105.842 36.2185 105.842 35.6185 122.5515 35.6185 122.5515 36.2185 194.055 36.2185 194.055 35.6945 141.8235 35.6945 141.8235 35.3215 37.835 35.3215 37.835 35.3185 0.3 35.3185 0.3 34.7185 14.994 34.7185 14.994 35.3185 37.835 35.3185 37.835 34.7215 104.4075 34.7215 104.4075 35.3215 141.8235 35.3215 141.8235 35.3185 104.6575 35.3185 104.6575 34.7185 122.5515 34.7185 122.5515 35.3185 141.8235 35.3185 141.8235 35.0945 159.2295 35.0945 159.2295 35.6945 159.7625 35.6945 159.7625 35.0945 174.756 35.0945 174.756 35.6945 194.055 35.6945 194.055 35.2195 175.419 35.2195 175.419 34.7945 141.8235 34.7945 141.8235 34.4185 0.3 34.4185 0.3 33.8185 25.842 33.8185 25.842 34.4185 36.414 34.4185 36.414 33.8185 122.5515 33.8185 122.5515 34.4185 141.8235 34.4185 141.8235 34.1945 174.756 34.1945 174.756 34.7945 175.419 34.7945 175.419 34.6615 193.149 34.6615 193.149 35.2195 194.055 35.2195 194.055 34.2115 175.419 34.2115 175.419 33.8945 141.8235 33.8945 141.8235 33.3795 0.3 33.3795 0.3 32.7795 122.5515 32.7795 122.5515 33.3795 141.8235 33.3795 141.8235 33.2945 159.2295 33.2945 159.2295 33.8945 159.7625 33.8945 159.7625 33.2945 174.756 33.2945 174.756 33.8945 175.419 33.8945 175.419 33.6535 183.361 33.6535 183.361 34.2115 183.811 34.2115 183.811 33.6535 193.149 33.6535 193.149 34.2115 194.055 34.2115 194.055 33.1495 176.661 33.1495 176.661 32.6995 191.907 32.6995 191.907 33.1495 194.055 33.1495 194.055 32.1955 175.419 32.1955 175.419 32.1795 0.3 32.1795 0.3 31.5795 122.5515 31.5795 122.5515 32.1795 175.419 32.1795 175.419 31.6375 184.757 31.6375 184.757 32.1955 185.207 32.1955 185.207 31.6375 193.149 31.6375 193.149 32.1955 194.055 32.1955 194.055 31.4255 160.4665 31.4255 160.4665 31.2795 0.3 31.2795 0.3 30.6795 104.4075 30.6795 104.4075 31.2795 104.6575 31.2795 104.6575 30.6795 122.5515 30.6795 122.5515 31.2795 160.4665 31.2795 160.4665 30.9755 172.52 30.9755 172.52 31.4255 194.055 31.4255 194.055 31.1335 176.661 31.1335 176.661 30.6835 191.907 30.6835 191.907 31.1335 194.055 31.1335 194.055 30.3795 0.3 30.3795 0.3 29.7795 122.5515 29.7795 122.5515 30.3795 194.055 30.3795 194.055 30.1795 175.419 30.1795 175.419 29.855 141.8235 29.855 141.8235 29.4795 0.3 29.4795 0.3 28.8795 14.331 28.8795 14.331 29.4795 104.6565 29.4795 104.6565 28.8795 122.5515 28.8795 122.5515 29.4795 141.8235 29.4795 141.8235 29.255 174.756 29.255 174.756 29.855 175.419 29.855 175.419 29.6215 183.361 29.6215 183.361 30.1795 183.811 30.1795 183.811 29.6215 193.149 29.6215 193.149 30.1795 194.055 30.1795 194.055 29.1175 176.661 29.1175 176.661 28.955 141.8235 28.955 141.8235 28.5795 0.3 28.5795 0.3 27.9795 122.5515 27.9795 122.5515 28.5795 141.8235 28.5795 141.8235 28.355 174.756 28.355 174.756 28.955 176.661 28.955 176.661 28.6675 191.907 28.6675 191.907 29.1175 194.055 29.1175 194.055 28.1635 175.419 28.1635 175.419 28.055 141.8235 28.055 141.8235 27.6795 0.3 27.6795 0.3 27.0795 104.4075 27.0795 104.4075 27.6795 104.6575 27.6795 104.6575 27.0795 122.5515 27.0795 122.5515 27.6795 141.8235 27.6795 141.8235 27.455 174.756 27.455 174.756 28.055 175.419 28.055 175.419 27.6055 184.757 27.6055 184.757 28.1635 185.207 28.1635 185.207 27.6055 193.149 27.6055 193.149 28.1635 194.055 28.1635 194.055 27.155 141.8235 27.155 141.8235 26.7795 0.3 26.7795 0.3 26.1795 122.5515 26.1795 122.5515 26.7795 141.8235 26.7795 141.8235 26.555 159.2295 26.555 159.2295 27.155 159.7625 27.155 159.7625 26.555 174.756 26.555 174.756 27.155 194.055 27.155 194.055 27.1015 176.661 27.1015 176.661 26.6515 191.907 26.6515 191.907 27.1015 194.055 27.1015 194.055 26.255 142.42 26.255 142.42 25.8795 0.3 25.8795 0.3 25.2795 104.4075 25.2795 104.4075 25.8795 142.42 25.8795 142.42 25.655 174.756 25.655 174.756 26.255 194.055 26.255 194.055 26.1475 175.419 26.1475 175.419 25.5895 183.361 25.5895 183.361 26.1475 183.811 26.1475 183.811 25.5895 193.149 25.5895 193.149 26.1475 194.055 26.1475 194.055 25.355 142.55 25.355 142.55 24.755 159.2295 24.755 159.2295 25.355 159.7625 25.355 159.7625 24.755 174.756 24.755 174.756 25.355 194.055 25.355 194.055 25.0855 176.661 25.0855 176.661 24.6375 36.414 24.6375 36.414 24.5795 0.3 24.5795 0.3 23.9795 36.1665 23.9795 36.1665 24.5795 36.414 24.5795 36.414 24.0575 104.4075 24.0575 104.4075 24.6375 104.6125 24.6375 104.6125 24.0375 122.5515 24.0375 122.5515 24.6375 176.661 24.6375 176.661 24.6355 191.907 24.6355 191.907 25.0855 194.055 25.0855 194.055 24.2705 141.8235 24.2705 141.8235 23.6795 0.3 23.6795 0.3 23.0795 6.225 23.0795 6.225 23.6795 141.8235 23.6795 141.8235 23.6705 159.2295 23.6705 159.2295 24.2705 159.7625 24.2705 159.7625 23.6705 174.756 23.6705 174.756 24.2705 194.055 24.2705 194.055 24.1315 175.419 24.1315 175.419 23.5735 184.757 23.5735 184.757 24.1315 185.207 24.1315 185.207 23.5735 193.149 23.5735 193.149 24.1315 194.055 24.1315 194.055 23.3705 141.8235 23.3705 141.8235 23.3375 29.1195 23.3375 29.1195 22.7795 0.3 22.7795 0.3 22.1795 6.225 22.1795 6.225 22.7795 29.1195 22.7795 29.1195 22.7375 36.1665 22.7375 36.1665 23.3375 36.414 23.3375 36.414 22.7575 104.4075 22.7575 104.4075 23.3375 104.6125 23.3375 104.6125 22.7375 122.5515 22.7375 122.5515 23.3375 141.8235 23.3375 141.8235 22.7705 174.756 22.7705 174.756 23.3705 194.055 23.3705 194.055 23.0695 176.661 23.0695 176.661 22.6195 191.907 22.6195 191.907 23.0695 194.055 23.0695 194.055 22.4705 141.8235 22.4705 141.8235 22.1375 124.627 22.1375 124.627 22.0375 36.414 22.0375 36.414 21.9575 16.3205 21.9575 16.3205 21.8795 0.3 21.8795 0.3 21.2795 14.8105 21.2795 14.8105 21.8795 16.3205 21.8795 16.3205 21.4575 36.1665 21.4575 36.1665 21.9575 36.414 21.9575 36.414 21.4575 104.4075 21.4575 104.4075 22.0375 104.6125 22.0375 104.6125 21.5375 122.5515 21.5375 122.5515 22.0375 124.627 22.0375 124.627 21.5375 141.574 21.5375 141.574 22.1375 141.8235 22.1375 141.8235 21.8705 159.2295 21.8705 159.2295 22.4705 159.7625 22.4705 159.7625 21.8705 174.756 21.8705 174.756 22.4705 194.055 22.4705 194.055 22.1155 175.419 22.1155 175.419 21.5575 183.361 21.5575 183.361 22.1155 183.811 22.1155 183.811 21.5575 193.149 21.5575 193.149 22.1155 194.055 22.1155 194.055 21.0535 176.661 21.0535 176.661 20.9795 0.3 20.9795 0.3 20.3795 146.198 20.3795 146.198 20.9795 176.661 20.9795 176.661 20.6035 191.907 20.6035 191.907 21.0535 194.055 21.0535 194.055 20.0995 175.419 20.0995 175.419 20.0015 160.4665 20.0015 160.4665 19.7795 0.3 19.7795 0.3 19.1795 104.4075 19.1795 104.4075 19.7795 160.4665 19.7795 160.4665 19.5515 172.52 19.5515 172.52 20.0015 175.419 20.0015 175.419 19.5415 184.757 19.5415 184.757 20.0995 185.207 20.0995 185.207 19.5415 193.149 19.5415 193.149 20.0995 194.055 20.0995 194.055 19.0375 176.661 19.0375 176.661 18.9795 36.414 18.9795 36.414 18.8795 6.475 18.8795 6.475 18.599 0.3 18.599 0.3 17.999 6.225 17.999 6.225 18.599 6.475 18.599 6.475 18.2795 12.393 18.2795 12.393 18.8795 12.643 18.8795 12.643 18.2795 29.657 18.2795 29.657 18.8795 36.414 18.8795 36.414 18.3795 104.4075 18.3795 104.4075 18.9795 176.661 18.9795 176.661 18.5875 191.907 18.5875 191.907 19.0375 194.055 19.0375 194.055 18.431 147.594 18.431 147.594 18.1815 120.928 18.1815 120.928 17.9795 6.475 17.9795 6.475 17.699 0.3 17.699 0.3 17.099 6.225 17.099 6.225 17.699 6.475 17.699 6.475 17.3795 12.393 17.3795 12.393 17.9795 12.643 17.9795 12.643 17.3795 25.6785 17.3795 25.6785 17.9795 120.928 17.9795 120.928 17.7315 146.1975 17.7315 146.1975 18.1815 147.594 18.1815 147.594 17.831 174.756 17.831 174.756 18.431 194.055 18.431 194.055 18.0835 175.419 18.0835 175.419 17.531 147.594 17.531 147.594 17.496 120.928 17.496 120.928 17.0795 6.475 17.0795 6.475 16.799 0.3 16.799 0.3 16.199 6.225 16.199 6.225 16.799 6.475 16.799 6.475 16.4795 12.393 16.4795 12.393 17.0795 12.643 17.0795 12.643 16.4795 25.6785 16.4795 25.6785 17.0795 120.928 17.0795 120.928 17.046 146.1975 17.046 146.1975 17.496 147.594 17.496 147.594 16.931 174.7565 16.931 174.7565 17.531 175.419 17.531 175.419 17.5255 183.361 17.5255 183.361 18.0835 183.811 18.0835 183.811 17.5255 193.149 17.5255 193.149 18.0835 194.055 18.0835 194.055 17.0215 176.661 17.0215 176.661 16.631 147.594 16.631 147.594 16.3895 36.414 16.3895 36.414 16.1795 6.4745 16.1795 6.4745 15.8165 0.3 15.8165 0.3 15.2165 6.225 15.2165 6.225 15.8165 6.4745 15.8165 6.4745 15.5795 17.2005 15.5795 17.2005 16.1795 17.47 16.1795 17.47 15.5795 25.6785 15.5795 25.6785 16.1795 36.414 16.1795 36.414 15.8095 146.198 15.8095 146.198 16.3895 147.594 16.3895 147.594 16.031 174.756 16.031 174.756 16.631 176.661 16.631 176.661 16.5715 191.907 16.5715 191.907 17.0215 194.055 17.0215 194.055 16.0675 175.419 16.0675 175.419 15.731 147.594 15.731 147.594 15.131 159.2295 15.131 159.2295 15.731 159.7625 15.731 159.7625 15.131 174.756 15.131 174.756 15.731 175.419 15.731 175.419 15.5095 184.757 15.5095 184.757 16.0675 185.207 16.0675 185.207 15.5095 193.149 15.5095 193.149 16.0675 194.055 16.0675 194.055 15.0895 6.475 15.0895 6.475 14.9165 0.3 14.9165 0.3 14.3165 6.225 14.3165 6.225 14.9165 6.475 14.9165 6.475 14.5095 146.1975 14.5095 146.1975 15.0895 194.055 15.0895 194.055 15.0055 176.661 15.0055 176.661 14.831 147.594 14.831 147.594 14.231 174.756 14.231 174.756 14.831 176.661 14.831 176.661 14.5555 191.907 14.5555 191.907 15.0055 194.055 15.0055 194.055 14.0515 175.419 14.0515 175.419 14.0165 0.3 14.0165 0.3 13.4165 6.225 13.4165 6.225 14.0165 175.419 14.0165 175.419 13.931 147.594 13.931 147.594 13.7895 6.475 13.7895 6.475 13.2095 146.1975 13.2095 146.1975 13.7895 147.594 13.7895 147.594 13.331 159.2295 13.331 159.2295 13.931 159.7625 13.931 159.7625 13.331 174.756 13.331 174.756 13.931 175.419 13.931 175.419 13.4935 183.361 13.4935 183.361 14.0515 183.811 14.0515 183.811 13.4935 193.149 13.4935 193.149 14.0515 194.055 14.0515 194.055 12.9895 176.661 12.9895 176.661 12.8465 147.594 12.8465 147.594 12.8165 0.3 12.8165 0.3 12.2165 25.6785 12.2165 25.6785 12.8165 122.232 12.8165 122.232 12.2165 146.1975 12.2165 146.1975 12.8165 147.594 12.8165 147.594 12.2465 159.2295 12.2465 159.2295 12.8465 159.7625 12.8465 159.7625 12.2465 174.756 12.2465 174.756 12.8465 176.661 12.8465 176.661 12.5395 191.907 12.5395 191.907 12.9895 194.055 12.9895 194.055 12.0355 175.419 12.0355 175.419 11.9465 147.594 11.9465 147.594 11.9165 0.3 11.9165 0.3 11.3165 6.225 11.3165 6.225 11.9165 125.927 11.9165 125.927 11.3165 146.1975 11.3165 146.1975 11.9165 147.594 11.9165 147.594 11.3465 174.756 11.3465 174.756 11.9465 175.419 11.9465 175.419 11.4775 184.757 11.4775 184.757 12.0355 185.207 12.0355 185.207 11.4775 193.149 11.4775 193.149 12.0355 194.055 12.0355 194.055 11.0465 147.594 11.0465 147.594 11.0165 0.3 11.0165 0.3 10.4165 6.225 10.4165 6.225 11.0165 125.8405 11.0165 125.8405 10.4165 146.1975 10.4165 146.1975 11.0165 147.594 11.0165 147.594 10.4465 159.2295 10.4465 159.2295 11.0465 159.7625 11.0465 159.7625 10.4465 174.756 10.4465 174.756 11.0465 194.055 11.0465 194.055 10.9735 176.661 10.9735 176.661 10.5235 191.907 10.5235 191.907 10.9735 194.055 10.9735 194.055 10.1365 0.3 10.1365 0.3 9.5365 146.1975 9.5365 146.1975 10.1365 194.055 10.1365 194.055 10.0195 175.419 10.0195 175.419 9.4615 183.361 9.4615 183.361 10.0195 183.811 10.0195 183.811 9.4615 193.149 9.4615 193.149 10.0195 194.055 10.0195 194.055 9.2365 0.3 9.2365 0.3 8.6365 146.1975 8.6365 146.1975 9.2365 194.055 9.2365 194.055 8.9575 176.661 8.9575 176.661 8.5775 160.4665 8.5775 160.4665 8.1275 172.52 8.1275 172.52 8.5775 176.661 8.5775 176.661 8.5075 191.907 8.5075 191.907 8.9575 194.055 8.9575 194.055 8.0365 0.3 8.0365 0.3 7.4365 146.1975 7.4365 146.1975 8.0365 194.055 8.0365 194.055 8.0035 175.419 8.0035 175.419 7.4455 184.757 7.4455 184.757 8.0035 185.207 8.0035 185.207 7.4455 193.149 7.4455 193.149 8.0035 194.055 8.0035 194.055 7.1365 0.3 7.1365 0.3 6.5365 146.1975 6.5365 146.1975 7.1365 194.055 7.1365 194.055 7.007 147.594 7.007 147.594 6.407 174.756 6.407 174.756 7.007 194.055 7.007 194.055 6.9415 176.661 6.9415 176.661 6.4915 191.907 6.4915 191.907 6.9415 194.055 6.9415 194.055 6.2565 0.3 6.2565 0.3 5.6565 146.1975 5.6565 146.1975 6.2565 194.055 6.2565 194.055 6.107 147.594 6.107 147.594 5.507 174.7565 5.507 174.7565 6.107 194.055 6.107 194.055 5.9875 175.419 5.9875 175.419 5.4565 36.414 5.4565 36.414 5.3565 0.3 5.3565 0.3 4.7565 6.225 4.7565 6.225 5.3565 36.414 5.3565 36.414 5.0065 146.1975 5.0065 146.1975 5.4565 175.419 5.4565 175.419 5.4295 183.361 5.4295 183.361 5.9875 183.811 5.9875 183.811 5.4295 193.149 5.4295 193.149 5.9875 194.055 5.9875 194.055 5.207 147.594 5.207 147.594 4.607 174.756 4.607 174.756 5.207 194.055 5.207 194.055 4.9255 176.661 4.9255 176.661 4.4765 0.3 4.4765 0.3 3.8765 6.225 3.8765 6.225 4.4765 36.414 4.4765 36.414 3.8765 146.1975 3.8765 146.1975 4.4765 176.661 4.4765 176.661 4.4755 191.907 4.4755 191.907 4.9255 194.055 4.9255 194.055 4.307 147.594 4.307 147.594 3.707 159.2295 3.707 159.2295 4.307 159.7625 4.307 159.7625 3.707 174.756 3.707 174.756 4.307 194.055 4.307 194.055 3.9715 175.419 3.9715 175.419 3.5765 0.3 3.5765 0.3 2.9765 6.225 2.9765 6.225 3.5765 36.414 3.5765 36.414 2.9765 146.1975 2.9765 146.1975 3.5765 175.419 3.5765 175.419 3.4135 184.757 3.4135 184.757 3.9715 185.207 3.9715 185.207 3.4135 193.149 3.4135 193.149 3.9715 194.055 3.9715 194.055 3.407 147.594 3.407 147.594 2.807 174.756 2.807 174.756 3.407 194.055 3.407 194.055 2.9635 175.419 2.9635 175.419 2.6965 0.3 2.6965 0.3 2.0965 6.225 2.0965 6.225 2.6965 36.414 2.6965 36.414 2.0965 146.1975 2.0965 146.1975 2.6965 175.419 2.6965 175.419 2.507 147.594 2.507 147.594 1.907 159.2295 1.907 159.2295 2.507 159.7625 2.507 159.7625 1.907 174.756 1.907 174.756 2.507 175.419 2.507 175.419 2.4055 193.149 2.4055 193.149 2.9635 194.055 2.9635 194.055 1.7965 0.3 1.7965 0.3 1.1965 146.1975 1.1965 146.1975 1.7965 194.055 1.7965 194.055 0.5965 0.3 0.5965 0.3 0.1465 146.1975 0.1465 146.1975 0.5965 194.055 0.5965 194.055 0 ;
  END
END dwc_lpddr5xphy_zcalio_ew

END LIBRARY
