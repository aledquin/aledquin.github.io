# LEF OUT API 
# Creation Date : Thu Dec 16 05:51:21 PST 2021
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_txrxdq_ns
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_txrxdq_ns 0 0 ;
  SYMMETRY X Y ;
  SIZE 38.16 BY 297 ;
  PIN DlySweepOut
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66536 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.76146 LAYER D6 ;
    ANTENNADIFFAREA 0.025272 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 18.17 0 18.25 0.08 ;
    END
  END DlySweepOut
  PIN DlySweepIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.33048 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.00798 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1071.91 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2470.1 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 18.46 0 18.54 0.08 ;
    END
  END DlySweepIn
  PIN CsrVrefDAC3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 22.868 75.21125 22.9 97.725 ;
    END
  END CsrVrefDAC3[6]
  PIN CsrVrefDAC3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 22.508 75.21125 22.54 97.725 ;
    END
  END CsrVrefDAC3[5]
  PIN CsrVrefDAC3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 22.148 75.21125 22.18 97.725 ;
    END
  END CsrVrefDAC3[4]
  PIN CsrVrefDAC3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 21.788 75.21125 21.82 97.725 ;
    END
  END CsrVrefDAC3[3]
  PIN CsrVrefDAC3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 21.428 75.21125 21.46 97.725 ;
    END
  END CsrVrefDAC3[2]
  PIN CsrVrefDAC3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 21.068 75.21125 21.1 97.725 ;
    END
  END CsrVrefDAC3[1]
  PIN CsrVrefDAC3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 562.248 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1274.6 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 20.708 75.21125 20.74 97.725 ;
    END
  END CsrVrefDAC3[0]
  PIN CsrVrefDAC2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 19.748 75.21125 19.78 97.702 ;
    END
  END CsrVrefDAC2[6]
  PIN CsrVrefDAC2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 19.388 75.21125 19.42 97.702 ;
    END
  END CsrVrefDAC2[5]
  PIN CsrVrefDAC2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 19.028 75.21125 19.06 97.702 ;
    END
  END CsrVrefDAC2[4]
  PIN CsrVrefDAC2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 18.668 75.21125 18.7 97.702 ;
    END
  END CsrVrefDAC2[3]
  PIN CsrVrefDAC2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 18.308 75.21125 18.34 97.702 ;
    END
  END CsrVrefDAC2[2]
  PIN CsrVrefDAC2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 564.47 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1281.26 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 17.948 75.21125 17.98 97.702 ;
    END
  END CsrVrefDAC2[1]
  PIN CsrVrefDAC2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7204399375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62329 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 562.248 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1274.6 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 17.588 75.21125 17.62 97.702 ;
    END
  END CsrVrefDAC2[0]
  PIN CsrVrefDAC1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7962479375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.79386 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 649.405 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1485.69 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 23.9105 75.21125 23.9425 98.6365 ;
    END
  END CsrVrefDAC1[6]
  PIN CsrVrefDAC1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79164 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.78349 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 647.849 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1485.69 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 23.8385 75.21125 23.8705 98.6365 ;
    END
  END CsrVrefDAC1[5]
  PIN CsrVrefDAC1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.771864 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.739 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 636.534 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1464.03 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 23.7665 75.21125 23.7985 98.6365 ;
    END
  END CsrVrefDAC1[4]
  PIN CsrVrefDAC1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7734 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.74245 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 640.831 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1476.69 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 23.6345 75.21125 23.6665 98.6365 ;
    END
  END CsrVrefDAC1[3]
  PIN CsrVrefDAC1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.790104 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.78004 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 660.442 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1525.03 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 23.5625 75.21125 23.5945 98.6365 ;
    END
  END CsrVrefDAC1[2]
  PIN CsrVrefDAC1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.794712 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.79041 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 672.664 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1557.03 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 23.4905 75.21125 23.5225 98.6365 ;
    END
  END CsrVrefDAC1[1]
  PIN CsrVrefDAC1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.780792 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.75909 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 657.529 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1525.51 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 23.4185 75.21125 23.4505 98.6365 ;
    END
  END CsrVrefDAC1[0]
  PIN CsrVrefDAC0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.798808 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.79962 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 691.38 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1609.03 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.6455 75.21125 16.6775 98.6365 ;
    END
  END CsrVrefDAC0[6]
  PIN CsrVrefDAC0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.797512 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.79671 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 680.898 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1579.22 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.7175 75.21125 16.7495 98.6365 ;
    END
  END CsrVrefDAC0[5]
  PIN CsrVrefDAC0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79484 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7906899375 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 669.355 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1547.03 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.7895 75.21125 16.8215 98.6365 ;
    END
  END CsrVrefDAC0[4]
  PIN CsrVrefDAC0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.793176 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.78695 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 657.849 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1514.14 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.9215 75.21125 16.9535 98.6365 ;
    END
  END CsrVrefDAC0[3]
  PIN CsrVrefDAC0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79164 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.78349 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 647.553 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1484.81 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.9935 75.21125 17.0255 98.6365 ;
    END
  END CsrVrefDAC0[2]
  PIN CsrVrefDAC0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.780792 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.75909 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 623.677 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1423.96 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 17.0655 75.21125 17.0975 98.6365 ;
    END
  END CsrVrefDAC0[1]
  PIN CsrVrefDAC0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.790104 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.78004 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 629.257 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1431.47 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 17.1375 75.21125 17.1695 98.6365 ;
    END
  END CsrVrefDAC0[0]
  PIN CsrSelAnalogVref
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.737896 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.66257 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 576.458 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1307.12 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 17.468 75.21125 17.5 98.2705 ;
    END
  END CsrSelAnalogVref
  PIN CsrRxCurrAdj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.759192 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.71049 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 619.201 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1421.36 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 24.2585 75.21125 24.2905 98.6365 ;
    END
  END CsrRxCurrAdj[7]
  PIN CsrRxCurrAdj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.763224 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.71956 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 631.529 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1457.68 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 24.1865 75.21125 24.2185 98.6365 ;
    END
  END CsrRxCurrAdj[6]
  PIN CsrRxCurrAdj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.76476 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.72301 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 645.275 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1497.69 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 24.1145 75.21125 24.1465 98.6365 ;
    END
  END CsrRxCurrAdj[5]
  PIN CsrRxCurrAdj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.767832 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.72993 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 661.868 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1544.36 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 24.0425 75.21125 24.0745 98.6365 ;
    END
  END CsrRxCurrAdj[4]
  PIN CsrRxCurrAdj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.76364 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.72049 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 658.752 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1539.11 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.25675 75.21125 16.28875 98.6365 ;
    END
  END CsrRxCurrAdj[3]
  PIN CsrRxCurrAdj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.759192 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.71049 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 643.437 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1494.07 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.32875 75.21125 16.36075 98.6365 ;
    END
  END CsrRxCurrAdj[2]
  PIN CsrRxCurrAdj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.771864 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.739 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 641.465 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1479.07 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.40075 75.21125 16.43275 98.6365 ;
    END
  END CsrRxCurrAdj[1]
  PIN CsrRxCurrAdj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.754872 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.70077 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 613.895 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1406.07 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 16.47275 75.21125 16.50475 98.6365 ;
    END
  END CsrRxCurrAdj[0]
  PIN CsrRxChPowerdown[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74636 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.68161 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 583.748 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1324.1 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 19.868 75.21125 19.9 97.702 ;
    END
  END CsrRxChPowerdown[3]
  PIN CsrRxChPowerdown[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74636 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.68161 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 589.655 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1341.82 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 19.508 75.21125 19.54 97.702 ;
    END
  END CsrRxChPowerdown[2]
  PIN CsrRxChPowerdown[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74636 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.68161 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 585.211 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1328.49 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 18.068 75.21125 18.1 97.702 ;
    END
  END CsrRxChPowerdown[1]
  PIN CsrRxChPowerdown[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74636 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.68161 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 583.507 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1323.37 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 17.708 75.21125 17.74 97.702 ;
    END
  END CsrRxChPowerdown[0]
  PIN CsrExtVrefRange
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7290799375 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.64273 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 591.877 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1358.49 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 20.348 75.21125 20.38 97.995 ;
    END
  END CsrExtVrefRange
  PIN CsrDfeCtrl[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.92056 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0856599375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1274.44 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 4117.02 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 36.62 0 36.7 0.08 ;
    END
  END CsrDfeCtrl[2]
  PIN CsrDfeCtrl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.92696 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.10006 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1244.7 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 3983.95 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 36.475 0 36.555 0.08 ;
    END
  END CsrDfeCtrl[1]
  PIN CsrDfeCtrl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93336 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1144599375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1235.07 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 3929.5 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 36.33 0 36.41 0.08 ;
    END
  END CsrDfeCtrl[0]
  PIN CsrTxChargeCancel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1204.22 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5397.97 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 269.16675 37.98 269.20675 ;
    END
  END CsrTxChargeCancel[3]
  PIN CsrTxChargeCancel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1197.51 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5369.49 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 269.00675 37.98 269.04675 ;
    END
  END CsrTxChargeCancel[2]
  PIN CsrTxChargeCancel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1202.9 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5393.59 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 268.84675 37.98 268.88675 ;
    END
  END CsrTxChargeCancel[1]
  PIN CsrTxChargeCancel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1183.09 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5317.59 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 268.68675 37.98 268.72675 ;
    END
  END CsrTxChargeCancel[0]
  PIN CsrTxCalBaseN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1260.31 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5640.32 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 257.86175 37.98 257.90175 ;
    END
  END CsrTxCalBaseN
  PIN atpg_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.69359 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.590699937 LAYER D6 ;
    ANTENNADIFFAREA 0.324 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0375839375 LAYER D6 ;
      ANTENNAMAXAREACAR 392.79 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 1161.36 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 37.215 0 37.295 0.08 ;
    END
  END atpg_mode
  PIN TxPowerdown[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05656 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14166 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 73.6301 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 222.695 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.6625 0 28.7425 0.08 ;
    END
  END TxPowerdown[1]
  PIN TxPowerdown[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 68.4128 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 198.639 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.5175 0 28.5975 0.08 ;
    END
  END TxPowerdown[0]
  PIN TxEq
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21376 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.49536 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0259199375 LAYER D6 ;
      ANTENNAMAXAREACAR 21.5715 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 60.6776 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.9375 0 28.0175 0.08 ;
    END
  END TxEq
  PIN TxEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.17056 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.39816 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0259199375 LAYER D6 ;
      ANTENNAMAXAREACAR 16.7297 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 48.0424 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.3725 0 28.4525 0.08 ;
    END
  END TxEn
  PIN TxDat
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.04096 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10656 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.020736 LAYER D6 ;
      ANTENNAMAXAREACAR 18.8628 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.302099938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.2275 0 28.3075 0.08 ;
    END
  END TxDat
  PIN TxClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10576 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2523599375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.011664 LAYER D6 ;
      ANTENNAMAXAREACAR 42.9762 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 138.026 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.0825 0 28.1625 0.08 ;
    END
  END TxClk
  PIN RxCoreLoopEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.38968 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.14118 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.047952 LAYER D6 ;
      ANTENNAMAXAREACAR 62.964799937 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 182.141 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 19.185 0 19.265 0.08 ;
    END
  END RxCoreLoopEn
  PIN FlyOverTriTx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D6 ;
      ANTENNAMAXAREACAR 45.7398 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 136.201 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.4625 0 27.5425 0.08 ;
    END
  END FlyOverTriTx
  PIN FlyOverEnTx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09936 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.23796 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 167.9 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 573.042 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 26.5375 0 26.6175 0.08 ;
    END
  END FlyOverEnTx
  PIN FlyOverDataTx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 90.1867 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 269.861 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.3175 0 27.3975 0.08 ;
    END
  END FlyOverDataTx
  PIN Ctlpipe_ODT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18748 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.43623 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D6 ;
      ANTENNAMAXAREACAR 151.155 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 433.289 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.6075 0 27.6875 0.08 ;
    END
  END Ctlpipe_ODT
  PIN CsrTxStrenEqLo480Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05656 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14166 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 63.173299937 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 138.625 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.0275 0 27.1075 0.08 ;
    END
  END CsrTxStrenEqLo480Pu
  PIN CsrTxStrenEqLo480Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.4358 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 72.0312 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.9525 0 29.0325 0.08 ;
    END
  END CsrTxStrenEqLo480Pd
  PIN CsrTxStrenEqLo240Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05656 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14166 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 63.173299937 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 138.625 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.8275 0 25.9075 0.08 ;
    END
  END CsrTxStrenEqLo240Pu
  PIN CsrTxStrenEqLo240Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.3779 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.770799938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 30.1525 0 30.2325 0.08 ;
    END
  END CsrTxStrenEqLo240Pd
  PIN CsrTxStrenEqLo120Pu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 63.0576 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 138.365 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 21.0275 0 21.1075 0.08 ;
    END
  END CsrTxStrenEqLo120Pu[3]
  PIN CsrTxStrenEqLo120Pu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 63.0576 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 138.365 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 22.2275 0 22.3075 0.08 ;
    END
  END CsrTxStrenEqLo120Pu[2]
  PIN CsrTxStrenEqLo120Pu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 63.0576 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 138.365 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 23.4275 0 23.5075 0.08 ;
    END
  END CsrTxStrenEqLo120Pu[1]
  PIN CsrTxStrenEqLo120Pu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 63.0576 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 138.365 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 24.6275 0 24.7075 0.08 ;
    END
  END CsrTxStrenEqLo120Pu[0]
  PIN CsrTxStrenEqLo120Pd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.3779 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.770799938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 34.9525 0 35.0325 0.08 ;
    END
  END CsrTxStrenEqLo120Pd[3]
  PIN CsrTxStrenEqLo120Pd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.3779 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.770799938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.7525 0 33.8325 0.08 ;
    END
  END CsrTxStrenEqLo120Pd[2]
  PIN CsrTxStrenEqLo120Pd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.3779 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.770799938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.5525 0 32.6325 0.08 ;
    END
  END CsrTxStrenEqLo120Pd[1]
  PIN CsrTxStrenEqLo120Pd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.3779 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.770799938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 31.3525 0 31.4325 0.08 ;
    END
  END CsrTxStrenEqLo120Pd[0]
  PIN CsrTxStrenEqHi480Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 65.4696 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 152.125 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 26.3725 0 26.4525 0.08 ;
    END
  END CsrTxStrenEqHi480Pu
  PIN CsrTxStrenEqHi480Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.5202 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.414 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.8075 0 28.8875 0.08 ;
    END
  END CsrTxStrenEqHi480Pd
  PIN CsrTxStrenEqHi240Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 65.4696 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 152.125 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.1725 0 25.2525 0.08 ;
    END
  END CsrTxStrenEqHi240Pu
  PIN CsrTxStrenEqHi240Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.5202 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.414 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 30.0075 0 30.0875 0.08 ;
    END
  END CsrTxStrenEqHi240Pd
  PIN CsrTxStrenEqHi120Pu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 65.4696 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 152.125 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 20.3725 0 20.4525 0.08 ;
    END
  END CsrTxStrenEqHi120Pu[3]
  PIN CsrTxStrenEqHi120Pu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 65.4696 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 152.125 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 21.5725 0 21.6525 0.08 ;
    END
  END CsrTxStrenEqHi120Pu[2]
  PIN CsrTxStrenEqHi120Pu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 65.4696 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 152.125 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 22.7725 0 22.8525 0.08 ;
    END
  END CsrTxStrenEqHi120Pu[1]
  PIN CsrTxStrenEqHi120Pu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 65.4696 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 152.125 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 23.9725 0 24.0525 0.08 ;
    END
  END CsrTxStrenEqHi120Pu[0]
  PIN CsrTxStrenEqHi120Pd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.5202 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.414 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 34.8075 0 34.8875 0.08 ;
    END
  END CsrTxStrenEqHi120Pd[3]
  PIN CsrTxStrenEqHi120Pd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.5202 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.414 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.6075 0 33.6875 0.08 ;
    END
  END CsrTxStrenEqHi120Pd[2]
  PIN CsrTxStrenEqHi120Pd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.5202 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.414 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.4075 0 32.4875 0.08 ;
    END
  END CsrTxStrenEqHi120Pd[1]
  PIN CsrTxStrenEqHi120Pd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 30.5202 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 71.414 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 31.2075 0 31.2875 0.08 ;
    END
  END CsrTxStrenEqHi120Pd[0]
  PIN CsrTxStren480Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 38.9592 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 96.430599938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 26.2275 0 26.3075 0.08 ;
    END
  END CsrTxStren480Pu
  PIN CsrTxStren480Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05656 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14166 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 28.0446 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 66.8592 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 29.6075 0 29.6875 0.08 ;
    END
  END CsrTxStren480Pd
  PIN CsrTxStren240Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 38.9592 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 96.430599938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.0275 0 25.1075 0.08 ;
    END
  END CsrTxStren240Pu
  PIN CsrTxStren240Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05656 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14166 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 28.0446 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 66.8592 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 30.8075 0 30.8875 0.08 ;
    END
  END CsrTxStren240Pd
  PIN CsrTxStren120Pu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 38.9592 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 96.430599938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 20.2275 0 20.3075 0.08 ;
    END
  END CsrTxStren120Pu[3]
  PIN CsrTxStren120Pu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 38.9592 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 96.430599938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 21.4275 0 21.5075 0.08 ;
    END
  END CsrTxStren120Pu[2]
  PIN CsrTxStren120Pu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 38.9592 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 96.430599938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 22.6275 0 22.7075 0.08 ;
    END
  END CsrTxStren120Pu[1]
  PIN CsrTxStren120Pu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 38.9592 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 96.430599938 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 23.8275 0 23.9075 0.08 ;
    END
  END CsrTxStren120Pu[0]
  PIN CsrTxStren120Pd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 28.0025 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 66.7645 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 35.6075 0 35.6875 0.08 ;
    END
  END CsrTxStren120Pd[3]
  PIN CsrTxStren120Pd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 28.0025 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 66.7645 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 34.4075 0 34.4875 0.08 ;
    END
  END CsrTxStren120Pd[2]
  PIN CsrTxStren120Pd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 28.0025 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 66.7645 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.2075 0 33.2875 0.08 ;
    END
  END CsrTxStren120Pd[1]
  PIN CsrTxStren120Pd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05616 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14076 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 28.0025 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 66.7645 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.0075 0 32.0875 0.08 ;
    END
  END CsrTxStren120Pd[0]
  PIN CsrTxOdtStren480Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 36.3059 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 101.615 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.1725 0 27.2525 0.08 ;
    END
  END CsrTxOdtStren480Pu
  PIN CsrTxOdtStren480Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 32.6377 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 87.4758 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 29.7525 0 29.8325 0.08 ;
    END
  END CsrTxOdtStren480Pd
  PIN CsrTxOdtStren240Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 36.3059 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 101.615 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.9725 0 26.0525 0.08 ;
    END
  END CsrTxOdtStren240Pu
  PIN CsrTxOdtStren240Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 32.6377 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 87.4758 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 30.9525 0 31.0325 0.08 ;
    END
  END CsrTxOdtStren240Pd
  PIN CsrTxOdtStren120Pu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 36.3059 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 101.615 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 21.1725 0 21.2525 0.08 ;
    END
  END CsrTxOdtStren120Pu[3]
  PIN CsrTxOdtStren120Pu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 36.3059 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 101.615 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 22.3725 0 22.4525 0.08 ;
    END
  END CsrTxOdtStren120Pu[2]
  PIN CsrTxOdtStren120Pu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 36.3059 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 101.615 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 23.5725 0 23.6525 0.08 ;
    END
  END CsrTxOdtStren120Pu[1]
  PIN CsrTxOdtStren120Pu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 36.3059 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 101.615 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 24.7725 0 24.8525 0.08 ;
    END
  END CsrTxOdtStren120Pu[0]
  PIN CsrTxOdtStren120Pd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 32.6377 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 87.4758 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 35.7525 0 35.8325 0.08 ;
    END
  END CsrTxOdtStren120Pd[3]
  PIN CsrTxOdtStren120Pd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 32.6377 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 87.4758 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 34.5525 0 34.6325 0.08 ;
    END
  END CsrTxOdtStren120Pd[2]
  PIN CsrTxOdtStren120Pd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 32.6377 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 87.4758 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.3525 0 33.4325 0.08 ;
    END
  END CsrTxOdtStren120Pd[1]
  PIN CsrTxOdtStren120Pd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06256 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15516 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 32.6377 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 87.4758 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.1525 0 32.2325 0.08 ;
    END
  END CsrTxOdtStren120Pd[0]
  PIN CsrReserved[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.04096 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10656 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 57.5837 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 179.028 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.6975 0 32.7775 0.08 ;
    END
  END CsrReserved[2]
  PIN CsrReserved[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.04096 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10656 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 69.4159 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 219.694 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 31.8625 0 31.9425 0.08 ;
    END
  END CsrReserved[1]
  PIN CsrReserved[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.04096 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10656 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 69.3834 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 219.389 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 31.624 0 31.704 0.08 ;
    END
  END CsrReserved[0]
  PIN dqrxamptst_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.92056 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0856599375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 349.189 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 1123.45 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 0.91775 0 0.99775 0.08 ;
    END
  END dqrxamptst_en
  PIN dqrxamptst3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.92696 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.10006 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 1.06275 0 1.14275 0.08 ;
    END
  END dqrxamptst3
  PIN dqrxamptst2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90776 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.05686 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 0.40425 0 0.48425 0.08 ;
    END
  END dqrxamptst2
  PIN dqrxamptst1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.27948 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.89323 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 1.315 0 1.395 0.08 ;
    END
  END dqrxamptst1
  PIN dqrxamptst0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91416 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.07126 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 0.54925 0 0.62925 0.08 ;
    END
  END dqrxamptst0
  PIN VREFA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.8 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 6.984 LAYER D8 ;
    ANTENNADIFFAREA 1.0752 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 0.18 143.52275 37.98 144.52275 ;
    END
  END VREFA
  PIN RxStandBy
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90136 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.04246 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1312.77 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 4316.75 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 1.46 0 1.54 0.08 ;
    END
  END RxStandBy
  PIN RxRcvDataOdd
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1481 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.59762 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 1.75 0 1.83 0.08 ;
    END
  END RxRcvDataOdd
  PIN RxRcvDataEven
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93336 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1144599375 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 1.605 0 1.685 0.08 ;
    END
  END RxRcvDataEven
  PIN RxPowerdown
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74636 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.68161 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 612.988 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1411.82 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 23.168 75.21125 23.2 97.725 ;
    END
  END RxPowerdown
  PIN RxPhase[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.32408 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.99358 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1087.83 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2564.24 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 18.605 0 18.685 0.08 ;
    END
  END RxPhase[6]
  PIN RxPhase[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.40248 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.16998 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1146.59 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2718.15 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 18.75 0 18.83 0.08 ;
    END
  END RxPhase[5]
  PIN RxPhase[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4088799375 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.18438 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1152.25 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2729.54 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 18.895 0 18.975 0.08 ;
    END
  END RxPhase[4]
  PIN RxPhase[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41528 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.19878 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1170.84 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2796.1 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 19.04 0 19.12 0.08 ;
    END
  END RxPhase[3]
  PIN RxPhase[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.33048 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.00798 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1103.98 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2628.66 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 19.765 0 19.845 0.08 ;
    END
  END RxPhase[2]
  PIN RxPhase[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.39608 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.15558 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1154.36 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2769.65 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 19.62 0 19.7 0.08 ;
    END
  END RxPhase[1]
  PIN RxPhase[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31128 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.96478 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1108.68 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2700.87 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 19.475 0 19.555 0.08 ;
    END
  END RxPhase[0]
  PIN RxParkOdd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29848 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.93598 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D6 ;
      ANTENNAMAXAREACAR 786.771 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 2400.21 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 36.78 0 36.86 0.08 ;
    END
  END RxParkOdd
  PIN RxParkEven
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30488 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.95038 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D6 ;
      ANTENNAMAXAREACAR 520.432 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 1197.26 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 19.91 0 19.99 0.08 ;
    END
  END RxParkEven
  PIN RxDllClkX
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.93 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5274 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 2122.54 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 1638.83 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 36.23 15.69525 38.16 16.69525 ;
    END
  END RxDllClkX
  PIN RxDllClkOutX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90136 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.04246 LAYER D6 ;
    ANTENNADIFFAREA 0.008424 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 37.65 0 37.73 0.08 ;
    END
  END RxDllClkOutX
  PIN RxDllClkOut
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90776 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.05686 LAYER D6 ;
    ANTENNADIFFAREA 0.008424 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 37.505 0 37.585 0.08 ;
    END
  END RxDllClkOut
  PIN RxDllClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.48798 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 2401.68 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2030.61 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 36.449 18.25925 38.16 19.25925 ;
    END
  END RxDllClk
  PIN RxDFEInit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91416 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.07126 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1295.76 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 4163.52 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 37.36 0 37.44 0.08 ;
    END
  END RxDFEInit
  PIN FlyOverEnRx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.737896 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.66257 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER M4 ;
      ANTENNAMAXAREACAR 578.68 LAYER M4 ;
      ANTENNAMAXSIDEAREACAR 1313.79 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 20.468 75.21125 20.5 98.2705 ;
    END
  END FlyOverEnRx
  PIN FlyOverDataRx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.00536 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.27646 LAYER D6 ;
    ANTENNADIFFAREA 0.033696 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 37.07 0 37.15 0.08 ;
    END
  END FlyOverDataRx
  PIN DlySweepSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29208 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.92158 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 1629.22 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 5063.45 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 36.925 0 37.005 0.08 ;
    END
  END DlySweepSel
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER D8 ;
        RECT 0.18 138.02275 37.98 138.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 154.82275 37.98 155.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 133.82275 37.98 134.62275 ;
        RECT 0.18 129.62275 37.98 130.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 125.42275 37.98 126.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 121.22275 37.98 122.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 5.793 37.98 6.393 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 117.02275 37.98 117.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 112.82275 37.98 113.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 108.62275 37.98 109.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 104.42275 37.98 105.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 36.44125 37.98 37.24125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 33.64125 37.98 34.44125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 30.84125 37.98 31.64125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 28.04125 37.98 28.84125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 25.24125 37.98 26.04125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 22.44125 37.98 23.24125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 19.64125 37.98 20.44125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 17.07725 37.98 17.87725 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 14.51325 37.98 15.31325 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 12.14925 37.98 12.94925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 9.78525 37.98 10.58525 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 66.62275 37.98 67.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 60.24125 37.98 61.04125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 56.04125 37.98 56.84125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 51.84125 37.98 52.64125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 47.64125 37.98 48.44125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 43.44125 37.98 44.24125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 163.354 37.98 164.154 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 169.138 37.98 169.938 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.15225 209.9165 37.98 210.7165 ;
        RECT 0.18 4.393 37.98 4.993 ;
    END
    PORT
      LAYER D8 ;
        RECT 20.18025 63.01275 37.98 63.81275 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 252.0685 37.98 252.8685 ;
        RECT 0.6 249.8585 37.98 250.6585 ;
        RECT 19.16175 243.176 37.98 243.976 ;
        RECT 0.6 240.6165 37.98 241.4165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 254.3215 17.4185 255.1215 ;
        RECT 0.6 247.30225 17.4185 248.10225 ;
        RECT 0.6 238.2165 17.4185 239.0165 ;
        RECT 0.6 234.9115 17.4185 235.7115 ;
        RECT 0.6 228.7165 16.33375 229.5165 ;
        RECT 0.6 226.5115 16.33375 227.3115 ;
        RECT 0.6 215.7165 17.4185 216.5165 ;
        RECT 0.6 212.4165 17.4185 213.2165 ;
        RECT 0.6 204.9165 16.33375 205.7165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 233.7165 37.98 234.5165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 237.1165 37.98 237.9165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 1.593 37.98 2.193 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 231.1165 37.98 231.9165 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.633 282.034 35.583 282.734 ;
        RECT 2.633 279.472 35.583 280.172 ;
        RECT 2.633 276.91 35.583 277.61 ;
        RECT 2.633 274.348 35.583 275.048 ;
        RECT 2.633 271.786 35.583 272.486 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 8.593 37.98 8.993 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 178.238 37.98 179.038 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 180.838 37.98 181.638 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 100.22275 37.98 101.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 97.42275 37.98 98.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 91.82275 37.98 92.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 87.62275 37.98 88.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 83.42275 37.98 84.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 79.22275 37.98 80.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 76.42275 37.98 77.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 73.62275 37.98 74.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 70.82275 37.98 71.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 39.24125 37.98 40.04125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 159.02275 37.98 159.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 150.62275 37.98 151.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 146.42275 37.98 147.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 142.22275 37.98 143.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 198.3165 16.33375 199.1165 ;
        RECT 0.6 173.638 16.33375 174.438 ;
        RECT 0.6 171.438 16.33375 172.238 ;
        RECT 0.6 168.038 16.33375 168.838 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 223.1165 37.98 223.9165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 220.5165 37.98 221.3165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 217.9165 37.98 218.7165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 7.193 37.98 7.793 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 2.993 37.98 3.593 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 207.3165 37.98 208.1165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 203.8165 37.98 204.6165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 268.02675 37.98 268.42675 ;
        RECT 0.6 262.86675 37.98 263.26675 ;
        RECT 0.6 261.32175 37.98 261.72175 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 201.6165 37.98 202.4165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 190.938 37.98 191.738 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 197.038 37.98 197.838 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 194.438 37.98 195.238 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 185.438 37.98 186.238 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 174.738 37.98 175.538 ;
    END
  END VSS
  PIN VSH
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 241.392 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 62.4817 LAYER D8 ;
    ANTENNADIFFAREA 57.633 LAYER D8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 4.80295 LAYER D8 ;
      ANTENNAMAXAREACAR 339.691 LAYER D8 ;
      ANTENNAMAXSIDEAREACAR 237.26 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 0.6 255.643 37.98 256.043 ;
        RECT 0.6 244.781 37.98 245.581 ;
    END
    PORT
      LAYER D8 ;
        RECT 17.054 227.6165 37.98 228.4165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 269.70675 37.98 270.10675 ;
        RECT 0.6 256.78025 37.98 257.58025 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 214.6165 37.98 215.4165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 204.9165 37.98 205.7165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 198.3165 37.98 199.1165 ;
        RECT 0.5205 187.633 37.98 188.433 ;
        RECT 0.6 183.238 37.98 184.038 ;
        RECT 19.16175 171.438 37.98 172.238 ;
    END
  END VSH
  PIN VIO_TIE_LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.35572 LAYER D6 ;
    ANTENNAPARTIALMETALAREA 0.58526 LAYER D7 ;
    ANTENNAPARTIALMETALAREA 0.0576 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4582999375 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.64087 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0864 LAYER D8 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S6 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S7 ;
    ANTENNADIFFAREA 0.16128 LAYER D7 ;
    ANTENNADIFFAREA 0.16128 LAYER S7 ;
    ANTENNADIFFAREA 0.16128 LAYER D8 ;
    PORT
      LAYER D6 ;
        RECT 23.307 257.01175 23.407 270.569 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.51 262.52175 19.75 262.76175 ;
    END
  END VIO_TIE_LO
  PIN VIO_TIE_HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.35572 LAYER D6 ;
    ANTENNAPARTIALMETALAREA 0.61246 LAYER D7 ;
    ANTENNAPARTIALMETALAREA 0.0576 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4582999375 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.76327 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0864 LAYER D8 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S6 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S7 ;
    ANTENNADIFFAREA 0.16128 LAYER D7 ;
    ANTENNADIFFAREA 0.16128 LAYER S7 ;
    ANTENNADIFFAREA 0.16128 LAYER D8 ;
    PORT
      LAYER D6 ;
        RECT 23.007 257.01175 23.107 270.569 ;
    END
    PORT
      LAYER D8 ;
        RECT 18.83 262.52175 19.07 262.76175 ;
    END
  END VIO_TIE_HI
  PIN VIO_PwrOk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.552 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8328 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2016 LAYER D5 ;
      ANTENNAMAXAREACAR 48.9171 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 38.9273 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 0.2 166.354 37.96 166.554 ;
    END
  END VIO_PwrOk
  PIN VIO_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.192 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 3.27456 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 2.338 63.332 19.53 64.332 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.165 293.318 35.995 294.338 ;
        RECT 2.165 290.756 35.995 291.776 ;
        RECT 2.165 288.194 35.995 289.214 ;
        RECT 2.165 285.632 35.995 286.652 ;
        RECT 2.633 280.592 35.583 281.612 ;
        RECT 2.633 278.03 35.583 279.05 ;
        RECT 2.633 275.468 35.583 276.488 ;
        RECT 2.633 272.906 35.583 273.926 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 251.4285 17.012 252.4285 ;
        RECT 2.338 242.568 17.012 243.568 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 224.39725 17.012 225.39725 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 210.266 17.012 211.266 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 189.3045 17.012 190.3045 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 175.058 17.012 176.058 ;
    END
  END VIO_PAD
  PIN VIO_FuncMode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2016 LAYER D7 ;
      ANTENNAMAXAREACAR 9.99107 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 41.3104 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 263.76675 37.98 263.80675 ;
    END
  END VIO_FuncMode
  PIN VIO_ForceLow
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08352 LAYER D6 ;
    ANTENNAPARTIALMETALAREA 0.73298 LAYER D7 ;
    ANTENNAPARTIALMETALAREA 0.0576 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 1.96835 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.30561 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0864 LAYER D8 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S6 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2016 LAYER D7 ;
      ANTENNAGATEAREA 0.2016 LAYER S7 ;
      ANTENNAGATEAREA 0.2016 LAYER D8 ;
      ANTENNAMAXAREACAR 4.31628 LAYER D7 ;
      ANTENNAMAXAREACAR 4.60199 LAYER D8 ;
      ANTENNAMAXSIDEAREACAR 19.042 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 19.4706 LAYER D8 ;
      ANTENNAMAXCUTCAR 0.0536706875 LAYER S7 ;
    PORT
      LAYER D8 ;
        RECT 19.17 262.52175 19.41 262.76175 ;
    END
    PORT
      LAYER D6 ;
        RECT 9.59575 259.73375 9.69575 270.569 ;
    END
  END VIO_ForceLow
  PIN VIO_CsrTxThermP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.6128 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 78.5137 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 265.80675 37.98 265.84675 ;
    END
  END VIO_CsrTxThermP[9]
  PIN VIO_CsrTxThermP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.2655 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 76.1692 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 265.12675 37.98 265.16675 ;
    END
  END VIO_CsrTxThermP[8]
  PIN VIO_CsrTxThermP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.104199937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 76.4377 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 265.04675 37.98 265.08675 ;
    END
  END VIO_CsrTxThermP[7]
  PIN VIO_CsrTxThermP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.674 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 74.5591 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 264.40675 37.98 264.44675 ;
    END
  END VIO_CsrTxThermP[6]
  PIN VIO_CsrTxThermP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.636 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 74.306799938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 264.32675 37.98 264.36675 ;
    END
  END VIO_CsrTxThermP[5]
  PIN VIO_CsrTxThermP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.5832 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 74.0836 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 264.24675 37.98 264.28675 ;
    END
  END VIO_CsrTxThermP[4]
  PIN VIO_CsrTxThermP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.44 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 73.3236 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 264.16675 37.98 264.20675 ;
    END
  END VIO_CsrTxThermP[3]
  PIN VIO_CsrTxThermP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.8139 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.7327 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 268.60675 37.98 268.64675 ;
    END
  END VIO_CsrTxThermP[30]
  PIN VIO_CsrTxThermP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.4617 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 73.1229 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 264.08675 37.98 264.12675 ;
    END
  END VIO_CsrTxThermP[2]
  PIN VIO_CsrTxThermP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.6417 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 78.9464 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 268.52675 37.98 268.56675 ;
    END
  END VIO_CsrTxThermP[29]
  PIN VIO_CsrTxThermP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.9297 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 80.1524 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.88675 37.98 267.92675 ;
    END
  END VIO_CsrTxThermP[28]
  PIN VIO_CsrTxThermP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.7987 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.3488 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.80675 37.98 267.84675 ;
    END
  END VIO_CsrTxThermP[27]
  PIN VIO_CsrTxThermP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.8641 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 78.7014 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.72675 37.98 267.76675 ;
    END
  END VIO_CsrTxThermP[26]
  PIN VIO_CsrTxThermP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.641 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 78.026 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.64675 37.98 267.68675 ;
    END
  END VIO_CsrTxThermP[25]
  PIN VIO_CsrTxThermP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.8657 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 84.1751 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.56675 37.98 267.60675 ;
    END
  END VIO_CsrTxThermP[24]
  PIN VIO_CsrTxThermP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.8522 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 84.186099938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.48675 37.98 267.52675 ;
    END
  END VIO_CsrTxThermP[23]
  PIN VIO_CsrTxThermP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.7995 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 82.793599938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.40675 37.98 267.44675 ;
    END
  END VIO_CsrTxThermP[22]
  PIN VIO_CsrTxThermP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.9226 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 83.2508 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.32675 37.98 267.36675 ;
    END
  END VIO_CsrTxThermP[21]
  PIN VIO_CsrTxThermP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.0786 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 80.5635 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.24675 37.98 267.28675 ;
    END
  END VIO_CsrTxThermP[20]
  PIN VIO_CsrTxThermP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.271 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 72.4332 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 264.00675 37.98 264.04675 ;
    END
  END VIO_CsrTxThermP[1]
  PIN VIO_CsrTxThermP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.6899 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 83.4591 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.16675 37.98 267.20675 ;
    END
  END VIO_CsrTxThermP[19]
  PIN VIO_CsrTxThermP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.572399937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 83.044799938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.08675 37.98 267.12675 ;
    END
  END VIO_CsrTxThermP[18]
  PIN VIO_CsrTxThermP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.486 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 82.7835 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 267.00675 37.98 267.04675 ;
    END
  END VIO_CsrTxThermP[17]
  PIN VIO_CsrTxThermP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.3082 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 81.958 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 266.92675 37.98 266.96675 ;
    END
  END VIO_CsrTxThermP[16]
  PIN VIO_CsrTxThermP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.2789 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 81.740099938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 266.84675 37.98 266.88675 ;
    END
  END VIO_CsrTxThermP[15]
  PIN VIO_CsrTxThermP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.1923 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 81.236599938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 266.76675 37.98 266.80675 ;
    END
  END VIO_CsrTxThermP[14]
  PIN VIO_CsrTxThermP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.8965 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.8012 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 266.12675 37.98 266.16675 ;
    END
  END VIO_CsrTxThermP[13]
  PIN VIO_CsrTxThermP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.8268 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.3787 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 266.04675 37.98 266.08675 ;
    END
  END VIO_CsrTxThermP[12]
  PIN VIO_CsrTxThermP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.7511 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 78.908 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 265.96675 37.98 266.00675 ;
    END
  END VIO_CsrTxThermP[11]
  PIN VIO_CsrTxThermP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.7807 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.154799938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 265.88675 37.98 265.92675 ;
    END
  END VIO_CsrTxThermP[10]
  PIN VIO_CsrTxThermP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.354099937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 72.4352 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 263.92675 37.98 263.96675 ;
    END
  END VIO_CsrTxThermP[0]
  PIN VIO_CsrTxCalBaseP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.1889 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 76.1671 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 263.60675 37.98 263.64675 ;
    END
  END VIO_CsrTxCalBaseP
  PIN VIO_CsrPreDriveMode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.916399937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 75.0438 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 263.84675 37.98 263.88675 ;
    END
  END VIO_CsrPreDriveMode[2]
  PIN VIO_CsrPreDriveMode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.973199937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 75.1849 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 263.68675 37.98 263.72675 ;
    END
  END VIO_CsrPreDriveMode[1]
  PIN VIO_CsrPreDriveMode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3024 LAYER D7 ;
      ANTENNAMAXAREACAR 6.41678 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 25.795899937 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 263.52675 37.98 263.56675 ;
    END
  END VIO_CsrPreDriveMode[0]
  PIN VDS3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.68 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 6.912 LAYER D8 ;
    ANTENNADIFFAREA 2.96654 LAYER D8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.628992 LAYER D8 ;
      ANTENNAMAXAREACAR 355.86 LAYER D8 ;
      ANTENNAMAXSIDEAREACAR 131.143 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 0.18 296.4 37.98 297 ;
    END
  END VDS3
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER D8 ;
        RECT 0.18 156.22275 37.98 157.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 139.42275 37.98 140.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 135.22275 37.98 136.02275 ;
        RECT 0.18 131.02275 37.98 131.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 126.82275 37.98 127.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 122.62275 37.98 123.42275 ;
        RECT 0.18 118.42275 37.98 119.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 114.22275 37.98 115.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 110.02275 37.98 110.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 105.82275 37.98 106.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 65.22275 37.98 66.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 61.64125 37.98 62.44125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 57.44125 37.98 58.24125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 53.24125 37.98 54.04125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 49.04125 37.98 49.84125 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.15225 211.2165 37.98 212.0165 ;
        RECT 0.18 44.84125 37.98 45.64125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 40.64125 37.98 41.44125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 179.538 37.98 180.338 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 176.938 37.98 177.738 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 170.338 16.33375 171.138 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 202.7165 16.33375 203.5165 ;
        RECT 0.6 200.5165 16.33375 201.3165 ;
        RECT 0.6 193.338 16.33375 194.138 ;
        RECT 0.6 186.538 16.33375 187.338 ;
        RECT 0.6 184.338 16.33375 185.138 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.165 294.76 35.995 295.46 ;
        RECT 2.165 292.198 35.995 292.898 ;
        RECT 2.165 289.636 35.995 290.336 ;
        RECT 2.165 287.074 35.995 287.774 ;
        RECT 2.165 284.512 35.995 285.212 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 248.753 37.98 249.553 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 253.1735 37.98 253.9735 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 245.873 37.98 246.673 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 236.0165 37.98 236.8165 ;
        RECT 0.6 232.4165 37.98 233.2165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 262.04175 37.98 262.42175 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 239.3165 37.98 240.1165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 166.938 37.98 167.738 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 172.538 37.98 173.338 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 101.62275 37.98 102.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 98.82275 37.98 99.62275 ;
        RECT 0.18 96.02275 37.98 96.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 93.22275 37.98 94.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 89.02275 37.98 89.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 84.82275 37.98 85.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 80.62275 37.98 81.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 77.82275 37.98 78.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 75.02275 37.98 75.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 72.22275 37.98 73.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 69.42275 37.98 70.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 164.754 37.98 165.554 ;
        RECT 0.18 160.42275 37.98 161.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 152.02275 37.98 152.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 147.82275 37.98 148.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 18.972 225.4165 37.98 226.2165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 227.6165 16.33375 228.4165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 221.8165 37.98 222.6165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 219.2165 37.98 220.0165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 229.8165 37.98 230.6165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 216.8165 37.98 217.6165 ;
        RECT 19.16175 189.833 37.98 190.633 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 208.6165 37.98 209.4165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 206.0165 37.98 206.8165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 199.4165 37.98 200.2165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 213.5165 37.98 214.3165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 266.26675 37.98 266.66675 ;
        RECT 0.6 264.54675 37.98 264.94675 ;
        RECT 0.6 259.96175 37.98 260.36175 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 195.738 37.98 196.538 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 192.238 37.98 193.038 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 182.138 37.98 182.938 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER D8 ;
        RECT 0.18 145.02275 37.98 145.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 140.82275 37.98 141.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 136.62275 37.98 137.42275 ;
        RECT 0.18 132.42275 37.98 133.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 128.22275 37.98 129.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 124.02275 37.98 124.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 119.82275 37.98 120.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 115.62275 37.98 116.42275 ;
        RECT 0.18 111.42275 37.98 112.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 107.22275 37.98 108.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 35.04125 37.98 35.84125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 32.24125 37.98 33.04125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 29.44125 37.98 30.24125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 26.64125 37.98 27.44125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 23.84125 37.98 24.64125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 21.04125 37.98 21.84125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 13.33125 37.98 14.13125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 68.02275 37.98 68.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 58.84125 37.98 59.64125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 54.64125 37.98 55.44125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 50.44125 37.98 51.24125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 46.24125 37.98 47.04125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 42.04125 37.98 42.84125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 10.96725 37.98 11.76725 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 6.493 37.98 7.093 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 5.093 37.98 5.693 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 7.893 37.98 8.493 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 3.693 37.98 4.293 ;
    END
    PORT
      LAYER D8 ;
        RECT 20.18025 64.11775 37.98 64.91775 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16525 254.3215 37.98 255.1215 ;
        RECT 19.16525 250.9635 37.98 251.7635 ;
        RECT 19.16525 247.25975 37.98 248.05975 ;
        RECT 19.16525 241.7165 37.98 242.5165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 234.9165 37.98 235.7165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 238.2165 37.98 239.0165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 2.293 37.98 2.893 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 103.02275 37.98 103.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 94.62275 37.98 95.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 90.42275 37.98 91.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 86.22275 37.98 87.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 82.02275 37.98 82.82275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 37.84125 37.98 38.64125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 161.82275 37.98 162.62275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 157.62275 37.98 158.42275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 153.42275 37.98 154.22275 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 149.22275 37.98 150.02275 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 228.7165 37.98 229.5165 ;
        RECT 19.16175 226.5165 37.98 227.3165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 215.7165 37.98 216.5165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 224.3165 37.98 225.1165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 212.4165 37.98 213.2165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 202.7165 37.98 203.5165 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 200.5165 37.98 201.3165 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 265.30675 37.98 265.70675 ;
        RECT 0.6 259.20175 37.98 259.60175 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 193.338 37.98 194.138 ;
        RECT 19.16175 188.738 37.98 189.538 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 184.338 37.98 185.138 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 186.538 37.98 187.338 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 170.338 37.98 171.138 ;
        RECT 19.16175 168.038 37.98 168.838 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 175.838 37.98 176.638 ;
        RECT 19.16175 173.638 37.98 174.438 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.18 0.893 37.98 1.493 ;
    END
  END VDD
  PIN TIE_LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.64065 LAYER D5 ;
    ANTENNAPARTIALMETALAREA 1.66117 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.612585 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.84003 LAYER D6 ;
    ANTENNAPARTIALCUTAREA 0.0064 LAYER S5 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.383616 LAYER D6 ;
      ANTENNAMAXAREACAR 30.9231 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 53.3299 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 23.607 257.01175 23.707 270.569 ;
    END
    PORT
      LAYER D5 ;
        RECT 20.887 257.31175 24.09025 257.51175 ;
    END
  END TIE_LO
  PIN TIE_HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5552999375 LAYER D5 ;
    ANTENNAPARTIALMETALAREA 1.35572 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.23577 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4582999375 LAYER D6 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S5 ;
    ANTENNADIFFAREA 0.008424 LAYER D5 ;
    ANTENNADIFFAREA 0.008424 LAYER S5 ;
    ANTENNADIFFAREA 0.008424 LAYER D6 ;
    PORT
      LAYER D5 ;
        RECT 20.967 269.75675 24.09025 269.95675 ;
    END
    PORT
      LAYER D6 ;
        RECT 23.907 257.01175 24.007 270.569 ;
    END
  END TIE_HI
  PIN CsrTxThermN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1314.38 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5772.87 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 259.06175 37.98 259.10175 ;
    END
  END CsrTxThermN[9]
  PIN CsrTxThermN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1291.11 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5674.81 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.98175 37.98 259.02175 ;
    END
  END CsrTxThermN[8]
  PIN CsrTxThermN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1251.5 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5628.53 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.90175 37.98 258.94175 ;
    END
  END CsrTxThermN[7]
  PIN CsrTxThermN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1255.63 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5632.66 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.82175 37.98 258.86175 ;
    END
  END CsrTxThermN[6]
  PIN CsrTxThermN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1258.67 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5556.43 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.74175 37.98 258.78175 ;
    END
  END CsrTxThermN[5]
  PIN CsrTxThermN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1266.82 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5684.65 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.66175 37.98 258.70175 ;
    END
  END CsrTxThermN[4]
  PIN CsrTxThermN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1254.64 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5634.13 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.58175 37.98 258.62175 ;
    END
  END CsrTxThermN[3]
  PIN CsrTxThermN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1238.82 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5550.97 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 261.90175 37.98 261.94175 ;
    END
  END CsrTxThermN[30]
  PIN CsrTxThermN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1283.52 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5719.42 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.50175 37.98 258.54175 ;
    END
  END CsrTxThermN[2]
  PIN CsrTxThermN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1234.09 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5552.08 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 261.82175 37.98 261.86175 ;
    END
  END CsrTxThermN[29]
  PIN CsrTxThermN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1252.92 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5580.35 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 261.18175 37.98 261.22175 ;
    END
  END CsrTxThermN[28]
  PIN CsrTxThermN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1254.33 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5579.8 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 261.10175 37.98 261.14175 ;
    END
  END CsrTxThermN[27]
  PIN CsrTxThermN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1263.56 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5612.47 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 261.02175 37.98 261.06175 ;
    END
  END CsrTxThermN[26]
  PIN CsrTxThermN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1273.03 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5636.61 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 260.94175 37.98 260.98175 ;
    END
  END CsrTxThermN[25]
  PIN CsrTxThermN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1191.13 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5341.33 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 260.86175 37.98 260.90175 ;
    END
  END CsrTxThermN[24]
  PIN CsrTxThermN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1247.55 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5579.17 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 260.78175 37.98 260.82175 ;
    END
  END CsrTxThermN[23]
  PIN CsrTxThermN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1235.41 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5503.72 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 260.70175 37.98 260.74175 ;
    END
  END CsrTxThermN[22]
  PIN CsrTxThermN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1255.59 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5596.73 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 260.62175 37.98 260.66175 ;
    END
  END CsrTxThermN[21]
  PIN CsrTxThermN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1249.48 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5590.13 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 260.54175 37.98 260.58175 ;
    END
  END CsrTxThermN[20]
  PIN CsrTxThermN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1236.4 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5527.08 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.42175 37.98 258.46175 ;
    END
  END CsrTxThermN[1]
  PIN CsrTxThermN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1243.39 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5576.03 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 260.46175 37.98 260.50175 ;
    END
  END CsrTxThermN[19]
  PIN CsrTxThermN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1247.13 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5591.42 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 259.78175 37.98 259.82175 ;
    END
  END CsrTxThermN[18]
  PIN CsrTxThermN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1240.21 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5539 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 259.70175 37.98 259.74175 ;
    END
  END CsrTxThermN[17]
  PIN CsrTxThermN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1330.43 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5949.4 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 263.44675 37.98 263.48675 ;
    END
  END CsrTxThermN[16]
  PIN CsrTxThermN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49526 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.73587 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1274.87 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5674.5 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 263.36675 37.9815 263.40675 ;
    END
  END CsrTxThermN[15]
  PIN CsrTxThermN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1345.01 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5796.25 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 257.94175 37.98 257.98175 ;
    END
  END CsrTxThermN[14]
  PIN CsrTxThermN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1318.71 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5748.84 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.02175 37.98 258.06175 ;
    END
  END CsrTxThermN[13]
  PIN CsrTxThermN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1336.95 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5810.76 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.10175 37.98 258.14175 ;
    END
  END CsrTxThermN[12]
  PIN CsrTxThermN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1303.61 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5668.79 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.18175 37.98 258.22175 ;
    END
  END CsrTxThermN[11]
  PIN CsrTxThermN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1326.55 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5785.31 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.26175 37.98 258.30175 ;
    END
  END CsrTxThermN[10]
  PIN CsrTxThermN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1276.72 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5729.31 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 258.34175 37.98 258.38175 ;
    END
  END CsrTxThermN[0]
  PIN CsrTxSrc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 606.455 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2723.3 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 269.56675 37.98 269.60675 ;
    END
  END CsrTxSrc[7]
  PIN CsrTxSrc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 608.794 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2727.03 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 269.48675 37.98 269.52675 ;
    END
  END CsrTxSrc[6]
  PIN CsrTxSrc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 614.789 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2757.18 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 269.40675 37.98 269.44675 ;
    END
  END CsrTxSrc[5]
  PIN CsrTxSrc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 610.997 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2742.82 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 269.32675 37.98 269.36675 ;
    END
  END CsrTxSrc[4]
  PIN CsrTxSrc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 601.531 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2700.86 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 269.24675 37.98 269.28675 ;
    END
  END CsrTxSrc[3]
  PIN CsrTxSrc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 599.259 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2685.22 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 269.08675 37.98 269.12675 ;
    END
  END CsrTxSrc[2]
  PIN CsrTxSrc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 607.318 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2725.79 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 268.92675 37.98 268.96675 ;
    END
  END CsrTxSrc[1]
  PIN CsrTxSrc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 596.986 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2677.44 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 268.76675 37.98 268.80675 ;
    END
  END CsrTxSrc[0]
  OBS
    LAYER M1 SPACING 0 ;
      RECT 0 0 38.16 297 ;
    LAYER M2 SPACING 0 ;
      RECT 0 0 38.16 297 ;
    LAYER M3 SPACING 0 ;
      RECT 0 0 38.16 297 ;
    LAYER M4 SPACING 0 ;
      POLYGON 0 0 0 297 38.16 297 38.16 98.6365 16.25675 98.6365 16.25675 75.21125 16.28875 75.21125 16.28875 98.6365 16.32875 98.6365 16.32875 75.21125 16.36075 75.21125 16.36075 98.6365 16.40075 98.6365 16.40075 75.21125 16.43275 75.21125 16.43275 98.6365 16.47275 98.6365 16.47275 75.21125 16.50475 75.21125 16.50475 98.6365 16.6455 98.6365 16.6455 75.21125 16.6775 75.21125 16.6775 98.6365 16.7175 98.6365 16.7175 75.21125 16.7495 75.21125 16.7495 98.6365 16.7895 98.6365 16.7895 75.21125 16.8215 75.21125 16.8215 98.6365 16.9215 98.6365 16.9215 75.21125 16.9535 75.21125 16.9535 98.6365 16.9935 98.6365 16.9935 75.21125 17.0255 75.21125 17.0255 98.6365 17.0655 98.6365 17.0655 75.21125 17.0975 75.21125 17.0975 98.6365 17.1375 98.6365 17.1375 75.21125 17.1695 75.21125 17.1695 98.6365 23.4185 98.6365 23.4185 98.2705 17.468 98.2705 17.468 75.21125 17.5 75.21125 17.5 98.2705 20.468 98.2705 20.468 97.995 20.348 97.995 20.348 97.702 17.588 97.702 17.588 75.21125 17.62 75.21125 17.62 97.702 17.708 97.702 17.708 75.21125 17.74 75.21125 17.74 97.702 17.948 97.702 17.948 75.21125 17.98 75.21125 17.98 97.702 18.068 97.702 18.068 75.21125 18.1 75.21125 18.1 97.702 18.308 97.702 18.308 75.21125 18.34 75.21125 18.34 97.702 18.668 97.702 18.668 75.21125 18.7 75.21125 18.7 97.702 19.028 97.702 19.028 75.21125 19.06 75.21125 19.06 97.702 19.388 97.702 19.388 75.21125 19.42 75.21125 19.42 97.702 19.508 97.702 19.508 75.21125 19.54 75.21125 19.54 97.702 19.748 97.702 19.748 75.21125 19.78 75.21125 19.78 97.702 19.868 97.702 19.868 75.21125 19.9 75.21125 19.9 97.702 20.348 97.702 20.348 75.21125 20.38 75.21125 20.38 97.995 20.468 97.995 20.468 75.21125 20.5 75.21125 20.5 98.2705 23.4185 98.2705 23.4185 97.725 20.708 97.725 20.708 75.21125 20.74 75.21125 20.74 97.725 21.068 97.725 21.068 75.21125 21.1 75.21125 21.1 97.725 21.428 97.725 21.428 75.21125 21.46 75.21125 21.46 97.725 21.788 97.725 21.788 75.21125 21.82 75.21125 21.82 97.725 22.148 97.725 22.148 75.21125 22.18 75.21125 22.18 97.725 22.508 97.725 22.508 75.21125 22.54 75.21125 22.54 97.725 22.868 97.725 22.868 75.21125 22.9 75.21125 22.9 97.725 23.168 97.725 23.168 75.21125 23.2 75.21125 23.2 97.725 23.4185 97.725 23.4185 75.21125 23.4505 75.21125 23.4505 98.6365 23.4905 98.6365 23.4905 75.21125 23.5225 75.21125 23.5225 98.6365 23.5625 98.6365 23.5625 75.21125 23.5945 75.21125 23.5945 98.6365 23.6345 98.6365 23.6345 75.21125 23.6665 75.21125 23.6665 98.6365 23.7665 98.6365 23.7665 75.21125 23.7985 75.21125 23.7985 98.6365 23.8385 98.6365 23.8385 75.21125 23.8705 75.21125 23.8705 98.6365 23.9105 98.6365 23.9105 75.21125 23.9425 75.21125 23.9425 98.6365 24.0425 98.6365 24.0425 75.21125 24.0745 75.21125 24.0745 98.6365 24.1145 98.6365 24.1145 75.21125 24.1465 75.21125 24.1465 98.6365 24.1865 98.6365 24.1865 75.21125 24.2185 75.21125 24.2185 98.6365 24.2585 98.6365 24.2585 75.21125 24.2905 75.21125 24.2905 98.6365 38.16 98.6365 38.16 0 ;
    LAYER D5 SPACING 0 ;
      RECT 0 0 38.16 75.21125 ;
      RECT 0 80.291 38.16 81.241 ;
      RECT 0 84.921 38.16 85.871 ;
      RECT 0 89.551 38.16 90.501 ;
      RECT 0 94.181 38.16 166.254 ;
      POLYGON 0 166.654 0 297 38.16 297 38.16 269.95675 20.967 269.95675 20.967 269.75675 24.09025 269.75675 24.09025 269.95675 38.16 269.95675 38.16 257.51175 20.887 257.51175 20.887 257.31175 24.09025 257.31175 24.09025 257.51175 38.16 257.51175 38.16 166.654 ;
    LAYER D6 SPACING 0 ;
      POLYGON 0 0 0 297 38.16 297 38.16 270.569 9.59575 270.569 9.59575 259.73375 9.69575 259.73375 9.69575 270.569 23.007 270.569 23.007 257.01175 23.107 257.01175 23.107 270.569 23.307 270.569 23.307 257.01175 23.407 257.01175 23.407 270.569 23.607 270.569 23.607 257.01175 23.707 257.01175 23.707 270.569 23.907 270.569 23.907 257.01175 24.007 257.01175 24.007 270.569 38.16 270.569 38.16 0 37.73 0 37.73 0.08 37.65 0.08 37.65 0 37.585 0 37.585 0.08 37.505 0.08 37.505 0 37.44 0 37.44 0.08 37.36 0.08 37.36 0 37.295 0 37.295 0.08 37.215 0.08 37.215 0 37.15 0 37.15 0.08 37.07 0.08 37.07 0 37.005 0 37.005 0.08 36.925 0.08 36.925 0 36.86 0 36.86 0.08 36.78 0.08 36.78 0 36.7 0 36.7 0.08 36.62 0.08 36.62 0 36.555 0 36.555 0.08 36.475 0.08 36.475 0 36.41 0 36.41 0.08 36.33 0.08 36.33 0 35.8325 0 35.8325 0.08 35.7525 0.08 35.7525 0 35.6875 0 35.6875 0.08 35.6075 0.08 35.6075 0 35.0325 0 35.0325 0.08 34.9525 0.08 34.9525 0 34.8875 0 34.8875 0.08 34.8075 0.08 34.8075 0 34.6325 0 34.6325 0.08 34.5525 0.08 34.5525 0 34.4875 0 34.4875 0.08 34.4075 0.08 34.4075 0 33.8325 0 33.8325 0.08 33.7525 0.08 33.7525 0 33.6875 0 33.6875 0.08 33.6075 0.08 33.6075 0 33.4325 0 33.4325 0.08 33.3525 0.08 33.3525 0 33.2875 0 33.2875 0.08 33.2075 0.08 33.2075 0 32.7775 0 32.7775 0.08 32.6975 0.08 32.6975 0 32.6325 0 32.6325 0.08 32.5525 0.08 32.5525 0 32.4875 0 32.4875 0.08 32.4075 0.08 32.4075 0 32.2325 0 32.2325 0.08 32.1525 0.08 32.1525 0 32.0875 0 32.0875 0.08 32.0075 0.08 32.0075 0 31.9425 0 31.9425 0.08 31.8625 0.08 31.8625 0 31.704 0 31.704 0.08 31.624 0.08 31.624 0 31.4325 0 31.4325 0.08 31.3525 0.08 31.3525 0 31.2875 0 31.2875 0.08 31.2075 0.08 31.2075 0 31.0325 0 31.0325 0.08 30.9525 0.08 30.9525 0 30.8875 0 30.8875 0.08 30.8075 0.08 30.8075 0 30.2325 0 30.2325 0.08 30.1525 0.08 30.1525 0 30.0875 0 30.0875 0.08 30.0075 0.08 30.0075 0 29.8325 0 29.8325 0.08 29.7525 0.08 29.7525 0 29.6875 0 29.6875 0.08 29.6075 0.08 29.6075 0 29.0325 0 29.0325 0.08 28.9525 0.08 28.9525 0 28.8875 0 28.8875 0.08 28.8075 0.08 28.8075 0 28.7425 0 28.7425 0.08 28.6625 0.08 28.6625 0 28.5975 0 28.5975 0.08 28.5175 0.08 28.5175 0 28.4525 0 28.4525 0.08 28.3725 0.08 28.3725 0 28.3075 0 28.3075 0.08 28.2275 0.08 28.2275 0 28.1625 0 28.1625 0.08 28.0825 0.08 28.0825 0 28.0175 0 28.0175 0.08 27.9375 0.08 27.9375 0 27.6875 0 27.6875 0.08 27.6075 0.08 27.6075 0 27.5425 0 27.5425 0.08 27.4625 0.08 27.4625 0 27.3975 0 27.3975 0.08 27.3175 0.08 27.3175 0 27.2525 0 27.2525 0.08 27.1725 0.08 27.1725 0 27.1075 0 27.1075 0.08 27.0275 0.08 27.0275 0 26.6175 0 26.6175 0.08 26.5375 0.08 26.5375 0 26.4525 0 26.4525 0.08 26.3725 0.08 26.3725 0 26.3075 0 26.3075 0.08 26.2275 0.08 26.2275 0 26.0525 0 26.0525 0.08 25.9725 0.08 25.9725 0 25.9075 0 25.9075 0.08 25.8275 0.08 25.8275 0 25.2525 0 25.2525 0.08 25.1725 0.08 25.1725 0 25.1075 0 25.1075 0.08 25.0275 0.08 25.0275 0 24.8525 0 24.8525 0.08 24.7725 0.08 24.7725 0 24.7075 0 24.7075 0.08 24.6275 0.08 24.6275 0 24.0525 0 24.0525 0.08 23.9725 0.08 23.9725 0 23.9075 0 23.9075 0.08 23.8275 0.08 23.8275 0 23.6525 0 23.6525 0.08 23.5725 0.08 23.5725 0 23.5075 0 23.5075 0.08 23.4275 0.08 23.4275 0 22.8525 0 22.8525 0.08 22.7725 0.08 22.7725 0 22.7075 0 22.7075 0.08 22.6275 0.08 22.6275 0 22.4525 0 22.4525 0.08 22.3725 0.08 22.3725 0 22.3075 0 22.3075 0.08 22.2275 0.08 22.2275 0 21.6525 0 21.6525 0.08 21.5725 0.08 21.5725 0 21.5075 0 21.5075 0.08 21.4275 0.08 21.4275 0 21.2525 0 21.2525 0.08 21.1725 0.08 21.1725 0 21.1075 0 21.1075 0.08 21.0275 0.08 21.0275 0 20.4525 0 20.4525 0.08 20.3725 0.08 20.3725 0 20.3075 0 20.3075 0.08 20.2275 0.08 20.2275 0 19.99 0 19.99 0.08 19.91 0.08 19.91 0 19.845 0 19.845 0.08 19.765 0.08 19.765 0 19.7 0 19.7 0.08 19.62 0.08 19.62 0 19.555 0 19.555 0.08 19.475 0.08 19.475 0 19.265 0 19.265 0.08 19.185 0.08 19.185 0 19.12 0 19.12 0.08 19.04 0.08 19.04 0 18.975 0 18.975 0.08 18.895 0.08 18.895 0 18.83 0 18.83 0.08 18.75 0.08 18.75 0 18.685 0 18.685 0.08 18.605 0.08 18.605 0 18.54 0 18.54 0.08 18.46 0.08 18.46 0 18.25 0 18.25 0.08 18.17 0.08 18.17 0 1.83 0 1.83 0.08 1.75 0.08 1.75 0 1.685 0 1.685 0.08 1.605 0.08 1.605 0 1.54 0 1.54 0.08 1.46 0.08 1.46 0 1.395 0 1.395 0.08 1.315 0.08 1.315 0 1.14275 0 1.14275 0.08 1.06275 0.08 1.06275 0 0.99775 0 0.99775 0.08 0.91775 0.08 0.91775 0 0.62925 0 0.62925 0.08 0.54925 0.08 0.54925 0 0.48425 0 0.48425 0.08 0.40425 0.08 0.40425 0 ;
    LAYER D7 SPACING 0 ;
      RECT 0 0 38.16 15.31325 ;
      RECT 0.18 17.07725 37.98 17.87725 ;
      RECT 0 19.64125 38.16 256.043 ;
      RECT 0 256.78025 38.16 257.58025 ;
      RECT 0.6 259.20175 37.98 259.60175 ;
      POLYGON 37.98 259.957 37.98 260.36175 0.6 260.36175 0.6 259.96175 23.78475 259.96175 23.78475 259.957 ;
      RECT 0.6 261.32175 37.98 261.72175 ;
      RECT 0.6 262.04175 37.98 262.42175 ;
      RECT 1.0855 262.58175 19.41 262.62175 ;
      RECT 19.51 262.58175 34.1415 262.62175 ;
      RECT 18.83 262.66175 34.1415 262.70175 ;
      RECT 0.6 262.86675 37.98 263.26675 ;
      RECT 0.6 264.54675 37.98 264.94675 ;
      POLYGON 37.98 265.302 37.98 265.70675 0.6 265.70675 0.6 265.30675 23.78475 265.30675 23.78475 265.302 ;
      RECT 0.6 266.26675 37.98 266.66675 ;
      RECT 0.6 268.02675 37.98 268.42675 ;
      RECT 0 269.7065 38.16 297 ;
  END
END dwc_ddrphy_txrxdq_ns

END LIBRARY
