# LEF OUT API 
# Creation Date : Wed Jul 15 04:13:24 PDT 2020
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_por
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_por 0 0 ;
  SYMMETRY X Y ;
  SIZE 32.604 BY 27.36 ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 0.3 23.4205 32.304 23.8705 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 26.6905 32.304 27.1405 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 7.9805 32.304 8.4305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 11.1805 32.304 11.6305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 14.3805 32.304 14.8305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 17.5805 32.304 18.0305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 1.5805 32.304 2.0305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 4.7805 32.304 5.2305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 20.0505 32.304 20.5005 ;
    END
  END VDD
  PIN PwrOk_VIO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 32.244 24.3005 32.604 24.6605 ;
    END
    PORT
      LAYER M8 ;
        RECT 24.614 24.2305 32.314 24.7305 ;
    END
  END PwrOk_VIO
  PIN PwrOkDlyd_VIO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M8 ;
        RECT 10.555 19.1905 20.1615 19.6905 ;
    END
    PORT
      LAYER M7 ;
        RECT 14.877 0 15.327 0.45 ;
    END
  END PwrOkDlyd_VIO
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 0.3 12.7805 32.304 13.2305 ;
    END
    PORT
      LAYER M8 ;
        RECT 20.497 19.1905 32.304 19.6905 ;
        RECT 0.3 19.1905 10.1235 19.6905 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 25.0905 32.314 25.5405 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 15.9805 32.304 16.4305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 9.5805 32.304 10.0305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 3.1805 32.304 3.6305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 6.3805 32.304 6.8305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 21.6605 32.304 22.2605 ;
    END
  END VDDQ
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M8 ;
        RECT 0.3 22.6205 32.304 23.0705 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 7.1805 32.304 7.6305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 11.9805 32.304 12.4305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 8.7805 32.304 9.2305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 15.1805 32.304 15.6305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 5.5805 32.304 6.0305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 2.3805 32.304 2.8305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 25.8905 32.304 26.3405 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 3.9805 32.304 4.4305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 16.7805 32.304 17.2305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 13.5805 32.304 14.0305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 10.3805 32.304 10.8305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 20.8505 32.304 21.3005 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 24.2305 24.314 24.7305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 18.3805 32.304 18.8305 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.3 0.7805 32.304 1.2305 ;
    END
  END VSS
  PIN DFTDatSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.5325 27.28 31.6125 27.36 ;
    END
  END DFTDatSel
  PIN ClrPORMemReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.9915 27.28 1.0715 27.36 ;
    END
  END ClrPORMemReset
  PIN MemResetLPullDown_VIO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 29.8905 0 29.9705 0.08 ;
    END
  END MemResetLPullDown_VIO
  PIN MemResetLPullUp_VIO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 27.8275 0 27.9075 0.08 ;
    END
  END MemResetLPullUp_VIO
  PIN DCTMemReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.7915 27.28 30.8715 27.36 ;
    END
  END DCTMemReset
  PIN Reset_X
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 32.1135 27.28 32.1935 27.36 ;
    END
  END Reset_X
  PIN SetDCTSanePulse
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.3725 27.28 31.4525 27.36 ;
    END
  END SetDCTSanePulse
  PIN PwrOk_VMEMP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.4105 27.28 0.4905 27.36 ;
    END
  END PwrOk_VMEMP
  PIN DCTSane
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.9985 27.28 21.0785 27.36 ;
    END
  END DCTSane
  PIN PORMemReset
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.4175 27.28 20.4975 27.36 ;
    END
  END PORMemReset
  PIN PwrOkDlyd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 0 22.8605 0.36 23.2205 ;
    END
  END PwrOkDlyd
  OBS
    LAYER M1 SPACING 0 ;
      RECT 0 0 32.604 27.36 ;
      RECT MASK 1 0.838 0.63 0.918 10.11 ;
      RECT MASK 1 28.062 0.63 28.142 10.11 ;
      RECT MASK 1 1.18 0.635 1.24 0.865 ;
      RECT MASK 1 1.512 0.635 1.572 0.865 ;
      RECT MASK 1 1.844 0.635 1.904 0.865 ;
      RECT MASK 1 2.176 0.635 2.236 0.865 ;
      RECT MASK 1 2.508 0.635 2.568 0.865 ;
      RECT MASK 1 2.84 0.635 2.9 0.865 ;
      RECT MASK 1 3.172 0.635 3.232 0.865 ;
      RECT MASK 1 3.504 0.635 3.564 0.865 ;
      RECT MASK 1 3.836 0.635 3.896 0.865 ;
      RECT MASK 1 4.168 0.635 4.228 0.865 ;
      RECT MASK 1 4.5 0.635 4.56 0.865 ;
      RECT MASK 1 4.832 0.635 4.892 0.865 ;
      RECT MASK 1 5.164 0.635 5.224 0.865 ;
      RECT MASK 1 5.496 0.635 5.556 0.865 ;
      RECT MASK 1 5.828 0.635 5.888 0.865 ;
      RECT MASK 1 6.16 0.635 6.22 0.865 ;
      RECT MASK 1 6.492 0.635 6.552 0.865 ;
      RECT MASK 1 6.824 0.635 6.884 0.865 ;
      RECT MASK 1 7.156 0.635 7.216 0.865 ;
      RECT MASK 1 7.488 0.635 7.548 0.865 ;
      RECT MASK 1 7.82 0.635 7.88 0.865 ;
      RECT MASK 1 8.152 0.635 8.212 0.865 ;
      RECT MASK 1 8.484 0.635 8.544 0.865 ;
      RECT MASK 1 8.816 0.635 8.876 0.865 ;
      RECT MASK 1 9.148 0.635 9.208 0.865 ;
      RECT MASK 1 9.48 0.635 9.54 0.865 ;
      RECT MASK 1 9.812 0.635 9.872 0.865 ;
      RECT MASK 1 10.144 0.635 10.204 0.865 ;
      RECT MASK 1 10.476 0.635 10.536 0.865 ;
      RECT MASK 1 10.808 0.635 10.868 0.865 ;
      RECT MASK 1 11.14 0.635 11.2 0.865 ;
      RECT MASK 1 11.472 0.635 11.532 0.865 ;
      RECT MASK 1 11.804 0.635 11.864 0.865 ;
      RECT MASK 1 12.136 0.635 12.196 0.865 ;
      RECT MASK 1 12.468 0.635 12.528 0.865 ;
      RECT MASK 1 12.8 0.635 12.86 0.865 ;
      RECT MASK 1 13.132 0.635 13.192 0.865 ;
      RECT MASK 1 13.464 0.635 13.524 0.865 ;
      RECT MASK 1 13.796 0.635 13.856 0.865 ;
      RECT MASK 1 14.128 0.635 14.188 0.865 ;
      RECT MASK 1 14.46 0.635 14.52 0.865 ;
      RECT MASK 1 14.792 0.635 14.852 0.865 ;
      RECT MASK 1 15.124 0.635 15.184 0.865 ;
      RECT MASK 1 15.456 0.635 15.516 0.865 ;
      RECT MASK 1 15.954 0.635 16.014 0.865 ;
      RECT MASK 1 16.286 0.635 16.346 0.865 ;
      RECT MASK 1 16.618 0.635 16.678 0.865 ;
      RECT MASK 1 16.95 0.635 17.01 0.865 ;
      RECT MASK 1 17.282 0.635 17.342 0.865 ;
      RECT MASK 1 17.614 0.635 17.674 0.865 ;
      RECT MASK 1 17.946 0.635 18.006 0.865 ;
      RECT MASK 1 18.278 0.635 18.338 0.865 ;
      RECT MASK 1 18.61 0.635 18.67 0.865 ;
      RECT MASK 1 18.942 0.635 19.002 0.865 ;
      RECT MASK 1 19.274 0.635 19.334 0.865 ;
      RECT MASK 1 19.606 0.635 19.666 0.865 ;
      RECT MASK 1 19.938 0.635 19.998 0.865 ;
      RECT MASK 1 20.27 0.635 20.33 0.865 ;
      RECT MASK 1 20.602 0.635 20.662 0.865 ;
      RECT MASK 1 20.934 0.635 20.994 0.865 ;
      RECT MASK 1 21.266 0.635 21.326 0.865 ;
      RECT MASK 1 21.598 0.635 21.658 0.865 ;
      RECT MASK 1 21.93 0.635 21.99 0.865 ;
      RECT MASK 1 22.262 0.635 22.322 0.865 ;
      RECT MASK 1 22.594 0.635 22.654 0.865 ;
      RECT MASK 1 22.926 0.635 22.986 0.865 ;
      RECT MASK 1 23.258 0.635 23.318 0.865 ;
      RECT MASK 1 23.59 0.635 23.65 0.865 ;
      RECT MASK 1 23.922 0.635 23.982 0.865 ;
      RECT MASK 1 24.254 0.635 24.314 0.865 ;
      RECT MASK 1 24.586 0.635 24.646 0.865 ;
      RECT MASK 1 24.918 0.635 24.978 0.865 ;
      RECT MASK 1 25.25 0.635 25.31 0.865 ;
      RECT MASK 1 25.582 0.635 25.642 0.865 ;
      RECT MASK 1 25.914 0.635 25.974 0.865 ;
      RECT MASK 1 26.246 0.635 26.306 0.865 ;
      RECT MASK 1 26.578 0.635 26.638 0.865 ;
      RECT MASK 1 26.91 0.635 26.97 0.865 ;
      RECT MASK 1 27.242 0.635 27.302 0.865 ;
      RECT MASK 1 27.574 0.635 27.634 0.865 ;
      RECT MASK 1 29.591 0.71 29.631 1.11 ;
      RECT MASK 1 29.812 0.71 29.852 1.52 ;
      RECT MASK 1 30.255 0.71 30.295 1.11 ;
      RECT MASK 1 30.476 0.71 30.516 1.52 ;
      RECT MASK 1 30.919 0.71 30.959 1.11 ;
      RECT MASK 1 31.14 0.71 31.18 1.52 ;
      RECT MASK 1 31.583 0.71 31.623 1.11 ;
      RECT MASK 1 31.804 0.765 31.844 1.52 ;
      RECT MASK 1 29.148 0.78 29.188 1.52 ;
      RECT MASK 1 29.372 1.155 29.406 1.875 ;
      RECT MASK 1 30.7 1.155 30.734 1.875 ;
      RECT MASK 1 30.036 1.275 30.07 1.875 ;
      RECT MASK 1 29.591 1.3525 29.631 1.915 ;
      RECT MASK 1 30.255 1.3525 30.295 1.915 ;
      RECT MASK 1 30.919 1.3525 30.959 1.915 ;
      RECT MASK 1 31.583 1.3525 31.623 1.915 ;
      RECT MASK 1 31.364 1.3545 31.398 1.875 ;
      RECT MASK 1 29.148 1.715 29.188 6.33 ;
      RECT MASK 1 29.812 1.715 29.852 6.33 ;
      RECT MASK 1 30.476 1.715 30.516 6.33 ;
      RECT MASK 1 31.14 1.715 31.18 6.33 ;
      RECT MASK 1 31.804 1.715 31.844 6.33 ;
      RECT MASK 1 31.583 2.208 31.623 2.952 ;
      RECT MASK 1 29.591 2.217 29.631 2.926 ;
      RECT MASK 1 30.255 2.217 30.295 2.926 ;
      RECT MASK 1 30.919 2.217 30.959 2.926 ;
      RECT MASK 1 29.369 3.305 29.409 10.135 ;
      RECT MASK 1 29.591 3.305 29.631 7.855 ;
      RECT MASK 1 30.033 3.305 30.073 10.135 ;
      RECT MASK 1 30.255 3.305 30.295 7.855 ;
      RECT MASK 1 30.697 3.305 30.737 10.135 ;
      RECT MASK 1 30.919 3.305 30.959 7.855 ;
      RECT MASK 1 31.361 3.305 31.401 10.135 ;
      RECT MASK 1 31.583 3.305 31.623 7.855 ;
      RECT MASK 1 29.148 6.51 29.188 8.882 ;
      RECT MASK 1 29.812 6.51 29.852 8.882 ;
      RECT MASK 1 30.476 6.51 30.516 8.882 ;
      RECT MASK 1 31.14 6.51 31.18 8.882 ;
      RECT MASK 1 31.804 6.51 31.844 8.882 ;
      RECT MASK 1 29.591 7.985 29.631 10.019 ;
      RECT MASK 1 30.255 7.985 30.295 10.019 ;
      RECT MASK 1 30.919 7.985 30.959 10.019 ;
      RECT MASK 1 31.583 7.985 31.623 10.019 ;
      RECT MASK 1 29.148 9.06 29.188 10.53 ;
      RECT MASK 1 29.812 9.06 29.852 10.53 ;
      RECT MASK 1 30.476 9.06 30.516 10.53 ;
      RECT MASK 1 31.14 9.06 31.18 10.53 ;
      RECT MASK 1 31.804 9.06 31.844 10.53 ;
      RECT MASK 1 26.91 9.1995 26.97 10.105 ;
      RECT MASK 1 27.242 9.1995 27.302 10.105 ;
      RECT MASK 1 7.986 9.505 8.046 14.285 ;
      RECT MASK 1 1.346 9.875 1.406 10.105 ;
      RECT MASK 1 1.678 9.875 1.738 10.105 ;
      RECT MASK 1 2.01 9.875 2.07 10.105 ;
      RECT MASK 1 2.342 9.875 2.402 10.105 ;
      RECT MASK 1 2.674 9.875 2.734 10.105 ;
      RECT MASK 1 3.006 9.875 3.066 10.105 ;
      RECT MASK 1 3.338 9.875 3.398 10.105 ;
      RECT MASK 1 3.67 9.875 3.73 10.105 ;
      RECT MASK 1 4.666 9.875 4.726 10.105 ;
      RECT MASK 1 4.998 9.875 5.058 10.105 ;
      RECT MASK 1 5.33 9.875 5.39 10.105 ;
      RECT MASK 1 5.662 9.875 5.722 10.105 ;
      RECT MASK 1 5.994 9.875 6.054 10.105 ;
      RECT MASK 1 6.326 9.875 6.386 10.105 ;
      RECT MASK 1 6.658 9.875 6.718 10.105 ;
      RECT MASK 1 6.99 9.875 7.05 10.105 ;
      RECT MASK 1 7.322 9.875 7.382 10.105 ;
      RECT MASK 1 7.654 9.875 7.714 10.105 ;
      RECT MASK 1 8.484 9.875 8.544 10.105 ;
      RECT MASK 1 8.816 9.875 8.876 10.105 ;
      RECT MASK 1 9.148 9.875 9.208 10.105 ;
      RECT MASK 1 9.48 9.875 9.54 10.105 ;
      RECT MASK 1 9.812 9.875 9.872 10.105 ;
      RECT MASK 1 10.144 9.875 10.204 10.105 ;
      RECT MASK 1 10.476 9.875 10.536 10.105 ;
      RECT MASK 1 10.808 9.875 10.868 10.105 ;
      RECT MASK 1 11.14 9.875 11.2 10.105 ;
      RECT MASK 1 11.472 9.875 11.532 10.105 ;
      RECT MASK 1 11.804 9.875 11.864 10.105 ;
      RECT MASK 1 12.136 9.875 12.196 10.105 ;
      RECT MASK 1 12.468 9.875 12.528 10.105 ;
      RECT MASK 1 12.8 9.875 12.86 10.105 ;
      RECT MASK 1 13.132 9.875 13.192 10.105 ;
      RECT MASK 1 13.464 9.875 13.524 10.105 ;
      RECT MASK 1 13.796 9.875 13.856 10.105 ;
      RECT MASK 1 14.128 9.875 14.188 10.105 ;
      RECT MASK 1 14.46 9.875 14.52 10.105 ;
      RECT MASK 1 14.792 9.875 14.852 10.105 ;
      RECT MASK 1 15.124 9.875 15.184 10.105 ;
      RECT MASK 1 15.954 9.875 16.014 10.105 ;
      RECT MASK 1 16.286 9.875 16.346 10.105 ;
      RECT MASK 1 16.618 9.875 16.678 10.105 ;
      RECT MASK 1 16.95 9.875 17.01 10.105 ;
      RECT MASK 1 17.282 9.875 17.342 10.105 ;
      RECT MASK 1 17.614 9.875 17.674 10.105 ;
      RECT MASK 1 17.946 9.875 18.006 10.105 ;
      RECT MASK 1 18.278 9.875 18.338 10.105 ;
      RECT MASK 1 18.61 9.875 18.67 10.105 ;
      RECT MASK 1 18.942 9.875 19.002 10.105 ;
      RECT MASK 1 19.274 9.875 19.334 10.105 ;
      RECT MASK 1 19.606 9.875 19.666 10.105 ;
      RECT MASK 1 19.938 9.875 19.998 10.105 ;
      RECT MASK 1 20.27 9.875 20.33 10.105 ;
      RECT MASK 1 20.602 9.875 20.662 10.105 ;
      RECT MASK 1 20.934 9.875 20.994 10.105 ;
      RECT MASK 1 21.266 9.875 21.326 10.105 ;
      RECT MASK 1 21.598 9.875 21.658 10.105 ;
      RECT MASK 1 21.93 9.875 21.99 10.105 ;
      RECT MASK 1 22.262 9.875 22.322 10.105 ;
      RECT MASK 1 22.594 9.875 22.654 10.105 ;
      RECT MASK 1 22.926 9.875 22.986 10.105 ;
      RECT MASK 1 23.258 9.875 23.318 10.105 ;
      RECT MASK 1 23.59 9.875 23.65 10.105 ;
      RECT MASK 1 23.922 9.875 23.982 10.105 ;
      RECT MASK 1 24.254 9.875 24.314 10.105 ;
      RECT MASK 1 24.586 9.875 24.646 10.105 ;
      RECT MASK 1 24.918 9.875 24.978 10.105 ;
      RECT MASK 1 25.25 9.875 25.31 10.105 ;
      RECT MASK 1 25.582 9.875 25.642 10.105 ;
      RECT MASK 1 25.914 9.875 25.974 10.105 ;
      RECT MASK 1 26.246 9.875 26.306 10.105 ;
      RECT MASK 1 26.578 9.875 26.638 10.105 ;
      RECT MASK 1 27.574 9.875 27.634 10.105 ;
      RECT MASK 1 10.664 10.255 10.724 16.81 ;
      RECT MASK 1 10.996 10.255 11.056 16.81 ;
      RECT MASK 1 11.686 10.255 11.746 10.565 ;
      RECT MASK 1 11.886 10.255 11.946 10.565 ;
      RECT MASK 1 12.086 10.255 12.146 10.565 ;
      RECT MASK 1 12.286 10.255 12.346 10.565 ;
      RECT MASK 1 12.486 10.255 12.546 10.565 ;
      RECT MASK 1 12.686 10.255 12.746 10.565 ;
      RECT MASK 1 12.886 10.255 12.946 10.565 ;
      RECT MASK 1 13.086 10.255 13.146 10.565 ;
      RECT MASK 1 13.286 10.255 13.346 10.565 ;
      RECT MASK 1 13.486 10.255 13.546 10.565 ;
      RECT MASK 1 13.686 10.255 13.746 10.565 ;
      RECT MASK 1 13.886 10.255 13.946 10.565 ;
      RECT MASK 1 14.086 10.255 14.146 10.565 ;
      RECT MASK 1 14.286 10.255 14.346 10.565 ;
      RECT MASK 1 14.486 10.255 14.546 10.565 ;
      RECT MASK 1 14.686 10.255 14.746 10.565 ;
      RECT MASK 1 14.886 10.255 14.946 10.565 ;
      RECT MASK 1 15.086 10.255 15.146 10.565 ;
      RECT MASK 1 15.286 10.255 15.346 10.565 ;
      RECT MASK 1 7.654 10.295 7.714 10.525 ;
      RECT MASK 1 8.318 10.295 8.378 12.565 ;
      RECT MASK 1 8.65 10.295 8.71 11.152 ;
      RECT MASK 1 8.982 10.295 9.042 11.152 ;
      RECT MASK 1 9.314 10.295 9.374 11.152 ;
      RECT MASK 1 9.646 10.295 9.706 10.525 ;
      RECT MASK 1 15.902 10.295 15.962 10.525 ;
      RECT MASK 1 16.102 10.295 16.162 10.525 ;
      RECT MASK 1 16.302 10.295 16.362 10.525 ;
      RECT MASK 1 16.502 10.295 16.562 10.525 ;
      RECT MASK 1 16.702 10.295 16.762 10.525 ;
      RECT MASK 1 16.902 10.295 16.962 10.525 ;
      RECT MASK 1 17.102 10.295 17.162 10.525 ;
      RECT MASK 1 17.302 10.295 17.362 10.525 ;
      RECT MASK 1 17.502 10.295 17.562 10.525 ;
      RECT MASK 1 17.702 10.295 17.762 10.525 ;
      RECT MASK 1 17.902 10.295 17.962 10.525 ;
      RECT MASK 1 18.102 10.295 18.162 10.525 ;
      RECT MASK 1 18.302 10.295 18.362 10.525 ;
      RECT MASK 1 18.502 10.295 18.562 10.525 ;
      RECT MASK 1 18.702 10.295 18.762 10.525 ;
      RECT MASK 1 18.902 10.295 18.962 10.525 ;
      RECT MASK 1 19.102 10.295 19.162 10.525 ;
      RECT MASK 1 19.302 10.295 19.362 10.525 ;
      RECT MASK 1 19.502 10.295 19.562 10.525 ;
      RECT MASK 1 19.702 10.295 19.762 10.525 ;
      RECT MASK 1 19.902 10.295 19.962 10.525 ;
      RECT MASK 1 20.102 10.295 20.162 10.525 ;
      RECT MASK 1 20.302 10.295 20.362 10.525 ;
      RECT MASK 1 20.502 10.295 20.562 10.525 ;
      RECT MASK 1 20.702 10.295 20.762 10.525 ;
      RECT MASK 1 20.902 10.295 20.962 10.525 ;
      RECT MASK 1 21.102 10.295 21.162 10.525 ;
      RECT MASK 1 21.302 10.295 21.362 10.525 ;
      RECT MASK 1 21.502 10.295 21.562 10.525 ;
      RECT MASK 1 21.702 10.295 21.762 10.525 ;
      RECT MASK 1 21.902 10.295 21.962 10.525 ;
      RECT MASK 1 22.102 10.295 22.162 10.525 ;
      RECT MASK 1 22.302 10.295 22.362 10.525 ;
      RECT MASK 1 22.502 10.295 22.562 10.525 ;
      RECT MASK 1 22.702 10.295 22.762 10.525 ;
      RECT MASK 1 22.902 10.295 22.962 10.525 ;
      RECT MASK 1 23.102 10.295 23.162 10.525 ;
      RECT MASK 1 23.302 10.295 23.362 10.525 ;
      RECT MASK 1 23.502 10.295 23.562 10.525 ;
      RECT MASK 1 23.702 10.295 23.762 10.525 ;
      RECT MASK 1 23.902 10.295 23.962 10.525 ;
      RECT MASK 1 24.102 10.295 24.162 10.525 ;
      RECT MASK 1 24.302 10.295 24.362 10.525 ;
      RECT MASK 1 24.502 10.295 24.562 10.525 ;
      RECT MASK 1 24.702 10.295 24.762 10.525 ;
      RECT MASK 1 27.846 10.295 27.906 10.525 ;
      RECT MASK 1 28.12 10.295 28.18 10.525 ;
      RECT MASK 1 28.394 10.295 28.454 10.525 ;
      RECT MASK 1 10.134 10.32 10.214 12.54 ;
      RECT MASK 1 10.83 10.375 10.89 16.81 ;
      RECT MASK 1 25.654 10.5 25.714 12.42 ;
      RECT MASK 1 25.928 10.5 25.988 12.42 ;
      RECT MASK 1 26.202 10.5 26.262 12.42 ;
      RECT MASK 1 26.476 10.5 26.536 12.42 ;
      RECT MASK 1 26.75 10.5 26.81 12.42 ;
      RECT MASK 1 27.024 10.5 27.084 12.42 ;
      RECT MASK 1 27.298 10.5 27.358 12.42 ;
      RECT MASK 1 11.769 10.693 11.829 10.941 ;
      RECT MASK 1 12.267 10.693 12.327 10.941 ;
      RECT MASK 1 12.765 10.693 12.825 10.946 ;
      RECT MASK 1 14.757 10.75 14.817 10.941 ;
      RECT MASK 1 13.097 10.752 13.157 10.946 ;
      RECT MASK 1 13.429 10.752 13.489 10.946 ;
      RECT MASK 1 13.761 10.752 13.821 10.946 ;
      RECT MASK 1 14.259 10.752 14.319 10.946 ;
      RECT MASK 1 15.255 10.752 15.315 10.946 ;
      RECT MASK 1 15.587 10.752 15.647 10.941 ;
      RECT MASK 1 15.919 10.752 15.979 10.941 ;
      RECT MASK 1 16.251 10.752 16.311 10.941 ;
      RECT MASK 1 17.247 10.752 17.307 10.946 ;
      RECT MASK 1 17.745 10.752 17.805 10.941 ;
      RECT MASK 1 18.409 10.752 18.469 10.946 ;
      RECT MASK 1 18.907 10.752 18.967 10.946 ;
      RECT MASK 1 19.239 10.752 19.299 10.946 ;
      RECT MASK 1 19.571 10.752 19.631 10.946 ;
      RECT MASK 1 20.069 10.752 20.129 10.946 ;
      RECT MASK 1 20.401 10.752 20.461 10.946 ;
      RECT MASK 1 20.899 10.752 20.959 10.946 ;
      RECT MASK 1 21.231 10.752 21.291 10.946 ;
      RECT MASK 1 21.563 10.752 21.623 10.946 ;
      RECT MASK 1 22.061 10.752 22.121 10.946 ;
      RECT MASK 1 22.393 10.752 22.453 10.946 ;
      RECT MASK 1 22.891 10.752 22.951 11.2385 ;
      RECT MASK 1 23.223 10.752 23.283 10.946 ;
      RECT MASK 1 23.555 10.752 23.615 11.2385 ;
      RECT MASK 1 24.053 10.752 24.113 11.2385 ;
      RECT MASK 1 24.453 10.752 24.513 11.2385 ;
      RECT MASK 1 24.653 10.752 24.713 11.2385 ;
      RECT MASK 1 12.101 10.958 12.161 11.782 ;
      RECT MASK 1 12.599 10.958 12.659 11.782 ;
      RECT MASK 1 15.089 10.958 15.149 11.782 ;
      RECT MASK 1 16.915 10.958 16.975 11.782 ;
      RECT MASK 1 18.077 10.958 18.137 11.782 ;
      RECT MASK 1 11.769 11.061 11.829 11.679 ;
      RECT MASK 1 12.267 11.061 12.327 11.679 ;
      RECT MASK 1 14.757 11.061 14.817 11.679 ;
      RECT MASK 1 12.765 11.066 12.825 11.674 ;
      RECT MASK 1 13.097 11.066 13.157 11.674 ;
      RECT MASK 1 13.429 11.066 13.489 11.674 ;
      RECT MASK 1 15.255 11.066 15.315 11.674 ;
      RECT MASK 1 15.587 11.066 15.647 11.674 ;
      RECT MASK 1 15.919 11.066 15.979 11.674 ;
      RECT MASK 1 16.583 11.066 16.643 11.674 ;
      RECT MASK 1 19.239 11.066 19.299 11.674 ;
      RECT MASK 1 21.231 11.066 21.291 11.674 ;
      RECT MASK 1 23.223 11.066 23.283 11.674 ;
      RECT MASK 1 11.162 11.092 11.222 12.67 ;
      RECT MASK 1 6.098 11.155 6.158 12.065 ;
      RECT MASK 1 13.761 11.217 13.821 11.648 ;
      RECT MASK 1 14.259 11.217 14.319 11.523 ;
      RECT MASK 1 16.251 11.217 16.311 11.41 ;
      RECT MASK 1 17.247 11.217 17.307 11.523 ;
      RECT MASK 1 4.082 11.275 4.142 11.585 ;
      RECT MASK 1 5.522 11.275 5.582 11.585 ;
      RECT MASK 1 6.386 11.275 6.446 11.585 ;
      RECT MASK 1 7.25 11.275 7.31 11.585 ;
      RECT MASK 1 2.93 11.281 2.99 15.575 ;
      RECT MASK 1 4.37 11.281 4.43 11.705 ;
      RECT MASK 1 5.234 11.281 5.294 11.705 ;
      RECT MASK 1 5.81 11.281 5.87 11.825 ;
      RECT MASK 1 8.65 11.285 8.71 11.579 ;
      RECT MASK 1 8.982 11.285 9.042 11.579 ;
      RECT MASK 1 9.314 11.285 9.374 11.579 ;
      RECT MASK 1 6.674 11.395 6.734 11.579 ;
      RECT MASK 1 8.65 11.708 8.71 12.565 ;
      RECT MASK 1 8.982 11.708 9.042 12.565 ;
      RECT MASK 1 9.314 11.708 9.374 12.565 ;
      RECT MASK 1 2.642 11.755 2.702 14.2855 ;
      RECT MASK 1 12.765 11.794 12.825 12.047 ;
      RECT MASK 1 13.097 11.794 13.157 11.988 ;
      RECT MASK 1 13.429 11.794 13.489 11.988 ;
      RECT MASK 1 13.761 11.794 13.821 11.988 ;
      RECT MASK 1 14.259 11.794 14.319 11.988 ;
      RECT MASK 1 15.255 11.794 15.315 11.988 ;
      RECT MASK 1 17.247 11.794 17.307 11.988 ;
      RECT MASK 1 18.409 11.794 18.469 11.988 ;
      RECT MASK 1 18.907 11.794 18.967 11.988 ;
      RECT MASK 1 19.239 11.794 19.299 11.988 ;
      RECT MASK 1 19.571 11.794 19.631 11.988 ;
      RECT MASK 1 20.069 11.794 20.129 11.988 ;
      RECT MASK 1 20.401 11.794 20.461 11.988 ;
      RECT MASK 1 20.899 11.794 20.959 11.988 ;
      RECT MASK 1 21.231 11.794 21.291 11.988 ;
      RECT MASK 1 21.563 11.794 21.623 11.988 ;
      RECT MASK 1 22.061 11.794 22.121 11.988 ;
      RECT MASK 1 22.393 11.794 22.453 11.988 ;
      RECT MASK 1 22.891 11.794 22.951 11.988 ;
      RECT MASK 1 23.223 11.794 23.283 11.988 ;
      RECT MASK 1 23.555 11.794 23.615 11.988 ;
      RECT MASK 1 24.053 11.794 24.113 11.988 ;
      RECT MASK 1 11.769 11.799 11.829 12.047 ;
      RECT MASK 1 12.267 11.799 12.327 12.047 ;
      RECT MASK 1 14.757 11.799 14.817 11.99 ;
      RECT MASK 1 15.587 11.799 15.647 11.988 ;
      RECT MASK 1 15.919 11.799 15.979 11.988 ;
      RECT MASK 1 16.251 11.799 16.311 11.988 ;
      RECT MASK 1 17.745 11.799 17.805 11.988 ;
      RECT MASK 1 4.082 11.995 4.142 14.029 ;
      RECT MASK 1 11.686 12.215 11.746 12.445 ;
      RECT MASK 1 11.886 12.215 11.946 12.445 ;
      RECT MASK 1 12.086 12.215 12.146 12.445 ;
      RECT MASK 1 12.286 12.215 12.346 12.445 ;
      RECT MASK 1 12.486 12.215 12.546 12.445 ;
      RECT MASK 1 12.686 12.215 12.746 12.445 ;
      RECT MASK 1 12.886 12.215 12.946 12.445 ;
      RECT MASK 1 13.086 12.215 13.146 12.445 ;
      RECT MASK 1 13.286 12.215 13.346 12.445 ;
      RECT MASK 1 13.486 12.215 13.546 12.445 ;
      RECT MASK 1 13.686 12.215 13.746 12.445 ;
      RECT MASK 1 13.886 12.215 13.946 12.445 ;
      RECT MASK 1 14.086 12.215 14.146 12.445 ;
      RECT MASK 1 14.286 12.215 14.346 12.445 ;
      RECT MASK 1 14.486 12.215 14.546 12.445 ;
      RECT MASK 1 14.686 12.215 14.746 12.445 ;
      RECT MASK 1 14.886 12.215 14.946 12.445 ;
      RECT MASK 1 15.086 12.215 15.146 12.445 ;
      RECT MASK 1 15.286 12.215 15.346 12.445 ;
      RECT MASK 1 15.486 12.215 15.546 12.445 ;
      RECT MASK 1 15.686 12.215 15.746 12.445 ;
      RECT MASK 1 15.886 12.215 15.946 12.445 ;
      RECT MASK 1 16.086 12.215 16.146 12.445 ;
      RECT MASK 1 16.286 12.215 16.346 12.445 ;
      RECT MASK 1 16.486 12.215 16.546 12.445 ;
      RECT MASK 1 16.686 12.215 16.746 12.445 ;
      RECT MASK 1 16.886 12.215 16.946 12.445 ;
      RECT MASK 1 17.086 12.215 17.146 12.445 ;
      RECT MASK 1 17.286 12.215 17.346 12.445 ;
      RECT MASK 1 17.486 12.215 17.546 12.445 ;
      RECT MASK 1 17.686 12.215 17.746 12.445 ;
      RECT MASK 1 17.886 12.215 17.946 12.445 ;
      RECT MASK 1 18.086 12.215 18.146 12.445 ;
      RECT MASK 1 18.286 12.215 18.346 12.445 ;
      RECT MASK 1 18.486 12.215 18.546 12.445 ;
      RECT MASK 1 18.686 12.215 18.746 12.445 ;
      RECT MASK 1 18.886 12.215 18.946 12.445 ;
      RECT MASK 1 19.086 12.215 19.146 12.445 ;
      RECT MASK 1 19.286 12.215 19.346 12.445 ;
      RECT MASK 1 19.486 12.215 19.546 12.445 ;
      RECT MASK 1 19.686 12.215 19.746 12.445 ;
      RECT MASK 1 19.886 12.215 19.946 12.445 ;
      RECT MASK 1 20.086 12.215 20.146 12.445 ;
      RECT MASK 1 20.286 12.215 20.346 12.445 ;
      RECT MASK 1 20.486 12.215 20.546 12.445 ;
      RECT MASK 1 20.686 12.215 20.746 12.445 ;
      RECT MASK 1 20.886 12.215 20.946 12.445 ;
      RECT MASK 1 21.086 12.215 21.146 12.445 ;
      RECT MASK 1 21.286 12.215 21.346 12.445 ;
      RECT MASK 1 21.486 12.215 21.546 12.445 ;
      RECT MASK 1 21.686 12.215 21.746 12.445 ;
      RECT MASK 1 21.886 12.215 21.946 12.445 ;
      RECT MASK 1 22.086 12.215 22.146 12.445 ;
      RECT MASK 1 22.286 12.215 22.346 12.445 ;
      RECT MASK 1 22.486 12.215 22.546 12.445 ;
      RECT MASK 1 22.686 12.215 22.746 12.445 ;
      RECT MASK 1 22.886 12.215 22.946 12.445 ;
      RECT MASK 1 23.086 12.215 23.146 12.445 ;
      RECT MASK 1 23.286 12.215 23.346 12.445 ;
      RECT MASK 1 23.486 12.215 23.546 12.445 ;
      RECT MASK 1 23.686 12.215 23.746 12.445 ;
      RECT MASK 1 23.886 12.215 23.946 12.445 ;
      RECT MASK 1 24.086 12.215 24.146 12.445 ;
      RECT MASK 1 24.286 12.215 24.346 12.445 ;
      RECT MASK 1 7.654 12.335 7.714 12.565 ;
      RECT MASK 1 9.646 12.335 9.706 12.565 ;
      RECT MASK 1 21.002 12.63 21.082 25.05 ;
      RECT MASK 1 21.178 12.63 21.238 12.87 ;
      RECT MASK 1 21.51 12.63 21.57 12.87 ;
      RECT MASK 1 21.842 12.63 21.902 12.87 ;
      RECT MASK 1 22.174 12.63 22.234 12.87 ;
      RECT MASK 1 22.506 12.63 22.566 12.87 ;
      RECT MASK 1 22.838 12.63 22.898 12.87 ;
      RECT MASK 1 23.17 12.63 23.23 12.87 ;
      RECT MASK 1 23.502 12.63 23.562 12.87 ;
      RECT MASK 1 23.834 12.63 23.894 12.87 ;
      RECT MASK 1 24.166 12.63 24.226 12.87 ;
      RECT MASK 1 24.498 12.63 24.558 12.87 ;
      RECT MASK 1 24.83 12.63 24.89 12.87 ;
      RECT MASK 1 25.162 12.63 25.222 12.87 ;
      RECT MASK 1 25.328 12.63 25.388 12.87 ;
      RECT MASK 1 25.494 12.63 25.554 12.87 ;
      RECT MASK 1 26.564 12.63 26.624 12.87 ;
      RECT MASK 1 26.73 12.63 26.79 12.87 ;
      RECT MASK 1 26.896 12.63 26.956 12.87 ;
      RECT MASK 1 27.228 12.63 27.288 12.87 ;
      RECT MASK 1 27.56 12.63 27.62 12.87 ;
      RECT MASK 1 27.892 12.63 27.952 12.87 ;
      RECT MASK 1 28.224 12.63 28.284 12.87 ;
      RECT MASK 1 28.556 12.63 28.616 12.87 ;
      RECT MASK 1 28.888 12.63 28.948 12.87 ;
      RECT MASK 1 29.22 12.63 29.28 12.87 ;
      RECT MASK 1 29.552 12.63 29.612 12.87 ;
      RECT MASK 1 29.884 12.63 29.944 12.87 ;
      RECT MASK 1 30.216 12.63 30.276 12.87 ;
      RECT MASK 1 30.548 12.63 30.608 12.87 ;
      RECT MASK 1 30.88 12.63 30.94 12.87 ;
      RECT MASK 1 31.212 12.63 31.272 12.87 ;
      RECT MASK 1 31.544 12.63 31.604 12.87 ;
      RECT MASK 1 0.838 12.72 0.918 15.03 ;
      RECT MASK 1 10.134 12.72 10.214 15 ;
      RECT MASK 1 7.654 12.73 7.714 12.985 ;
      RECT MASK 1 8.318 12.73 8.378 15.025 ;
      RECT MASK 1 8.65 12.73 8.71 13.612 ;
      RECT MASK 1 8.982 12.73 9.042 13.612 ;
      RECT MASK 1 9.314 12.73 9.374 13.612 ;
      RECT MASK 1 9.646 12.73 9.706 12.985 ;
      RECT MASK 1 21.842 13.05 21.902 15.74 ;
      RECT MASK 1 22.838 13.05 22.898 16.05 ;
      RECT MASK 1 24.83 13.05 24.89 15.74 ;
      RECT MASK 1 13.936 13.17 13.996 17.37 ;
      RECT MASK 1 14.434 13.17 14.494 14.068 ;
      RECT MASK 1 13.53 13.255 13.59 16.145 ;
      RECT MASK 1 17.24 13.34 17.3 13.59 ;
      RECT MASK 1 18.453 13.34 18.487 13.65 ;
      RECT MASK 1 18.653 13.34 18.687 13.65 ;
      RECT MASK 1 18.853 13.34 18.887 13.65 ;
      RECT MASK 1 19.053 13.34 19.087 13.65 ;
      RECT MASK 1 19.253 13.34 19.287 13.65 ;
      RECT MASK 1 22.174 13.35 22.234 15.44 ;
      RECT MASK 1 24.166 13.35 24.226 19.5 ;
      RECT MASK 1 24.498 13.35 24.558 15.44 ;
      RECT MASK 1 21.51 13.45 21.57 16.7 ;
      RECT MASK 1 18.114 13.5 18.174 14.174 ;
      RECT MASK 1 19.666 13.5 19.726 14.174 ;
      RECT MASK 1 23.668 13.55 23.728 23.463 ;
      RECT MASK 1 30.9865 13.63 31.0865 18.5735 ;
      RECT MASK 1 3.218 13.751 3.278 14.405 ;
      RECT MASK 1 5.234 13.751 5.294 14.405 ;
      RECT MASK 1 6.386 13.751 6.446 14.405 ;
      RECT MASK 1 6.962 13.751 7.022 14.405 ;
      RECT MASK 1 7.2445 13.751 7.3045 14.405 ;
      RECT MASK 1 8.65 13.751 8.71 14.029 ;
      RECT MASK 1 8.982 13.751 9.042 14.029 ;
      RECT MASK 1 9.314 13.751 9.374 14.029 ;
      RECT MASK 1 16.242 13.834 16.302 14.5815 ;
      RECT MASK 1 12.534 13.838 12.594 15.022 ;
      RECT MASK 1 12.866 13.838 12.926 15.022 ;
      RECT MASK 1 14.102 13.838 14.162 14.47 ;
      RECT MASK 1 6.674 13.849 6.734 14.029 ;
      RECT MASK 1 18.44 13.96 18.5 14.845 ;
      RECT MASK 1 18.64 13.96 18.7 14.845 ;
      RECT MASK 1 15.172 14.03 15.232 14.825 ;
      RECT MASK 1 16.74 14.15 16.8 14.369 ;
      RECT MASK 1 17.546 14.155 17.606 14.8595 ;
      RECT MASK 1 8.65 14.168 8.71 15.025 ;
      RECT MASK 1 8.982 14.168 9.042 15.025 ;
      RECT MASK 1 9.314 14.168 9.374 15.025 ;
      RECT MASK 1 16.9005 14.39 16.9605 14.604 ;
      RECT MASK 1 17.239 14.39 17.299 14.604 ;
      RECT MASK 1 13.198 14.515 13.258 17.765 ;
      RECT MASK 1 16.242 14.6195 16.302 15.0255 ;
      RECT MASK 1 18.114 14.72 18.174 15.82 ;
      RECT MASK 1 19.666 14.72 19.726 15.82 ;
      RECT MASK 1 18.954 14.725 19.014 15.09 ;
      RECT MASK 1 19.26 14.725 19.32 15.815 ;
      RECT MASK 1 14.102 14.736 14.162 15.022 ;
      RECT MASK 1 14.434 14.736 14.494 15.022 ;
      RECT MASK 1 17.239 14.75 17.299 15.022 ;
      RECT MASK 1 17.806 14.792 17.866 15.748 ;
      RECT MASK 1 7.986 14.795 8.046 15.025 ;
      RECT MASK 1 9.646 14.795 9.706 15.025 ;
      RECT MASK 1 18.453 15.21 18.487 15.33 ;
      RECT MASK 1 18.653 15.21 18.687 15.33 ;
      RECT MASK 1 18.853 15.21 18.887 15.33 ;
      RECT MASK 1 19.053 15.21 19.087 15.33 ;
      RECT MASK 1 2.088 15.24 2.268 20.25 ;
      RECT MASK 1 0.852 15.33 0.892 16.8 ;
      RECT MASK 1 1.516 15.33 1.556 16.8 ;
      RECT MASK 1 2.48 15.351 2.54 15.609 ;
      RECT MASK 1 2.646 15.351 2.706 15.609 ;
      RECT MASK 1 3.144 15.351 3.204 15.609 ;
      RECT MASK 1 3.31 15.351 3.37 15.609 ;
      RECT MASK 1 3.476 15.351 3.536 15.609 ;
      RECT MASK 1 3.642 15.351 3.702 15.609 ;
      RECT MASK 1 3.808 15.351 3.868 15.609 ;
      RECT MASK 1 3.974 15.351 4.034 15.609 ;
      RECT MASK 1 4.14 15.351 4.2 15.609 ;
      RECT MASK 1 4.306 15.351 4.366 15.609 ;
      RECT MASK 1 4.472 15.351 4.532 15.609 ;
      RECT MASK 1 4.638 15.351 4.698 15.609 ;
      RECT MASK 1 4.804 15.351 4.864 15.609 ;
      RECT MASK 1 4.97 15.351 5.03 15.609 ;
      RECT MASK 1 5.136 15.351 5.196 15.609 ;
      RECT MASK 1 5.302 15.351 5.362 15.609 ;
      RECT MASK 1 5.468 15.351 5.528 15.609 ;
      RECT MASK 1 5.634 15.351 5.694 15.609 ;
      RECT MASK 1 5.8 15.351 5.86 15.609 ;
      RECT MASK 1 5.966 15.351 6.026 15.609 ;
      RECT MASK 1 6.132 15.351 6.192 15.609 ;
      RECT MASK 1 6.298 15.351 6.358 15.609 ;
      RECT MASK 1 6.464 15.351 6.524 15.609 ;
      RECT MASK 1 6.63 15.351 6.69 15.609 ;
      RECT MASK 1 6.796 15.351 6.856 15.609 ;
      RECT MASK 1 6.962 15.351 7.022 15.609 ;
      RECT MASK 1 7.128 15.351 7.188 15.609 ;
      RECT MASK 1 7.294 15.351 7.354 15.609 ;
      RECT MASK 1 7.46 15.351 7.52 15.609 ;
      RECT MASK 1 7.626 15.351 7.686 15.609 ;
      RECT MASK 1 7.792 15.351 7.852 15.609 ;
      RECT MASK 1 7.958 15.351 8.018 15.609 ;
      RECT MASK 1 8.124 15.351 8.184 15.609 ;
      RECT MASK 1 8.29 15.351 8.35 15.609 ;
      RECT MASK 1 8.456 15.351 8.516 15.609 ;
      RECT MASK 1 8.622 15.351 8.682 15.609 ;
      RECT MASK 1 8.788 15.351 8.848 15.609 ;
      RECT MASK 1 8.954 15.351 9.014 15.609 ;
      RECT MASK 1 9.12 15.351 9.18 15.609 ;
      RECT MASK 1 9.286 15.351 9.346 15.609 ;
      RECT MASK 1 9.452 15.351 9.512 15.609 ;
      RECT MASK 1 9.618 15.351 9.678 15.609 ;
      RECT MASK 1 9.784 15.351 9.844 15.609 ;
      RECT MASK 1 9.95 15.351 10.01 15.609 ;
      RECT MASK 1 10.116 15.351 10.176 15.609 ;
      RECT MASK 1 10.282 15.351 10.342 15.609 ;
      RECT MASK 1 18.954 15.45 19.014 15.815 ;
      RECT MASK 1 1.295 15.481 1.335 17.875 ;
      RECT MASK 1 16.242 15.5145 16.302 15.9205 ;
      RECT MASK 1 12.534 15.518 12.594 16.702 ;
      RECT MASK 1 12.866 15.518 12.926 16.702 ;
      RECT MASK 1 14.102 15.518 14.162 15.804 ;
      RECT MASK 1 14.434 15.518 14.494 15.804 ;
      RECT MASK 1 17.239 15.518 17.299 15.79 ;
      RECT MASK 1 17.546 15.6805 17.606 16.385 ;
      RECT MASK 1 18.44 15.695 18.5 16.58 ;
      RECT MASK 1 18.64 15.695 18.7 16.58 ;
      RECT MASK 1 15.172 15.715 15.232 16.51 ;
      RECT MASK 1 1.073 15.725 1.113 22.555 ;
      RECT MASK 1 2.718 15.75 2.778 20.37 ;
      RECT MASK 1 2.992 15.75 3.052 20.37 ;
      RECT MASK 1 3.266 15.75 3.326 20.37 ;
      RECT MASK 1 3.54 15.75 3.6 20.37 ;
      RECT MASK 1 3.814 15.75 3.874 20.37 ;
      RECT MASK 1 4.088 15.75 4.148 20.37 ;
      RECT MASK 1 4.362 15.75 4.422 18.78 ;
      RECT MASK 1 4.636 15.75 4.696 18.78 ;
      RECT MASK 1 4.91 15.75 4.97 18.78 ;
      RECT MASK 1 5.184 15.75 5.244 18.78 ;
      RECT MASK 1 5.458 15.75 5.518 18.78 ;
      RECT MASK 1 5.732 15.75 5.792 18.78 ;
      RECT MASK 1 6.006 15.75 6.066 18.78 ;
      RECT MASK 1 6.28 15.75 6.34 17.19 ;
      RECT MASK 1 6.554 15.75 6.614 17.19 ;
      RECT MASK 1 6.828 15.75 6.888 17.19 ;
      RECT MASK 1 7.102 15.75 7.162 17.19 ;
      RECT MASK 1 7.376 15.75 7.436 17.19 ;
      RECT MASK 1 7.65 15.75 7.71 17.19 ;
      RECT MASK 1 7.924 15.75 7.984 17.19 ;
      RECT MASK 1 8.198 15.75 8.258 17.19 ;
      RECT MASK 1 8.472 15.75 8.532 17.19 ;
      RECT MASK 1 8.746 15.75 8.806 17.19 ;
      RECT MASK 1 9.02 15.75 9.08 17.19 ;
      RECT MASK 1 9.294 15.75 9.354 17.19 ;
      RECT MASK 1 9.568 15.75 9.628 17.19 ;
      RECT MASK 1 9.842 15.75 9.902 17.19 ;
      RECT MASK 1 10.116 15.75 10.176 17.19 ;
      RECT MASK 1 10.39 15.75 10.45 17.245 ;
      RECT MASK 1 23.502 15.87 23.562 16.15 ;
      RECT MASK 1 23.834 15.87 23.894 16.15 ;
      RECT MASK 1 24.498 15.87 24.558 16.15 ;
      RECT MASK 1 24.83 15.87 24.89 16.15 ;
      RECT MASK 1 22.506 15.925 22.566 16.45 ;
      RECT MASK 1 16.9005 15.936 16.9605 16.15 ;
      RECT MASK 1 17.239 15.936 17.299 16.15 ;
      RECT MASK 1 16.242 15.9585 16.302 16.706 ;
      RECT MASK 1 14.102 16.07 14.162 16.702 ;
      RECT MASK 1 21.842 16.17 21.902 16.9 ;
      RECT MASK 1 22.174 16.17 22.234 16.9 ;
      RECT MASK 1 16.74 16.171 16.8 16.39 ;
      RECT MASK 1 18.114 16.366 18.174 17.04 ;
      RECT MASK 1 19.666 16.366 19.726 17.04 ;
      RECT MASK 1 22.838 16.37 22.898 17.1 ;
      RECT MASK 1 20.686 16.405 20.746 21.8485 ;
      RECT MASK 1 14.434 16.472 14.494 17.37 ;
      RECT MASK 1 22.506 16.62 22.566 17 ;
      RECT MASK 1 18.453 16.89 18.487 17.2 ;
      RECT MASK 1 18.653 16.89 18.687 17.2 ;
      RECT MASK 1 18.853 16.89 18.887 17.2 ;
      RECT MASK 1 19.053 16.89 19.087 17.2 ;
      RECT MASK 1 19.253 16.89 19.287 17.2 ;
      RECT MASK 1 23.502 16.92 23.562 17.61 ;
      RECT MASK 1 23.834 16.92 23.894 17.61 ;
      RECT MASK 1 24.498 16.92 24.558 17.61 ;
      RECT MASK 1 24.83 16.92 24.89 17.61 ;
      RECT MASK 1 17.24 16.95 17.3 17.2 ;
      RECT MASK 1 0.852 16.978 0.892 19.35 ;
      RECT MASK 1 1.516 16.978 1.556 19.35 ;
      RECT MASK 1 30.4885 16.99 30.5885 20.21 ;
      RECT MASK 1 23.17 17.02 23.23 20.36 ;
      RECT MASK 1 6.28 17.34 6.34 18.815 ;
      RECT MASK 1 21.842 17.37 21.902 18.275 ;
      RECT MASK 1 22.174 17.37 22.234 18.275 ;
      RECT MASK 1 22.506 17.37 22.566 18.275 ;
      RECT MASK 1 22.838 17.37 22.898 18.275 ;
      RECT MASK 1 23.502 17.79 23.562 18.275 ;
      RECT MASK 1 1.295 18.005 1.335 22.555 ;
      RECT MASK 1 7.367 18.017 7.427 18.803 ;
      RECT MASK 1 7.865 18.017 7.925 18.803 ;
      RECT MASK 1 8.363 18.017 8.423 18.803 ;
      RECT MASK 1 9.027 18.017 9.087 18.808 ;
      RECT MASK 1 9.359 18.017 9.419 18.947 ;
      RECT MASK 1 9.608 18.017 9.668 18.947 ;
      RECT MASK 1 9.774 18.017 9.834 18.947 ;
      RECT MASK 1 9.94 18.017 10 18.723 ;
      RECT MASK 1 10.106 18.017 10.166 18.947 ;
      RECT MASK 1 10.272 18.017 10.332 18.947 ;
      RECT MASK 1 10.438 18.017 10.498 18.947 ;
      RECT MASK 1 10.604 18.017 10.664 18.641 ;
      RECT MASK 1 10.77 18.017 10.83 18.947 ;
      RECT MASK 1 10.936 18.017 10.996 18.947 ;
      RECT MASK 1 11.102 18.017 11.162 18.947 ;
      RECT MASK 1 11.268 18.017 11.328 18.723 ;
      RECT MASK 1 11.434 18.017 11.494 18.947 ;
      RECT MASK 1 11.6 18.017 11.66 18.947 ;
      RECT MASK 1 11.766 18.017 11.826 18.947 ;
      RECT MASK 1 11.932 18.017 11.992 18.641 ;
      RECT MASK 1 12.098 18.017 12.158 18.947 ;
      RECT MASK 1 12.264 18.017 12.324 18.947 ;
      RECT MASK 1 12.43 18.017 12.49 18.947 ;
      RECT MASK 1 12.596 18.017 12.656 18.723 ;
      RECT MASK 1 12.762 18.017 12.822 18.947 ;
      RECT MASK 1 12.928 18.017 12.988 18.947 ;
      RECT MASK 1 13.094 18.017 13.154 18.947 ;
      RECT MASK 1 13.26 18.017 13.32 18.641 ;
      RECT MASK 1 13.426 18.017 13.486 18.947 ;
      RECT MASK 1 13.592 18.017 13.652 18.947 ;
      RECT MASK 1 13.758 18.017 13.818 18.947 ;
      RECT MASK 1 13.924 18.017 13.984 18.723 ;
      RECT MASK 1 14.09 18.017 14.15 18.947 ;
      RECT MASK 1 14.256 18.017 14.316 18.947 ;
      RECT MASK 1 14.422 18.017 14.482 18.947 ;
      RECT MASK 1 14.588 18.017 14.648 18.641 ;
      RECT MASK 1 14.754 18.017 14.814 18.947 ;
      RECT MASK 1 14.92 18.017 14.98 18.947 ;
      RECT MASK 1 15.086 18.017 15.146 18.947 ;
      RECT MASK 1 15.252 18.017 15.312 18.723 ;
      RECT MASK 1 15.418 18.017 15.478 18.947 ;
      RECT MASK 1 15.584 18.017 15.644 18.947 ;
      RECT MASK 1 15.75 18.017 15.81 18.947 ;
      RECT MASK 1 15.916 18.017 15.976 18.641 ;
      RECT MASK 1 16.082 18.017 16.142 18.947 ;
      RECT MASK 1 16.248 18.017 16.308 18.947 ;
      RECT MASK 1 16.414 18.017 16.474 18.947 ;
      RECT MASK 1 16.58 18.017 16.64 18.723 ;
      RECT MASK 1 16.746 18.017 16.806 18.947 ;
      RECT MASK 1 16.912 18.017 16.972 18.947 ;
      RECT MASK 1 17.078 18.017 17.138 18.947 ;
      RECT MASK 1 17.244 18.017 17.304 18.641 ;
      RECT MASK 1 17.41 18.017 17.47 18.947 ;
      RECT MASK 1 17.576 18.017 17.636 18.947 ;
      RECT MASK 1 17.742 18.017 17.802 18.947 ;
      RECT MASK 1 17.908 18.017 17.968 18.723 ;
      RECT MASK 1 18.074 18.017 18.134 18.947 ;
      RECT MASK 1 18.24 18.017 18.3 18.947 ;
      RECT MASK 1 18.406 18.017 18.466 18.947 ;
      RECT MASK 1 18.572 18.017 18.632 18.641 ;
      RECT MASK 1 18.738 18.017 18.798 18.947 ;
      RECT MASK 1 18.904 18.017 18.964 18.947 ;
      RECT MASK 1 19.07 18.017 19.13 18.947 ;
      RECT MASK 1 19.236 18.017 19.296 18.723 ;
      RECT MASK 1 19.402 18.017 19.462 18.947 ;
      RECT MASK 1 19.568 18.017 19.628 18.947 ;
      RECT MASK 1 19.734 18.017 19.794 18.947 ;
      RECT MASK 1 19.9 18.017 19.96 18.641 ;
      RECT MASK 1 20.066 18.017 20.126 18.947 ;
      RECT MASK 1 23.502 18.67 23.562 19.12 ;
      RECT MASK 1 7.699 18.728 7.759 19.552 ;
      RECT MASK 1 8.197 18.728 8.257 19.552 ;
      RECT MASK 1 8.695 18.728 8.755 19.552 ;
      RECT MASK 1 10.604 18.803 10.664 19.477 ;
      RECT MASK 1 11.932 18.803 11.992 19.477 ;
      RECT MASK 1 13.26 18.803 13.32 19.477 ;
      RECT MASK 1 14.588 18.803 14.648 19.477 ;
      RECT MASK 1 15.916 18.803 15.976 19.477 ;
      RECT MASK 1 17.244 18.803 17.304 19.477 ;
      RECT MASK 1 18.572 18.803 18.632 19.477 ;
      RECT MASK 1 19.9 18.803 19.96 19.477 ;
      RECT MASK 1 4.362 18.93 4.422 20.37 ;
      RECT MASK 1 7.367 18.9865 7.427 19.293 ;
      RECT MASK 1 7.865 18.9865 7.925 19.293 ;
      RECT MASK 1 8.363 18.9865 8.423 19.293 ;
      RECT MASK 1 9.027 18.987 9.087 19.552 ;
      RECT MASK 1 5.502 19.015 5.542 19.445 ;
      RECT MASK 1 5.702 19.015 5.742 19.46 ;
      RECT MASK 1 5.902 19.015 5.942 19.445 ;
      RECT MASK 1 6.102 19.015 6.142 19.445 ;
      RECT MASK 1 6.302 19.015 6.342 19.445 ;
      RECT MASK 1 20.274 19.357 20.334 21.002 ;
      RECT MASK 1 9.359 19.367 9.419 20.261 ;
      RECT MASK 1 9.608 19.367 9.668 20.237 ;
      RECT MASK 1 9.774 19.367 9.834 20.237 ;
      RECT MASK 1 10.106 19.367 10.166 20.237 ;
      RECT MASK 1 10.272 19.367 10.332 20.237 ;
      RECT MASK 1 10.438 19.367 10.498 20.237 ;
      RECT MASK 1 10.77 19.367 10.83 20.237 ;
      RECT MASK 1 10.936 19.367 10.996 20.237 ;
      RECT MASK 1 11.102 19.367 11.162 20.237 ;
      RECT MASK 1 11.434 19.367 11.494 20.237 ;
      RECT MASK 1 11.6 19.367 11.66 20.237 ;
      RECT MASK 1 11.766 19.367 11.826 20.237 ;
      RECT MASK 1 12.098 19.367 12.158 20.237 ;
      RECT MASK 1 12.264 19.367 12.324 20.237 ;
      RECT MASK 1 12.43 19.367 12.49 20.237 ;
      RECT MASK 1 12.762 19.367 12.822 20.237 ;
      RECT MASK 1 12.928 19.367 12.988 20.237 ;
      RECT MASK 1 13.094 19.367 13.154 20.237 ;
      RECT MASK 1 13.426 19.367 13.486 20.237 ;
      RECT MASK 1 13.592 19.367 13.652 20.237 ;
      RECT MASK 1 13.758 19.367 13.818 20.237 ;
      RECT MASK 1 14.09 19.367 14.15 20.237 ;
      RECT MASK 1 14.256 19.367 14.316 20.237 ;
      RECT MASK 1 14.422 19.367 14.482 20.237 ;
      RECT MASK 1 14.754 19.367 14.814 20.237 ;
      RECT MASK 1 14.92 19.367 14.98 20.237 ;
      RECT MASK 1 15.086 19.367 15.146 20.237 ;
      RECT MASK 1 15.418 19.367 15.478 20.237 ;
      RECT MASK 1 15.584 19.367 15.644 20.237 ;
      RECT MASK 1 15.75 19.367 15.81 20.237 ;
      RECT MASK 1 16.082 19.367 16.142 20.237 ;
      RECT MASK 1 16.248 19.367 16.308 20.237 ;
      RECT MASK 1 16.414 19.367 16.474 20.237 ;
      RECT MASK 1 16.746 19.367 16.806 20.237 ;
      RECT MASK 1 16.912 19.367 16.972 20.237 ;
      RECT MASK 1 17.078 19.367 17.138 20.237 ;
      RECT MASK 1 17.41 19.367 17.47 20.237 ;
      RECT MASK 1 17.576 19.367 17.636 20.237 ;
      RECT MASK 1 17.742 19.367 17.802 20.237 ;
      RECT MASK 1 18.074 19.367 18.134 20.237 ;
      RECT MASK 1 18.24 19.367 18.3 20.237 ;
      RECT MASK 1 18.406 19.367 18.466 20.147 ;
      RECT MASK 1 18.738 19.367 18.798 20.237 ;
      RECT MASK 1 18.904 19.367 18.964 20.237 ;
      RECT MASK 1 19.07 19.367 19.13 20.237 ;
      RECT MASK 1 19.402 19.367 19.462 20.237 ;
      RECT MASK 1 19.568 19.367 19.628 20.237 ;
      RECT MASK 1 19.734 19.367 19.794 20.237 ;
      RECT MASK 1 20.066 19.367 20.126 20.237 ;
      RECT MASK 1 7.367 19.477 7.427 20.261 ;
      RECT MASK 1 7.865 19.477 7.925 20.261 ;
      RECT MASK 1 8.363 19.477 8.423 20.261 ;
      RECT MASK 1 23.834 19.52 23.894 19.8 ;
      RECT MASK 1 0.852 19.53 0.892 24.145 ;
      RECT MASK 1 1.516 19.53 1.556 24.145 ;
      RECT MASK 1 9.94 19.562 10 20.237 ;
      RECT MASK 1 11.268 19.562 11.328 20.237 ;
      RECT MASK 1 12.596 19.562 12.656 20.237 ;
      RECT MASK 1 13.924 19.562 13.984 20.237 ;
      RECT MASK 1 15.252 19.562 15.312 20.237 ;
      RECT MASK 1 16.58 19.562 16.64 20.237 ;
      RECT MASK 1 17.908 19.562 17.968 20.237 ;
      RECT MASK 1 19.236 19.562 19.296 20.237 ;
      RECT MASK 1 10.604 19.639 10.664 20.237 ;
      RECT MASK 1 11.932 19.639 11.992 20.237 ;
      RECT MASK 1 13.26 19.639 13.32 20.237 ;
      RECT MASK 1 14.588 19.639 14.648 20.237 ;
      RECT MASK 1 15.916 19.639 15.976 20.237 ;
      RECT MASK 1 17.244 19.639 17.304 20.237 ;
      RECT MASK 1 18.572 19.639 18.632 20.147 ;
      RECT MASK 1 19.9 19.639 19.96 20.237 ;
      RECT MASK 1 5.702 19.72 5.742 20.1685 ;
      RECT MASK 1 5.502 19.735 5.542 20.1685 ;
      RECT MASK 1 5.902 19.735 5.942 20.1685 ;
      RECT MASK 1 6.102 19.735 6.142 20.1685 ;
      RECT MASK 1 6.302 19.735 6.342 20.1685 ;
      RECT MASK 1 23.834 19.98 23.894 20.97 ;
      RECT MASK 1 21.842 20.125 21.902 20.97 ;
      RECT MASK 1 22.174 20.125 22.234 20.97 ;
      RECT MASK 1 22.506 20.125 22.566 20.97 ;
      RECT MASK 1 22.838 20.125 22.898 20.97 ;
      RECT MASK 1 23.502 20.125 23.562 20.97 ;
      RECT MASK 1 14.547 20.381 14.607 21.002 ;
      RECT MASK 1 14.879 20.381 14.939 20.752 ;
      RECT MASK 1 15.377 20.381 15.437 21.002 ;
      RECT MASK 1 16.041 20.381 16.101 21.002 ;
      RECT MASK 1 16.539 20.381 16.599 20.636 ;
      RECT MASK 1 17.037 20.381 17.097 21.002 ;
      RECT MASK 1 17.452 20.381 17.512 21.002 ;
      RECT MASK 1 17.618 20.381 17.678 21.002 ;
      RECT MASK 1 17.784 20.381 17.844 20.636 ;
      RECT MASK 1 17.95 20.381 18.01 21.002 ;
      RECT MASK 1 18.116 20.381 18.176 21.002 ;
      RECT MASK 1 18.282 20.381 18.342 21.002 ;
      RECT MASK 1 18.614 20.381 18.674 21.002 ;
      RECT MASK 1 18.78 20.381 18.84 21.002 ;
      RECT MASK 1 18.946 20.381 19.006 21.002 ;
      RECT MASK 1 19.112 20.381 19.172 20.636 ;
      RECT MASK 1 19.278 20.381 19.338 21.002 ;
      RECT MASK 1 19.444 20.381 19.504 21.002 ;
      RECT MASK 1 19.61 20.381 19.67 21.002 ;
      RECT MASK 1 19.942 20.381 20.002 21.002 ;
      RECT MASK 1 20.108 20.381 20.168 21.002 ;
      RECT MASK 1 3.498 20.49 3.558 24.111 ;
      RECT MASK 1 15.709 20.648 15.769 21.472 ;
      RECT MASK 1 11.763 20.7 11.823 21.51 ;
      RECT MASK 1 12.095 20.7 12.155 21.51 ;
      RECT MASK 1 12.676 20.7 12.736 21.51 ;
      RECT MASK 1 13.008 20.7 13.068 21.51 ;
      RECT MASK 1 13.34 20.7 13.4 21.51 ;
      RECT MASK 1 23.17 20.73 23.23 20.97 ;
      RECT MASK 1 24.166 20.73 24.226 20.97 ;
      RECT MASK 1 24.498 20.73 24.558 20.97 ;
      RECT MASK 1 24.83 20.73 24.89 20.97 ;
      RECT MASK 1 16.539 20.756 16.599 21.364 ;
      RECT MASK 1 14.879 20.907 14.939 21.305 ;
      RECT MASK 1 4.27 20.915 4.33 22.558 ;
      RECT MASK 1 5.496 20.915 5.556 22.558 ;
      RECT MASK 1 2.403 20.94 2.437 21.15 ;
      RECT MASK 1 2.631 20.94 2.665 21.7 ;
      RECT MASK 1 2.859 20.94 2.893 21.15 ;
      RECT MASK 1 3.074 20.94 3.134 21.56 ;
      RECT MASK 1 14.132 21.2225 14.192 22.3375 ;
      RECT MASK 1 20.44 21.2225 20.5 22.3375 ;
      RECT MASK 1 6.056 21.235 6.116 21.508 ;
      RECT MASK 1 6.388 21.235 6.448 21.508 ;
      RECT MASK 1 6.72 21.235 6.78 21.508 ;
      RECT MASK 1 7.052 21.235 7.112 21.508 ;
      RECT MASK 1 7.384 21.235 7.444 21.508 ;
      RECT MASK 1 7.716 21.235 7.776 21.508 ;
      RECT MASK 1 8.048 21.235 8.108 21.508 ;
      RECT MASK 1 8.38 21.235 8.44 21.508 ;
      RECT MASK 1 8.712 21.235 8.772 21.508 ;
      RECT MASK 1 9.044 21.235 9.104 21.508 ;
      RECT MASK 1 9.376 21.235 9.436 21.508 ;
      RECT MASK 1 10.103 21.278 10.163 22.019 ;
      RECT MASK 1 10.767 21.278 10.827 22.015 ;
      RECT MASK 1 11.099 21.278 11.159 21.785 ;
      RECT MASK 1 11.431 21.278 11.491 22.462 ;
      RECT MASK 1 5.145 21.289 5.205 22.286 ;
      RECT MASK 1 12.344 21.475 12.404 22.505 ;
      RECT MASK 1 14.335 21.484 14.395 22.309 ;
      RECT MASK 1 14.713 21.484 14.773 22.309 ;
      RECT MASK 1 14.879 21.484 14.939 21.678 ;
      RECT MASK 1 16.041 21.484 16.101 22.309 ;
      RECT MASK 1 16.539 21.484 16.599 22.076 ;
      RECT MASK 1 17.037 21.484 17.097 22.309 ;
      RECT MASK 1 17.452 21.484 17.512 22.265 ;
      RECT MASK 1 17.618 21.484 17.678 22.265 ;
      RECT MASK 1 17.784 21.484 17.844 22.076 ;
      RECT MASK 1 17.95 21.484 18.01 22.265 ;
      RECT MASK 1 18.116 21.484 18.176 22.265 ;
      RECT MASK 1 18.282 21.484 18.342 22.265 ;
      RECT MASK 1 18.614 21.484 18.674 22.265 ;
      RECT MASK 1 18.78 21.484 18.84 22.265 ;
      RECT MASK 1 18.946 21.484 19.006 22.265 ;
      RECT MASK 1 19.112 21.484 19.172 22.081 ;
      RECT MASK 1 19.278 21.484 19.338 22.265 ;
      RECT MASK 1 19.444 21.484 19.504 22.265 ;
      RECT MASK 1 19.61 21.484 19.67 22.265 ;
      RECT MASK 1 19.942 21.484 20.002 22.265 ;
      RECT MASK 1 20.108 21.484 20.168 22.309 ;
      RECT MASK 1 20.274 21.484 20.334 22.309 ;
      RECT MASK 1 15.377 21.489 15.437 22.071 ;
      RECT MASK 1 15.045 21.592 15.105 21.968 ;
      RECT MASK 1 15.709 21.592 15.769 21.968 ;
      RECT MASK 1 18.448 21.592 18.508 21.968 ;
      RECT MASK 1 19.776 21.592 19.836 21.967 ;
      RECT MASK 1 10.435 21.628 10.495 21.946 ;
      RECT MASK 1 13.34 21.63 13.4 22.15 ;
      RECT MASK 1 11.763 21.715 11.823 22.112 ;
      RECT MASK 1 2.161 21.725 2.221 21.905 ;
      RECT MASK 1 9.771 21.734 9.831 22.51 ;
      RECT MASK 1 13.838 21.74 13.898 24.005 ;
      RECT MASK 1 22.53 21.8915 22.59 22.82 ;
      RECT MASK 1 22.73 21.8915 22.79 22.82 ;
      RECT MASK 1 22.93 21.8915 22.99 22.82 ;
      RECT MASK 1 23.93 21.898 23.99 22.82 ;
      RECT MASK 1 24.13 21.898 24.19 22.82 ;
      RECT MASK 1 12.012 21.93 12.072 22.112 ;
      RECT MASK 1 11.099 21.955 11.159 22.462 ;
      RECT MASK 1 2.161 22.075 2.221 22.8 ;
      RECT MASK 1 3.074 22.075 3.134 22.8 ;
      RECT MASK 1 15.045 22.088 15.105 22.912 ;
      RECT MASK 1 15.709 22.088 15.769 22.912 ;
      RECT MASK 1 2.631 22.16 2.665 22.8 ;
      RECT MASK 1 6.056 22.195 6.116 22.462 ;
      RECT MASK 1 10.435 22.195 10.495 23.645 ;
      RECT MASK 1 10.767 22.195 10.827 23.645 ;
      RECT MASK 1 12.676 22.195 12.736 23.645 ;
      RECT MASK 1 13.008 22.195 13.068 23.645 ;
      RECT MASK 1 16.539 22.196 16.599 22.804 ;
      RECT MASK 1 6.388 22.232 6.448 23.608 ;
      RECT MASK 1 6.72 22.232 6.78 22.462 ;
      RECT MASK 1 7.052 22.232 7.112 23.608 ;
      RECT MASK 1 7.384 22.232 7.444 23.608 ;
      RECT MASK 1 7.716 22.232 7.776 23.608 ;
      RECT MASK 1 8.048 22.232 8.108 23.608 ;
      RECT MASK 1 8.38 22.232 8.44 23.608 ;
      RECT MASK 1 8.712 22.232 8.772 23.608 ;
      RECT MASK 1 9.044 22.232 9.104 23.608 ;
      RECT MASK 1 9.376 22.232 9.436 23.608 ;
      RECT MASK 1 10.103 22.232 10.163 22.505 ;
      RECT MASK 1 11.763 22.232 11.823 23.608 ;
      RECT MASK 1 12.095 22.232 12.155 23.608 ;
      RECT MASK 1 13.34 22.27 13.4 23.57 ;
      RECT MASK 1 4.813 22.427 4.873 22.835 ;
      RECT MASK 1 2.403 22.59 2.437 22.8 ;
      RECT MASK 1 2.859 22.59 2.893 22.8 ;
      RECT MASK 1 14.335 22.685 14.395 23.516 ;
      RECT MASK 1 14.713 22.685 14.773 23.516 ;
      RECT MASK 1 15.377 22.685 15.437 23.179 ;
      RECT MASK 1 16.041 22.685 16.101 23.516 ;
      RECT MASK 1 17.037 22.685 17.097 23.516 ;
      RECT MASK 1 17.452 22.685 17.512 23.179 ;
      RECT MASK 1 17.618 22.685 17.678 23.179 ;
      RECT MASK 1 17.95 22.685 18.01 23.179 ;
      RECT MASK 1 18.116 22.685 18.176 23.179 ;
      RECT MASK 1 18.282 22.685 18.342 23.179 ;
      RECT MASK 1 18.614 22.685 18.674 23.179 ;
      RECT MASK 1 18.78 22.685 18.84 23.179 ;
      RECT MASK 1 18.946 22.685 19.006 23.179 ;
      RECT MASK 1 19.278 22.685 19.338 23.179 ;
      RECT MASK 1 19.444 22.685 19.504 23.179 ;
      RECT MASK 1 19.61 22.685 19.67 23.179 ;
      RECT MASK 1 19.942 22.685 20.002 23.408 ;
      RECT MASK 1 20.274 22.685 20.334 23.516 ;
      RECT MASK 1 16.539 22.924 16.599 23.516 ;
      RECT MASK 1 17.784 22.924 17.844 23.179 ;
      RECT MASK 1 19.112 22.924 19.172 23.179 ;
      RECT MASK 1 1.295 22.934 1.335 23.643 ;
      RECT MASK 1 22.53 23 22.59 23.8845 ;
      RECT MASK 1 22.73 23 22.79 23.8845 ;
      RECT MASK 1 22.93 23 22.99 23.8845 ;
      RECT MASK 1 23.93 23 23.99 23.8815 ;
      RECT MASK 1 24.13 23 24.19 23.8815 ;
      RECT MASK 1 4.813 23.005 4.873 23.413 ;
      RECT MASK 1 15.709 23.033 15.769 23.516 ;
      RECT MASK 1 2.161 23.04 2.221 23.705 ;
      RECT MASK 1 2.403 23.04 2.437 23.25 ;
      RECT MASK 1 2.631 23.04 2.665 23.705 ;
      RECT MASK 1 2.859 23.04 2.893 23.25 ;
      RECT MASK 1 3.074 23.04 3.134 23.705 ;
      RECT MASK 1 15.211 23.261 15.271 23.516 ;
      RECT MASK 1 4.27 23.282 4.33 24.925 ;
      RECT MASK 1 5.496 23.282 5.556 24.925 ;
      RECT MASK 1 17.369 23.322 17.429 23.516 ;
      RECT MASK 1 17.867 23.322 17.927 23.516 ;
      RECT MASK 1 18.365 23.322 18.425 23.516 ;
      RECT MASK 1 18.697 23.322 18.757 23.516 ;
      RECT MASK 1 19.195 23.322 19.255 23.516 ;
      RECT MASK 1 19.693 23.322 19.753 23.516 ;
      RECT MASK 1 9.771 23.33 9.831 24.106 ;
      RECT MASK 1 10.103 23.335 10.163 23.608 ;
      RECT MASK 1 12.344 23.335 12.404 24.365 ;
      RECT MASK 1 6.056 23.378 6.116 23.645 ;
      RECT MASK 1 6.72 23.378 6.78 23.608 ;
      RECT MASK 1 11.099 23.378 11.159 23.885 ;
      RECT MASK 1 11.431 23.378 11.491 24.562 ;
      RECT MASK 1 5.145 23.554 5.205 24.551 ;
      RECT MASK 1 15.211 23.636 15.271 24.244 ;
      RECT MASK 1 16.539 23.636 16.599 24.244 ;
      RECT MASK 1 17.867 23.636 17.927 24.244 ;
      RECT MASK 1 19.195 23.636 19.255 24.244 ;
      RECT MASK 1 13.34 23.69 13.4 24.21 ;
      RECT MASK 1 11.763 23.728 11.823 24.125 ;
      RECT MASK 1 12.012 23.728 12.072 23.91 ;
      RECT MASK 1 10.103 23.821 10.163 24.562 ;
      RECT MASK 1 10.767 23.825 10.827 24.562 ;
      RECT MASK 1 10.435 23.894 10.495 24.212 ;
      RECT MASK 1 1.076 23.9 1.11 24.5055 ;
      RECT MASK 1 1.295 23.945 1.335 24.5075 ;
      RECT MASK 1 11.099 24.055 11.159 24.562 ;
      RECT MASK 1 14.132 24.1025 14.192 25.2175 ;
      RECT MASK 1 20.44 24.1025 20.5 25.2175 ;
      RECT MASK 1 2.631 24.14 2.665 24.9 ;
      RECT MASK 1 14.713 24.147 14.773 24.956 ;
      RECT MASK 1 15.709 24.147 15.769 24.956 ;
      RECT MASK 1 16.041 24.147 16.101 24.956 ;
      RECT MASK 1 17.037 24.147 17.097 24.956 ;
      RECT MASK 1 17.369 24.147 17.429 24.956 ;
      RECT MASK 1 18.365 24.147 18.425 24.956 ;
      RECT MASK 1 18.697 24.147 18.757 24.956 ;
      RECT MASK 1 19.693 24.147 19.753 24.956 ;
      RECT MASK 1 20.191 24.147 20.251 24.956 ;
      RECT MASK 1 3.074 24.28 3.134 24.9 ;
      RECT MASK 1 11.763 24.33 11.823 25.14 ;
      RECT MASK 1 12.095 24.33 12.155 25.14 ;
      RECT MASK 1 12.676 24.33 12.736 25.14 ;
      RECT MASK 1 13.008 24.33 13.068 25.14 ;
      RECT MASK 1 13.34 24.33 13.4 25.14 ;
      RECT MASK 1 6.056 24.332 6.116 24.605 ;
      RECT MASK 1 6.388 24.332 6.448 24.605 ;
      RECT MASK 1 6.72 24.332 6.78 24.605 ;
      RECT MASK 1 7.052 24.332 7.112 24.605 ;
      RECT MASK 1 7.384 24.332 7.444 24.605 ;
      RECT MASK 1 7.716 24.332 7.776 24.605 ;
      RECT MASK 1 8.048 24.332 8.108 24.605 ;
      RECT MASK 1 8.38 24.332 8.44 24.605 ;
      RECT MASK 1 8.712 24.332 8.772 24.605 ;
      RECT MASK 1 9.044 24.332 9.104 24.605 ;
      RECT MASK 1 9.376 24.332 9.436 24.605 ;
      RECT MASK 1 0.852 24.34 0.892 25.15 ;
      RECT MASK 1 1.516 24.34 1.556 25.15 ;
      RECT MASK 1 15.211 24.364 15.271 24.956 ;
      RECT MASK 1 16.539 24.364 16.599 24.956 ;
      RECT MASK 1 17.867 24.364 17.927 24.956 ;
      RECT MASK 1 19.195 24.364 19.255 24.956 ;
      RECT MASK 1 2.403 24.69 2.437 24.9 ;
      RECT MASK 1 2.859 24.69 2.893 24.9 ;
      RECT MASK 1 21.178 24.81 21.238 25.05 ;
      RECT MASK 1 21.51 24.81 21.57 25.05 ;
      RECT MASK 1 21.842 24.81 21.902 25.05 ;
      RECT MASK 1 22.174 24.81 22.234 25.05 ;
      RECT MASK 1 22.506 24.81 22.566 25.05 ;
      RECT MASK 1 22.838 24.81 22.898 25.05 ;
      RECT MASK 1 23.17 24.81 23.23 25.05 ;
      RECT MASK 1 23.502 24.81 23.562 25.05 ;
      RECT MASK 1 23.834 24.81 23.894 25.05 ;
      RECT MASK 1 24.166 24.81 24.226 25.05 ;
      RECT MASK 1 24.498 24.81 24.558 25.05 ;
      RECT MASK 1 24.83 24.81 24.89 25.05 ;
      RECT MASK 1 25.162 24.81 25.222 25.05 ;
      RECT MASK 1 25.494 24.81 25.554 25.05 ;
      RECT MASK 1 26.398 24.81 26.458 25.05 ;
      RECT MASK 1 26.73 24.81 26.79 25.05 ;
      RECT MASK 1 27.062 24.81 27.122 25.05 ;
      RECT MASK 1 27.394 24.81 27.454 25.05 ;
      RECT MASK 1 27.726 24.81 27.786 25.05 ;
      RECT MASK 1 28.058 24.81 28.118 25.05 ;
      RECT MASK 1 28.39 24.81 28.45 25.05 ;
      RECT MASK 1 28.722 24.81 28.782 25.05 ;
      RECT MASK 1 29.054 24.81 29.114 25.05 ;
      RECT MASK 1 29.386 24.81 29.446 25.05 ;
      RECT MASK 1 29.718 24.81 29.778 25.05 ;
      RECT MASK 1 30.05 24.81 30.11 25.05 ;
      RECT MASK 1 30.382 24.81 30.442 25.05 ;
      RECT MASK 1 30.714 24.81 30.774 25.05 ;
      RECT MASK 1 31.046 24.81 31.106 25.05 ;
      RECT MASK 1 31.378 24.81 31.438 25.05 ;
      RECT MASK 1 1.295 24.835 1.335 25.095 ;
      RECT MASK 1 15.211 25.076 15.271 25.684 ;
      RECT MASK 1 16.539 25.076 16.599 25.684 ;
      RECT MASK 1 17.867 25.076 17.927 25.684 ;
      RECT MASK 1 19.195 25.076 19.255 25.684 ;
      RECT MASK 1 21.849 25.2 21.909 26.64 ;
      RECT MASK 1 22.123 25.2 22.183 26.64 ;
      RECT MASK 1 22.397 25.2 22.457 26.64 ;
      RECT MASK 1 22.671 25.2 22.731 26.64 ;
      RECT MASK 1 22.945 25.2 23.005 26.64 ;
      RECT MASK 1 23.219 25.2 23.279 26.64 ;
      RECT MASK 1 23.493 25.2 23.553 26.64 ;
      RECT MASK 1 23.767 25.2 23.827 26.64 ;
      RECT MASK 1 24.041 25.2 24.101 26.64 ;
      RECT MASK 1 24.315 25.2 24.375 26.64 ;
      RECT MASK 1 24.589 25.2 24.649 26.64 ;
      RECT MASK 1 24.863 25.2 24.923 26.64 ;
      RECT MASK 1 6.774 25.26 6.834 26.64 ;
      RECT MASK 1 7.048 25.26 7.108 26.64 ;
      RECT MASK 1 7.322 25.26 7.382 26.64 ;
      RECT MASK 1 7.596 25.26 7.656 26.64 ;
      RECT MASK 1 7.87 25.26 7.93 26.64 ;
      RECT MASK 1 8.144 25.26 8.204 26.64 ;
      RECT MASK 1 8.418 25.26 8.478 26.64 ;
      RECT MASK 1 8.692 25.26 8.752 26.64 ;
      RECT MASK 1 8.966 25.26 9.026 26.64 ;
      RECT MASK 1 9.24 25.26 9.3 26.64 ;
      RECT MASK 1 9.514 25.26 9.574 26.64 ;
      RECT MASK 1 9.788 25.26 9.848 26.64 ;
      RECT MASK 1 10.062 25.26 10.122 26.64 ;
      RECT MASK 1 10.336 25.26 10.396 26.64 ;
      RECT MASK 1 10.61 25.26 10.67 26.64 ;
      RECT MASK 1 10.884 25.26 10.944 26.64 ;
      RECT MASK 1 11.158 25.26 11.218 26.64 ;
      RECT MASK 1 11.432 25.26 11.492 26.64 ;
      RECT MASK 1 11.706 25.26 11.766 26.64 ;
      RECT MASK 1 11.98 25.26 12.04 26.64 ;
      RECT MASK 1 12.254 25.26 12.314 26.64 ;
      RECT MASK 1 12.528 25.26 12.588 26.64 ;
      RECT MASK 1 14.713 25.5885 14.773 26.46 ;
      RECT MASK 1 15.709 25.5885 15.769 26.46 ;
      RECT MASK 1 16.041 25.5885 16.101 26.46 ;
      RECT MASK 1 17.037 25.5885 17.097 26.46 ;
      RECT MASK 1 17.369 25.5885 17.429 26.46 ;
      RECT MASK 1 18.365 25.5885 18.425 26.46 ;
      RECT MASK 1 18.697 25.5885 18.757 26.46 ;
      RECT MASK 1 19.693 25.5885 19.753 26.46 ;
      RECT MASK 1 20.191 25.5885 20.251 26.46 ;
      RECT MASK 1 15.211 25.804 15.271 26.46 ;
      RECT MASK 1 16.539 25.804 16.599 26.46 ;
      RECT MASK 1 17.867 25.804 17.927 26.46 ;
      RECT MASK 1 19.195 25.804 19.255 26.46 ;
    LAYER M2 SPACING 0 ;
      RECT 0 0 32.604 27.36 ;
    LAYER M1 SPACING 0 ;
      RECT MASK 2 1.346 0.635 1.406 0.865 ;
      RECT MASK 2 1.678 0.635 1.738 0.865 ;
      RECT MASK 2 2.01 0.635 2.07 0.865 ;
      RECT MASK 2 2.342 0.635 2.402 0.865 ;
      RECT MASK 2 2.674 0.635 2.734 0.865 ;
      RECT MASK 2 3.006 0.635 3.066 0.865 ;
      RECT MASK 2 3.338 0.635 3.398 0.865 ;
      RECT MASK 2 3.67 0.635 3.73 0.865 ;
      RECT MASK 2 4.002 0.635 4.062 0.865 ;
      RECT MASK 2 4.334 0.635 4.394 0.865 ;
      RECT MASK 2 4.666 0.635 4.726 0.865 ;
      RECT MASK 2 4.998 0.635 5.058 0.865 ;
      RECT MASK 2 5.33 0.635 5.39 0.865 ;
      RECT MASK 2 5.662 0.635 5.722 0.865 ;
      RECT MASK 2 5.994 0.635 6.054 0.865 ;
      RECT MASK 2 6.326 0.635 6.386 0.865 ;
      RECT MASK 2 6.658 0.635 6.718 0.865 ;
      RECT MASK 2 6.99 0.635 7.05 0.865 ;
      RECT MASK 2 7.322 0.635 7.382 0.865 ;
      RECT MASK 2 7.654 0.635 7.714 0.865 ;
      RECT MASK 2 7.986 0.635 8.046 0.865 ;
      RECT MASK 2 8.318 0.635 8.378 0.865 ;
      RECT MASK 2 8.65 0.635 8.71 0.865 ;
      RECT MASK 2 8.982 0.635 9.042 0.865 ;
      RECT MASK 2 9.314 0.635 9.374 0.865 ;
      RECT MASK 2 9.646 0.635 9.706 0.865 ;
      RECT MASK 2 9.978 0.635 10.038 0.865 ;
      RECT MASK 2 10.31 0.635 10.37 0.865 ;
      RECT MASK 2 10.642 0.635 10.702 0.865 ;
      RECT MASK 2 10.974 0.635 11.034 0.865 ;
      RECT MASK 2 11.306 0.635 11.366 0.865 ;
      RECT MASK 2 11.638 0.635 11.698 0.865 ;
      RECT MASK 2 11.97 0.635 12.03 0.865 ;
      RECT MASK 2 12.302 0.635 12.362 0.865 ;
      RECT MASK 2 12.634 0.635 12.694 0.865 ;
      RECT MASK 2 12.966 0.635 13.026 0.865 ;
      RECT MASK 2 13.298 0.635 13.358 0.865 ;
      RECT MASK 2 13.63 0.635 13.69 0.865 ;
      RECT MASK 2 13.962 0.635 14.022 0.865 ;
      RECT MASK 2 14.294 0.635 14.354 0.865 ;
      RECT MASK 2 14.626 0.635 14.686 0.865 ;
      RECT MASK 2 14.958 0.635 15.018 0.865 ;
      RECT MASK 2 15.29 0.635 15.35 0.865 ;
      RECT MASK 2 15.622 0.635 15.682 0.865 ;
      RECT MASK 2 15.788 0.635 15.848 0.865 ;
      RECT MASK 2 16.12 0.635 16.18 0.865 ;
      RECT MASK 2 16.452 0.635 16.512 0.865 ;
      RECT MASK 2 16.784 0.635 16.844 0.865 ;
      RECT MASK 2 17.116 0.635 17.176 0.865 ;
      RECT MASK 2 17.448 0.635 17.508 0.865 ;
      RECT MASK 2 17.78 0.635 17.84 0.865 ;
      RECT MASK 2 18.112 0.635 18.172 0.865 ;
      RECT MASK 2 18.444 0.635 18.504 0.865 ;
      RECT MASK 2 18.776 0.635 18.836 0.865 ;
      RECT MASK 2 19.108 0.635 19.168 0.865 ;
      RECT MASK 2 19.44 0.635 19.5 0.865 ;
      RECT MASK 2 19.772 0.635 19.832 0.865 ;
      RECT MASK 2 20.104 0.635 20.164 0.865 ;
      RECT MASK 2 20.436 0.635 20.496 0.865 ;
      RECT MASK 2 20.768 0.635 20.828 0.865 ;
      RECT MASK 2 21.1 0.635 21.16 0.865 ;
      RECT MASK 2 21.432 0.635 21.492 0.865 ;
      RECT MASK 2 21.764 0.635 21.824 0.865 ;
      RECT MASK 2 22.096 0.635 22.156 0.865 ;
      RECT MASK 2 22.428 0.635 22.488 0.865 ;
      RECT MASK 2 22.76 0.635 22.82 0.865 ;
      RECT MASK 2 23.092 0.635 23.152 0.865 ;
      RECT MASK 2 23.424 0.635 23.484 0.865 ;
      RECT MASK 2 23.756 0.635 23.816 0.865 ;
      RECT MASK 2 24.088 0.635 24.148 0.865 ;
      RECT MASK 2 24.42 0.635 24.48 0.865 ;
      RECT MASK 2 24.752 0.635 24.812 0.865 ;
      RECT MASK 2 25.084 0.635 25.144 0.865 ;
      RECT MASK 2 25.416 0.635 25.476 0.865 ;
      RECT MASK 2 25.748 0.635 25.808 0.865 ;
      RECT MASK 2 26.08 0.635 26.14 0.865 ;
      RECT MASK 2 26.412 0.635 26.472 0.865 ;
      RECT MASK 2 26.744 0.635 26.804 0.865 ;
      RECT MASK 2 27.076 0.635 27.136 0.865 ;
      RECT MASK 2 27.408 0.635 27.468 0.865 ;
      RECT MASK 2 27.74 0.635 27.8 0.865 ;
      RECT MASK 2 29.48 0.71 29.52 1.541 ;
      RECT MASK 2 30.144 0.71 30.184 1.541 ;
      RECT MASK 2 30.808 0.71 30.848 1.541 ;
      RECT MASK 2 31.472 0.71 31.512 1.541 ;
      RECT MASK 2 31.251 0.96 31.291 7.255 ;
      RECT MASK 2 31.693 1 31.733 7.735 ;
      RECT MASK 2 29.259 1.189 29.299 7.255 ;
      RECT MASK 2 29.701 1.189 29.741 7.735 ;
      RECT MASK 2 29.923 1.189 29.963 7.255 ;
      RECT MASK 2 30.365 1.189 30.405 7.735 ;
      RECT MASK 2 30.587 1.189 30.627 7.255 ;
      RECT MASK 2 31.029 1.189 31.069 7.735 ;
      RECT MASK 2 29.48 1.579 29.52 6.33 ;
      RECT MASK 2 30.144 1.579 30.184 6.33 ;
      RECT MASK 2 30.808 1.579 30.848 6.33 ;
      RECT MASK 2 31.472 1.579 31.512 6.33 ;
      RECT MASK 2 29.48 7.145 29.52 7.37 ;
      RECT MASK 2 30.144 7.145 30.184 7.37 ;
      RECT MASK 2 30.808 7.145 30.848 7.37 ;
      RECT MASK 2 31.472 7.145 31.512 7.37 ;
      RECT MASK 2 29.48 7.625 29.52 7.85 ;
      RECT MASK 2 30.144 7.625 30.184 7.85 ;
      RECT MASK 2 30.808 7.625 30.848 7.85 ;
      RECT MASK 2 31.472 7.625 31.512 7.85 ;
      RECT MASK 2 29.48 8.225 29.52 9.775 ;
      RECT MASK 2 30.144 8.225 30.184 9.775 ;
      RECT MASK 2 30.808 8.225 30.848 9.775 ;
      RECT MASK 2 31.472 8.225 31.512 9.775 ;
      RECT MASK 2 1.9605 9.1995 2.0205 9.695 ;
      RECT MASK 2 2.738 9.1995 2.798 9.575 ;
      RECT MASK 2 3.512 9.1995 3.572 9.695 ;
      RECT MASK 2 14.74 9.1995 14.8 9.575 ;
      RECT MASK 2 15.455 9.1995 15.515 10.445 ;
      RECT MASK 2 7.82 9.385 7.88 15.025 ;
      RECT MASK 2 8.152 9.385 8.212 15.025 ;
      RECT MASK 2 4.226 9.505 4.286 12.065 ;
      RECT MASK 2 1.18 9.875 1.24 10.105 ;
      RECT MASK 2 1.512 9.875 1.572 10.105 ;
      RECT MASK 2 1.844 9.875 1.904 10.105 ;
      RECT MASK 2 2.176 9.875 2.236 10.105 ;
      RECT MASK 2 2.508 9.875 2.568 10.105 ;
      RECT MASK 2 2.84 9.875 2.9 10.105 ;
      RECT MASK 2 3.172 9.875 3.232 10.105 ;
      RECT MASK 2 3.504 9.875 3.564 10.105 ;
      RECT MASK 2 3.836 9.875 3.896 10.105 ;
      RECT MASK 2 4.5 9.875 4.56 10.105 ;
      RECT MASK 2 4.832 9.875 4.892 10.105 ;
      RECT MASK 2 5.164 9.875 5.224 10.105 ;
      RECT MASK 2 5.496 9.875 5.556 10.105 ;
      RECT MASK 2 5.828 9.875 5.888 10.105 ;
      RECT MASK 2 6.16 9.875 6.22 10.105 ;
      RECT MASK 2 6.492 9.875 6.552 10.105 ;
      RECT MASK 2 6.824 9.875 6.884 10.105 ;
      RECT MASK 2 7.156 9.875 7.216 10.105 ;
      RECT MASK 2 7.488 9.875 7.548 10.105 ;
      RECT MASK 2 8.318 9.875 8.378 10.105 ;
      RECT MASK 2 8.65 9.875 8.71 10.105 ;
      RECT MASK 2 8.982 9.875 9.042 10.105 ;
      RECT MASK 2 9.314 9.875 9.374 10.105 ;
      RECT MASK 2 9.646 9.875 9.706 10.105 ;
      RECT MASK 2 9.978 9.875 10.038 10.105 ;
      RECT MASK 2 10.31 9.875 10.37 10.105 ;
      RECT MASK 2 10.642 9.875 10.702 10.105 ;
      RECT MASK 2 10.974 9.875 11.034 10.105 ;
      RECT MASK 2 11.306 9.875 11.366 10.105 ;
      RECT MASK 2 11.638 9.875 11.698 10.105 ;
      RECT MASK 2 11.97 9.875 12.03 10.105 ;
      RECT MASK 2 12.302 9.875 12.362 10.105 ;
      RECT MASK 2 12.634 9.875 12.694 10.105 ;
      RECT MASK 2 12.966 9.875 13.026 10.105 ;
      RECT MASK 2 13.298 9.875 13.358 10.105 ;
      RECT MASK 2 13.63 9.875 13.69 10.105 ;
      RECT MASK 2 13.962 9.875 14.022 10.105 ;
      RECT MASK 2 14.294 9.875 14.354 10.105 ;
      RECT MASK 2 14.626 9.875 14.686 10.105 ;
      RECT MASK 2 14.958 9.875 15.018 10.105 ;
      RECT MASK 2 15.29 9.875 15.35 10.105 ;
      RECT MASK 2 15.788 9.875 15.848 10.105 ;
      RECT MASK 2 16.12 9.875 16.18 10.105 ;
      RECT MASK 2 16.452 9.875 16.512 10.105 ;
      RECT MASK 2 16.784 9.875 16.844 10.105 ;
      RECT MASK 2 17.116 9.875 17.176 10.105 ;
      RECT MASK 2 17.448 9.875 17.508 10.105 ;
      RECT MASK 2 17.78 9.875 17.84 10.105 ;
      RECT MASK 2 18.112 9.875 18.172 10.105 ;
      RECT MASK 2 18.444 9.875 18.504 10.105 ;
      RECT MASK 2 18.776 9.875 18.836 10.105 ;
      RECT MASK 2 19.108 9.875 19.168 10.105 ;
      RECT MASK 2 19.44 9.875 19.5 10.105 ;
      RECT MASK 2 19.772 9.875 19.832 10.105 ;
      RECT MASK 2 20.104 9.875 20.164 10.105 ;
      RECT MASK 2 20.436 9.875 20.496 10.105 ;
      RECT MASK 2 20.768 9.875 20.828 10.105 ;
      RECT MASK 2 21.1 9.875 21.16 10.105 ;
      RECT MASK 2 21.432 9.875 21.492 10.105 ;
      RECT MASK 2 21.764 9.875 21.824 10.105 ;
      RECT MASK 2 22.096 9.875 22.156 10.105 ;
      RECT MASK 2 22.428 9.875 22.488 10.105 ;
      RECT MASK 2 22.76 9.875 22.82 10.105 ;
      RECT MASK 2 23.092 9.875 23.152 10.105 ;
      RECT MASK 2 23.424 9.875 23.484 10.105 ;
      RECT MASK 2 23.756 9.875 23.816 10.105 ;
      RECT MASK 2 24.088 9.875 24.148 10.105 ;
      RECT MASK 2 24.42 9.875 24.48 10.105 ;
      RECT MASK 2 24.752 9.875 24.812 10.105 ;
      RECT MASK 2 25.084 9.875 25.144 10.105 ;
      RECT MASK 2 25.416 9.875 25.476 10.105 ;
      RECT MASK 2 25.748 9.875 25.808 10.105 ;
      RECT MASK 2 26.08 9.875 26.14 10.105 ;
      RECT MASK 2 26.412 9.875 26.472 10.105 ;
      RECT MASK 2 26.744 9.875 26.804 10.105 ;
      RECT MASK 2 27.076 9.875 27.136 10.105 ;
      RECT MASK 2 27.408 9.875 27.468 10.105 ;
      RECT MASK 2 27.74 9.875 27.8 10.105 ;
      RECT MASK 2 0.838 10.29 0.918 12.54 ;
      RECT MASK 2 1.058 10.295 1.118 10.525 ;
      RECT MASK 2 1.346 10.295 1.406 10.525 ;
      RECT MASK 2 1.634 10.295 1.694 12.565 ;
      RECT MASK 2 1.922 10.295 1.982 12.565 ;
      RECT MASK 2 2.21 10.295 2.27 12.565 ;
      RECT MASK 2 2.498 10.295 2.558 10.525 ;
      RECT MASK 2 2.786 10.295 2.846 12.565 ;
      RECT MASK 2 3.074 10.295 3.134 10.525 ;
      RECT MASK 2 3.362 10.295 3.422 12.565 ;
      RECT MASK 2 3.65 10.295 3.71 10.525 ;
      RECT MASK 2 3.938 10.295 3.998 12.565 ;
      RECT MASK 2 4.514 10.295 4.574 10.525 ;
      RECT MASK 2 4.802 10.295 4.862 12.565 ;
      RECT MASK 2 5.09 10.295 5.15 10.525 ;
      RECT MASK 2 5.378 10.295 5.438 10.525 ;
      RECT MASK 2 5.666 10.295 5.726 12.565 ;
      RECT MASK 2 5.954 10.295 6.014 10.525 ;
      RECT MASK 2 6.242 10.295 6.302 10.525 ;
      RECT MASK 2 6.53 10.295 6.59 12.565 ;
      RECT MASK 2 6.818 10.295 6.878 11.509 ;
      RECT MASK 2 7.106 10.295 7.166 12.565 ;
      RECT MASK 2 7.394 10.295 7.454 12.565 ;
      RECT MASK 2 8.484 10.295 8.544 12.565 ;
      RECT MASK 2 8.816 10.295 8.876 10.525 ;
      RECT MASK 2 9.148 10.295 9.208 10.525 ;
      RECT MASK 2 9.48 10.295 9.54 12.565 ;
      RECT MASK 2 9.812 10.295 9.872 10.525 ;
      RECT MASK 2 25.791 10.295 25.851 12.42 ;
      RECT MASK 2 26.065 10.295 26.125 12.42 ;
      RECT MASK 2 26.339 10.295 26.399 12.42 ;
      RECT MASK 2 26.613 10.295 26.673 12.42 ;
      RECT MASK 2 26.887 10.295 26.947 12.42 ;
      RECT MASK 2 27.161 10.295 27.221 12.42 ;
      RECT MASK 2 24.984 10.5 25.064 12.21 ;
      RECT MASK 2 27.972 10.5 28.052 12.21 ;
      RECT MASK 2 11.935 10.693 11.995 10.941 ;
      RECT MASK 2 12.433 10.693 12.493 10.941 ;
      RECT MASK 2 14.923 10.75 14.983 10.941 ;
      RECT MASK 2 16.5 10.752 16.56 10.941 ;
      RECT MASK 2 16.749 10.752 16.809 10.941 ;
      RECT MASK 2 17.911 10.752 17.971 10.941 ;
      RECT MASK 2 18.243 10.752 18.303 10.941 ;
      RECT MASK 2 18.658 10.752 18.718 10.946 ;
      RECT MASK 2 19.82 10.752 19.88 10.946 ;
      RECT MASK 2 20.65 10.752 20.71 10.946 ;
      RECT MASK 2 21.812 10.752 21.872 10.946 ;
      RECT MASK 2 22.642 10.752 22.702 11.2385 ;
      RECT MASK 2 23.804 10.752 23.864 11.2385 ;
      RECT MASK 2 2.498 10.928 2.558 11.152 ;
      RECT MASK 2 3.074 10.928 3.134 11.152 ;
      RECT MASK 2 3.65 10.928 3.71 11.152 ;
      RECT MASK 2 4.514 10.928 4.574 11.945 ;
      RECT MASK 2 5.09 10.928 5.15 11.945 ;
      RECT MASK 2 5.378 10.928 5.438 12.065 ;
      RECT MASK 2 5.954 10.928 6.014 11.932 ;
      RECT MASK 2 6.242 10.928 6.302 11.932 ;
      RECT MASK 2 8.816 10.928 8.876 14.392 ;
      RECT MASK 2 9.148 10.928 9.208 14.392 ;
      RECT MASK 2 12.931 10.958 12.991 11.782 ;
      RECT MASK 2 13.263 10.958 13.323 11.782 ;
      RECT MASK 2 13.595 10.958 13.655 11.782 ;
      RECT MASK 2 13.927 10.958 13.987 11.782 ;
      RECT MASK 2 14.425 10.958 14.485 11.782 ;
      RECT MASK 2 15.421 10.958 15.481 11.782 ;
      RECT MASK 2 15.753 10.958 15.813 11.782 ;
      RECT MASK 2 16.085 10.958 16.145 11.782 ;
      RECT MASK 2 17.413 10.958 17.473 11.782 ;
      RECT MASK 2 20.235 10.958 20.295 11.782 ;
      RECT MASK 2 22.227 10.958 22.287 11.782 ;
      RECT MASK 2 24.219 10.958 24.279 11.782 ;
      RECT MASK 2 4.658 11.035 4.718 11.825 ;
      RECT MASK 2 4.946 11.035 5.006 11.825 ;
      RECT MASK 2 11.935 11.061 11.995 11.679 ;
      RECT MASK 2 12.433 11.061 12.493 11.679 ;
      RECT MASK 2 14.923 11.061 14.983 11.679 ;
      RECT MASK 2 17.911 11.061 17.971 11.679 ;
      RECT MASK 2 16.749 11.217 16.809 11.615 ;
      RECT MASK 2 6.962 11.275 7.022 11.585 ;
      RECT MASK 2 16.417 11.378 16.477 11.615 ;
      RECT MASK 2 2.498 11.708 2.558 11.932 ;
      RECT MASK 2 3.074 11.708 3.134 11.932 ;
      RECT MASK 2 3.65 11.708 3.71 11.932 ;
      RECT MASK 2 6.818 11.708 6.878 11.932 ;
      RECT MASK 2 18.658 11.794 18.718 11.988 ;
      RECT MASK 2 19.82 11.794 19.88 11.988 ;
      RECT MASK 2 20.65 11.794 20.71 11.988 ;
      RECT MASK 2 21.812 11.794 21.872 11.988 ;
      RECT MASK 2 22.642 11.794 22.702 11.988 ;
      RECT MASK 2 23.804 11.794 23.864 11.988 ;
      RECT MASK 2 11.935 11.799 11.995 12.047 ;
      RECT MASK 2 12.433 11.799 12.493 12.047 ;
      RECT MASK 2 14.923 11.799 14.983 11.99 ;
      RECT MASK 2 16.5 11.799 16.56 11.988 ;
      RECT MASK 2 16.749 11.799 16.809 11.988 ;
      RECT MASK 2 17.911 11.799 17.971 11.988 ;
      RECT MASK 2 18.243 11.799 18.303 11.988 ;
      RECT MASK 2 1.058 12.335 1.118 12.565 ;
      RECT MASK 2 1.346 12.335 1.406 12.565 ;
      RECT MASK 2 2.498 12.335 2.558 12.565 ;
      RECT MASK 2 3.074 12.335 3.134 12.565 ;
      RECT MASK 2 3.65 12.335 3.71 12.565 ;
      RECT MASK 2 4.226 12.335 4.286 12.565 ;
      RECT MASK 2 4.514 12.335 4.574 12.565 ;
      RECT MASK 2 5.09 12.335 5.15 12.565 ;
      RECT MASK 2 5.378 12.335 5.438 12.565 ;
      RECT MASK 2 5.954 12.335 6.014 12.565 ;
      RECT MASK 2 6.242 12.335 6.302 12.565 ;
      RECT MASK 2 6.818 12.335 6.878 12.565 ;
      RECT MASK 2 9.812 12.335 9.872 12.565 ;
      RECT MASK 2 21.344 12.63 21.404 12.87 ;
      RECT MASK 2 21.676 12.63 21.736 15.64 ;
      RECT MASK 2 22.008 12.63 22.068 12.87 ;
      RECT MASK 2 22.34 12.63 22.4 12.87 ;
      RECT MASK 2 22.672 12.63 22.732 12.87 ;
      RECT MASK 2 23.004 12.63 23.064 12.87 ;
      RECT MASK 2 23.336 12.63 23.396 12.87 ;
      RECT MASK 2 23.668 12.63 23.728 12.87 ;
      RECT MASK 2 24 12.63 24.06 12.87 ;
      RECT MASK 2 24.332 12.63 24.392 12.87 ;
      RECT MASK 2 24.664 12.63 24.724 12.87 ;
      RECT MASK 2 24.996 12.63 25.056 15.64 ;
      RECT MASK 2 25.65 12.63 25.73 25.05 ;
      RECT MASK 2 26.222 12.63 26.302 25.05 ;
      RECT MASK 2 26.398 12.63 26.458 12.87 ;
      RECT MASK 2 27.062 12.63 27.122 12.87 ;
      RECT MASK 2 27.394 12.63 27.454 12.87 ;
      RECT MASK 2 27.726 12.63 27.786 12.87 ;
      RECT MASK 2 28.058 12.63 28.118 12.87 ;
      RECT MASK 2 28.39 12.63 28.45 12.87 ;
      RECT MASK 2 28.722 12.63 28.782 12.87 ;
      RECT MASK 2 29.054 12.63 29.114 12.87 ;
      RECT MASK 2 29.386 12.63 29.446 12.87 ;
      RECT MASK 2 29.718 12.63 29.778 12.87 ;
      RECT MASK 2 30.05 12.63 30.11 12.87 ;
      RECT MASK 2 30.382 12.63 30.442 12.87 ;
      RECT MASK 2 30.714 12.63 30.774 12.87 ;
      RECT MASK 2 31.046 12.63 31.106 12.87 ;
      RECT MASK 2 31.378 12.63 31.438 12.87 ;
      RECT MASK 2 31.7 12.63 31.78 25.05 ;
      RECT MASK 2 1.058 12.73 1.118 12.985 ;
      RECT MASK 2 1.346 12.73 1.406 12.985 ;
      RECT MASK 2 1.634 12.73 1.694 15.025 ;
      RECT MASK 2 1.922 12.73 1.982 15.025 ;
      RECT MASK 2 2.21 12.73 2.27 15.025 ;
      RECT MASK 2 2.498 12.73 2.558 15.025 ;
      RECT MASK 2 2.786 12.73 2.846 13.612 ;
      RECT MASK 2 3.074 12.73 3.134 15.025 ;
      RECT MASK 2 3.362 12.73 3.422 15.025 ;
      RECT MASK 2 3.65 12.73 3.71 12.985 ;
      RECT MASK 2 3.938 12.73 3.998 12.985 ;
      RECT MASK 2 4.226 12.73 4.286 12.985 ;
      RECT MASK 2 4.514 12.73 4.574 15.025 ;
      RECT MASK 2 4.802 12.73 4.862 12.985 ;
      RECT MASK 2 5.09 12.73 5.15 12.985 ;
      RECT MASK 2 5.378 12.73 5.438 15.025 ;
      RECT MASK 2 5.666 12.73 5.726 12.985 ;
      RECT MASK 2 5.954 12.73 6.014 12.985 ;
      RECT MASK 2 6.242 12.73 6.302 12.985 ;
      RECT MASK 2 6.53 12.73 6.59 15.025 ;
      RECT MASK 2 6.818 12.73 6.878 13.612 ;
      RECT MASK 2 7.106 12.73 7.166 15.025 ;
      RECT MASK 2 7.394 12.73 7.454 15.025 ;
      RECT MASK 2 8.484 12.73 8.544 15.025 ;
      RECT MASK 2 9.48 12.73 9.54 15.025 ;
      RECT MASK 2 9.812 12.73 9.872 12.985 ;
      RECT MASK 2 20.806 13.0575 20.866 22.5 ;
      RECT MASK 2 13.696 13.135 13.756 14.705 ;
      RECT MASK 2 22.672 13.15 22.732 15.64 ;
      RECT MASK 2 24 13.15 24.06 15.64 ;
      RECT MASK 2 14.766 13.17 14.826 17.37 ;
      RECT MASK 2 15.91 13.17 15.97 17.37 ;
      RECT MASK 2 16.242 13.17 16.302 13.532 ;
      RECT MASK 2 16.574 13.17 16.634 17.37 ;
      RECT MASK 2 22.008 13.25 22.068 15.54 ;
      RECT MASK 2 24.664 13.25 24.724 15.54 ;
      RECT MASK 2 12.368 13.26 12.428 13.985 ;
      RECT MASK 2 12.7 13.26 12.76 14.088 ;
      RECT MASK 2 13.032 13.26 13.092 13.985 ;
      RECT MASK 2 13.364 13.26 13.424 14.1475 ;
      RECT MASK 2 15.338 13.26 15.398 14.1475 ;
      RECT MASK 2 18.353 13.34 18.387 13.65 ;
      RECT MASK 2 18.553 13.34 18.587 13.65 ;
      RECT MASK 2 18.753 13.34 18.787 13.65 ;
      RECT MASK 2 18.953 13.34 18.987 13.65 ;
      RECT MASK 2 19.153 13.34 19.187 13.65 ;
      RECT MASK 2 19.353 13.34 19.387 13.65 ;
      RECT MASK 2 19.54 13.34 19.6 13.59 ;
      RECT MASK 2 3.65 13.388 3.71 14.392 ;
      RECT MASK 2 3.938 13.388 3.998 14.392 ;
      RECT MASK 2 4.226 13.388 4.286 14.392 ;
      RECT MASK 2 4.802 13.388 4.862 14.392 ;
      RECT MASK 2 5.09 13.388 5.15 14.392 ;
      RECT MASK 2 5.666 13.388 5.726 13.612 ;
      RECT MASK 2 5.954 13.388 6.014 13.612 ;
      RECT MASK 2 6.242 13.388 6.302 14.392 ;
      RECT MASK 2 23.336 13.45 23.396 15.34 ;
      RECT MASK 2 22.34 13.55 22.4 15.24 ;
      RECT MASK 2 6.098 13.751 6.158 14.285 ;
      RECT MASK 2 14.268 13.838 14.328 14.124 ;
      RECT MASK 2 14.6 13.838 14.66 14.124 ;
      RECT MASK 2 16.076 13.838 16.136 14.105 ;
      RECT MASK 2 16.408 13.838 16.468 14.105 ;
      RECT MASK 2 19.14 13.955 19.2 14.935 ;
      RECT MASK 2 18.24 13.96 18.3 14.845 ;
      RECT MASK 2 18.84 13.96 18.9 14.845 ;
      RECT MASK 2 15.504 14.03 15.564 14.825 ;
      RECT MASK 2 17.426 14.0325 17.486 14.8595 ;
      RECT MASK 2 19.54 14.045 19.6 14.845 ;
      RECT MASK 2 12.368 14.105 12.428 14.755 ;
      RECT MASK 2 2.786 14.168 2.846 14.392 ;
      RECT MASK 2 5.666 14.168 5.726 14.392 ;
      RECT MASK 2 5.954 14.168 6.014 14.392 ;
      RECT MASK 2 6.818 14.168 6.878 14.392 ;
      RECT MASK 2 14.434 14.188 14.494 14.571 ;
      RECT MASK 2 17.94 14.188 18 14.6965 ;
      RECT MASK 2 14.268 14.289 14.328 14.672 ;
      RECT MASK 2 27.3345 14.3445 27.4345 23.3435 ;
      RECT MASK 2 14.6 14.39 14.66 15.065 ;
      RECT MASK 2 13.364 14.7125 13.424 15.8275 ;
      RECT MASK 2 15.338 14.7125 15.398 15.8275 ;
      RECT MASK 2 17.94 14.7345 18 15.065 ;
      RECT MASK 2 16.076 14.755 16.136 15.022 ;
      RECT MASK 2 16.408 14.755 16.468 15.022 ;
      RECT MASK 2 12.7 14.772 12.76 15.768 ;
      RECT MASK 2 14.268 14.792 14.328 15.748 ;
      RECT MASK 2 17.632 14.792 17.692 15.748 ;
      RECT MASK 2 1.058 14.795 1.118 15.025 ;
      RECT MASK 2 1.346 14.795 1.406 15.025 ;
      RECT MASK 2 2.786 14.795 2.846 15.025 ;
      RECT MASK 2 3.65 14.795 3.71 15.025 ;
      RECT MASK 2 3.938 14.795 3.998 15.025 ;
      RECT MASK 2 4.226 14.795 4.286 15.025 ;
      RECT MASK 2 4.802 14.795 4.862 15.025 ;
      RECT MASK 2 5.09 14.795 5.15 15.025 ;
      RECT MASK 2 5.666 14.795 5.726 15.025 ;
      RECT MASK 2 5.954 14.795 6.014 15.025 ;
      RECT MASK 2 6.242 14.795 6.302 15.025 ;
      RECT MASK 2 6.818 14.795 6.878 15.025 ;
      RECT MASK 2 7.654 14.795 7.714 15.025 ;
      RECT MASK 2 8.816 14.795 8.876 15.025 ;
      RECT MASK 2 9.148 14.795 9.208 15.025 ;
      RECT MASK 2 9.812 14.795 9.872 15.025 ;
      RECT MASK 2 12.368 14.875 12.428 15.665 ;
      RECT MASK 2 13.032 14.875 13.092 15.665 ;
      RECT MASK 2 18.353 15.21 18.387 15.33 ;
      RECT MASK 2 18.553 15.21 18.587 15.33 ;
      RECT MASK 2 18.753 15.21 18.787 15.33 ;
      RECT MASK 2 18.953 15.21 18.987 15.33 ;
      RECT MASK 2 19.453 15.21 19.487 15.33 ;
      RECT MASK 2 14.6 15.475 14.66 16.15 ;
      RECT MASK 2 17.94 15.475 18 15.8055 ;
      RECT MASK 2 16.076 15.518 16.136 15.785 ;
      RECT MASK 2 16.408 15.518 16.468 15.785 ;
      RECT MASK 2 19.14 15.605 19.2 16.585 ;
      RECT MASK 2 17.426 15.6805 17.486 16.5075 ;
      RECT MASK 2 18.24 15.695 18.3 16.58 ;
      RECT MASK 2 18.84 15.695 18.9 16.58 ;
      RECT MASK 2 19.54 15.695 19.6 16.495 ;
      RECT MASK 2 15.504 15.715 15.564 16.51 ;
      RECT MASK 2 2.855 15.75 2.915 20.37 ;
      RECT MASK 2 3.129 15.75 3.189 20.37 ;
      RECT MASK 2 3.403 15.75 3.463 20.37 ;
      RECT MASK 2 3.677 15.75 3.737 20.37 ;
      RECT MASK 2 3.951 15.75 4.011 20.37 ;
      RECT MASK 2 4.225 15.75 4.285 20.37 ;
      RECT MASK 2 4.499 15.75 4.559 18.847 ;
      RECT MASK 2 4.773 15.75 4.833 18.847 ;
      RECT MASK 2 5.047 15.75 5.107 18.847 ;
      RECT MASK 2 5.321 15.75 5.381 18.847 ;
      RECT MASK 2 5.595 15.75 5.655 18.847 ;
      RECT MASK 2 5.869 15.75 5.929 18.847 ;
      RECT MASK 2 6.143 15.75 6.203 18.815 ;
      RECT MASK 2 6.417 15.75 6.477 17.277 ;
      RECT MASK 2 6.691 15.75 6.751 17.277 ;
      RECT MASK 2 6.965 15.75 7.025 17.277 ;
      RECT MASK 2 7.239 15.75 7.299 17.277 ;
      RECT MASK 2 7.513 15.75 7.573 17.277 ;
      RECT MASK 2 7.787 15.75 7.847 17.277 ;
      RECT MASK 2 8.061 15.75 8.121 17.277 ;
      RECT MASK 2 8.335 15.75 8.395 17.277 ;
      RECT MASK 2 8.609 15.75 8.669 17.277 ;
      RECT MASK 2 8.883 15.75 8.943 17.277 ;
      RECT MASK 2 9.157 15.75 9.217 17.277 ;
      RECT MASK 2 9.431 15.75 9.491 17.277 ;
      RECT MASK 2 9.705 15.75 9.765 17.277 ;
      RECT MASK 2 9.979 15.75 10.039 17.277 ;
      RECT MASK 2 10.253 15.75 10.313 17.245 ;
      RECT MASK 2 12.368 15.785 12.428 16.435 ;
      RECT MASK 2 17.94 15.8435 18 16.352 ;
      RECT MASK 2 14.268 15.868 14.328 16.251 ;
      RECT MASK 2 21.676 15.87 21.736 16.15 ;
      RECT MASK 2 22.672 15.87 22.732 20.06 ;
      RECT MASK 2 23.336 15.87 23.396 16.15 ;
      RECT MASK 2 24 15.87 24.06 16.15 ;
      RECT MASK 2 24.332 15.87 24.392 16.15 ;
      RECT MASK 2 24.664 15.87 24.724 16.15 ;
      RECT MASK 2 24.996 15.87 25.056 16.15 ;
      RECT MASK 2 14.434 15.969 14.494 16.352 ;
      RECT MASK 2 22.008 15.97 22.068 17.1 ;
      RECT MASK 2 22.34 15.97 22.4 20.56 ;
      RECT MASK 2 1.184 16.085 1.224 17.635 ;
      RECT MASK 2 23.004 16.17 23.064 16.9 ;
      RECT MASK 2 13.364 16.3925 13.424 17.28 ;
      RECT MASK 2 15.338 16.3925 15.398 17.28 ;
      RECT MASK 2 14.268 16.416 14.328 16.702 ;
      RECT MASK 2 14.6 16.416 14.66 16.702 ;
      RECT MASK 2 16.076 16.435 16.136 16.702 ;
      RECT MASK 2 16.408 16.435 16.468 16.702 ;
      RECT MASK 2 12.7 16.452 12.76 17.28 ;
      RECT MASK 2 12.368 16.555 12.428 17.28 ;
      RECT MASK 2 13.032 16.555 13.092 17.28 ;
      RECT MASK 2 18.353 16.89 18.387 17.2 ;
      RECT MASK 2 18.553 16.89 18.587 17.2 ;
      RECT MASK 2 18.753 16.89 18.787 17.2 ;
      RECT MASK 2 18.953 16.89 18.987 17.2 ;
      RECT MASK 2 19.153 16.89 19.187 17.2 ;
      RECT MASK 2 19.353 16.89 19.387 17.2 ;
      RECT MASK 2 21.676 16.92 21.736 18.37 ;
      RECT MASK 2 23.336 16.92 23.396 17.61 ;
      RECT MASK 2 24 16.92 24.06 17.61 ;
      RECT MASK 2 24.332 16.92 24.392 17.61 ;
      RECT MASK 2 24.664 16.92 24.724 17.61 ;
      RECT MASK 2 24.996 16.92 25.056 17.61 ;
      RECT MASK 2 19.54 16.95 19.6 17.2 ;
      RECT MASK 2 16.242 17.008 16.302 17.37 ;
      RECT MASK 2 22.008 17.37 22.068 18.275 ;
      RECT MASK 2 23.004 17.37 23.064 18.275 ;
      RECT MASK 2 6.82 17.675 6.86 20.565 ;
      RECT MASK 2 1.184 18.01 1.224 18.235 ;
      RECT MASK 2 7.533 18.017 7.593 18.713 ;
      RECT MASK 2 8.031 18.017 8.091 18.713 ;
      RECT MASK 2 8.529 18.017 8.589 18.713 ;
      RECT MASK 2 8.861 18.017 8.921 18.947 ;
      RECT MASK 2 1.405 18.125 1.445 24.671 ;
      RECT MASK 2 1.184 18.49 1.224 18.715 ;
      RECT MASK 2 21.676 18.54 21.736 18.82 ;
      RECT MASK 2 0.963 18.605 1.003 24.671 ;
      RECT MASK 2 9.193 18.716 9.253 19.225 ;
      RECT MASK 2 7.533 18.895 7.593 19.385 ;
      RECT MASK 2 8.031 18.895 8.091 19.385 ;
      RECT MASK 2 8.529 18.895 8.589 19.385 ;
      RECT MASK 2 9.94 18.895 10 19.385 ;
      RECT MASK 2 11.268 18.895 11.328 19.385 ;
      RECT MASK 2 12.596 18.895 12.656 19.385 ;
      RECT MASK 2 13.924 18.895 13.984 19.385 ;
      RECT MASK 2 15.252 18.895 15.312 19.385 ;
      RECT MASK 2 16.58 18.895 16.64 19.385 ;
      RECT MASK 2 17.908 18.895 17.968 19.385 ;
      RECT MASK 2 19.236 18.895 19.296 19.385 ;
      RECT MASK 2 5.602 19.31 5.642 20.49 ;
      RECT MASK 2 5.802 19.31 5.842 19.87 ;
      RECT MASK 2 6.002 19.31 6.042 19.87 ;
      RECT MASK 2 6.202 19.31 6.242 20.565 ;
      RECT MASK 2 20.44 19.357 20.5 21.002 ;
      RECT MASK 2 8.861 19.367 8.921 20.261 ;
      RECT MASK 2 9.193 19.472 9.253 20.261 ;
      RECT MASK 2 21.676 19.52 21.736 19.8 ;
      RECT MASK 2 1.184 19.53 1.224 24.281 ;
      RECT MASK 2 7.533 19.569 7.593 20.261 ;
      RECT MASK 2 8.031 19.569 8.091 20.261 ;
      RECT MASK 2 8.529 19.569 8.589 20.261 ;
      RECT MASK 2 21.676 19.98 21.736 20.97 ;
      RECT MASK 2 22.008 20.125 22.068 20.97 ;
      RECT MASK 2 23.004 20.125 23.064 20.97 ;
      RECT MASK 2 23.336 20.125 23.396 20.97 ;
      RECT MASK 2 18.448 20.292 18.508 21.472 ;
      RECT MASK 2 14.132 20.381 14.192 21.0725 ;
      RECT MASK 2 14.381 20.381 14.441 20.997 ;
      RECT MASK 2 14.713 20.381 14.773 20.997 ;
      RECT MASK 2 15.211 20.381 15.271 20.997 ;
      RECT MASK 2 15.543 20.381 15.603 20.631 ;
      RECT MASK 2 15.875 20.381 15.935 20.997 ;
      RECT MASK 2 16.29 20.381 16.35 21.002 ;
      RECT MASK 2 16.788 20.381 16.848 21.002 ;
      RECT MASK 2 15.045 20.648 15.105 21.472 ;
      RECT MASK 2 17.203 20.648 17.263 21.472 ;
      RECT MASK 2 19.776 20.648 19.836 21.472 ;
      RECT MASK 2 6.222 20.7 6.282 21.51 ;
      RECT MASK 2 6.554 20.7 6.614 21.51 ;
      RECT MASK 2 6.886 20.7 6.946 21.51 ;
      RECT MASK 2 7.218 20.7 7.278 21.51 ;
      RECT MASK 2 7.55 20.7 7.61 21.51 ;
      RECT MASK 2 7.882 20.7 7.942 21.51 ;
      RECT MASK 2 8.214 20.7 8.274 21.51 ;
      RECT MASK 2 8.546 20.7 8.606 21.51 ;
      RECT MASK 2 8.878 20.7 8.938 21.51 ;
      RECT MASK 2 9.21 20.7 9.27 21.51 ;
      RECT MASK 2 10.601 20.7 10.661 21.508 ;
      RECT MASK 2 11.265 20.7 11.325 21.51 ;
      RECT MASK 2 11.597 20.7 11.657 21.51 ;
      RECT MASK 2 22.34 20.73 22.4 20.97 ;
      RECT MASK 2 22.672 20.73 22.732 20.97 ;
      RECT MASK 2 24 20.73 24.06 20.97 ;
      RECT MASK 2 24.332 20.73 24.392 20.97 ;
      RECT MASK 2 24.664 20.73 24.724 20.97 ;
      RECT MASK 2 24.996 20.73 25.056 20.97 ;
      RECT MASK 2 15.543 20.751 15.603 21.369 ;
      RECT MASK 2 17.784 20.815 17.844 21.305 ;
      RECT MASK 2 19.112 20.815 19.172 21.305 ;
      RECT MASK 2 2.237 20.94 2.297 21.56 ;
      RECT MASK 2 2.517 20.94 2.551 21.15 ;
      RECT MASK 2 2.745 20.94 2.779 21.15 ;
      RECT MASK 2 9.937 21.235 9.997 22.107 ;
      RECT MASK 2 12.215 21.235 12.275 21.703 ;
      RECT MASK 2 12.51 21.235 12.57 22.462 ;
      RECT MASK 2 12.842 21.235 12.902 22.462 ;
      RECT MASK 2 4.104 21.278 4.164 22.558 ;
      RECT MASK 2 5.33 21.278 5.39 22.558 ;
      RECT MASK 2 9.542 21.278 9.602 21.545 ;
      RECT MASK 2 10.269 21.278 10.329 22.797 ;
      RECT MASK 2 11.929 21.278 11.989 21.545 ;
      RECT MASK 2 13.174 21.278 13.234 22.462 ;
      RECT MASK 2 2.789 21.31 2.849 22.34 ;
      RECT MASK 2 5.828 21.392 5.888 21.931 ;
      RECT MASK 2 2.447 21.4 2.507 22.43 ;
      RECT MASK 2 14.547 21.484 14.607 22.309 ;
      RECT MASK 2 15.211 21.484 15.271 22.309 ;
      RECT MASK 2 16.29 21.484 16.35 22.309 ;
      RECT MASK 2 16.788 21.484 16.848 22.309 ;
      RECT MASK 2 15.543 21.489 15.603 22.071 ;
      RECT MASK 2 15.875 21.489 15.935 22.071 ;
      RECT MASK 2 17.203 21.592 17.263 21.968 ;
      RECT MASK 2 9.293 21.633 9.353 22.006 ;
      RECT MASK 2 6.222 21.729 6.282 22.107 ;
      RECT MASK 2 10.933 21.734 10.993 22.107 ;
      RECT MASK 2 11.265 21.734 11.325 22.006 ;
      RECT MASK 2 14.879 21.882 14.939 22.071 ;
      RECT MASK 2 22.63 21.8915 22.69 22.82 ;
      RECT MASK 2 22.83 21.8915 22.89 22.82 ;
      RECT MASK 2 24.03 21.898 24.09 22.82 ;
      RECT MASK 2 23.83 21.9005 23.89 22.82 ;
      RECT MASK 2 5.662 21.931 5.722 22.317 ;
      RECT MASK 2 5.828 22.052 5.888 22.317 ;
      RECT MASK 2 17.203 22.088 17.263 22.912 ;
      RECT MASK 2 18.448 22.088 18.508 22.912 ;
      RECT MASK 2 19.776 22.088 19.836 22.912 ;
      RECT MASK 2 23.568 22.1755 23.628 23.6825 ;
      RECT MASK 2 11.597 22.19 11.657 23.65 ;
      RECT MASK 2 14.879 22.191 14.939 22.809 ;
      RECT MASK 2 15.543 22.191 15.603 22.809 ;
      RECT MASK 2 11.265 22.195 11.325 23.645 ;
      RECT MASK 2 6.222 22.232 6.282 22.505 ;
      RECT MASK 2 6.554 22.232 6.614 22.505 ;
      RECT MASK 2 6.886 22.232 6.946 22.505 ;
      RECT MASK 2 7.218 22.232 7.278 22.505 ;
      RECT MASK 2 7.55 22.232 7.61 22.505 ;
      RECT MASK 2 7.882 22.232 7.942 22.505 ;
      RECT MASK 2 8.214 22.232 8.274 22.505 ;
      RECT MASK 2 8.546 22.232 8.606 22.505 ;
      RECT MASK 2 8.878 22.232 8.938 22.505 ;
      RECT MASK 2 9.21 22.232 9.27 22.505 ;
      RECT MASK 2 9.542 22.232 9.602 22.505 ;
      RECT MASK 2 11.929 22.232 11.989 22.505 ;
      RECT MASK 2 17.784 22.255 17.844 22.745 ;
      RECT MASK 2 19.112 22.255 19.172 22.745 ;
      RECT MASK 2 13.672 22.425 13.732 23.885 ;
      RECT MASK 2 4.647 22.427 4.707 22.835 ;
      RECT MASK 2 4.979 22.427 5.039 22.835 ;
      RECT MASK 2 2.517 22.59 2.551 22.8 ;
      RECT MASK 2 2.745 22.59 2.779 22.8 ;
      RECT MASK 2 14.132 22.6625 14.192 23.7775 ;
      RECT MASK 2 20.44 22.6625 20.5 23.7775 ;
      RECT MASK 2 14.535 22.685 14.595 23.516 ;
      RECT MASK 2 15.211 22.685 15.271 23.118 ;
      RECT MASK 2 15.875 22.685 15.935 23.179 ;
      RECT MASK 2 16.29 22.685 16.35 23.516 ;
      RECT MASK 2 16.788 22.685 16.848 23.516 ;
      RECT MASK 2 20.108 22.685 20.168 23.516 ;
      RECT MASK 2 14.879 22.929 14.939 23.118 ;
      RECT MASK 2 15.543 22.929 15.603 23.179 ;
      RECT MASK 2 22.63 23 22.69 23.8845 ;
      RECT MASK 2 22.83 23 22.89 23.8845 ;
      RECT MASK 2 23.83 23 23.89 23.8815 ;
      RECT MASK 2 24.03 23 24.09 23.8815 ;
      RECT MASK 2 4.647 23.005 4.707 23.413 ;
      RECT MASK 2 4.979 23.005 5.039 23.413 ;
      RECT MASK 2 2.517 23.04 2.551 23.25 ;
      RECT MASK 2 2.745 23.04 2.779 23.25 ;
      RECT MASK 2 10.269 23.043 10.329 24.562 ;
      RECT MASK 2 14.962 23.261 15.022 23.516 ;
      RECT MASK 2 4.104 23.282 4.164 24.562 ;
      RECT MASK 2 5.33 23.282 5.39 24.562 ;
      RECT MASK 2 15.46 23.322 15.52 23.516 ;
      RECT MASK 2 17.618 23.322 17.678 23.516 ;
      RECT MASK 2 18.116 23.322 18.176 23.516 ;
      RECT MASK 2 18.946 23.322 19.006 23.516 ;
      RECT MASK 2 19.444 23.322 19.504 23.516 ;
      RECT MASK 2 6.222 23.335 6.282 23.608 ;
      RECT MASK 2 6.554 23.335 6.614 23.608 ;
      RECT MASK 2 6.886 23.335 6.946 23.608 ;
      RECT MASK 2 7.218 23.335 7.278 23.608 ;
      RECT MASK 2 7.55 23.335 7.61 23.608 ;
      RECT MASK 2 7.882 23.335 7.942 23.608 ;
      RECT MASK 2 8.214 23.335 8.274 23.608 ;
      RECT MASK 2 8.546 23.335 8.606 23.608 ;
      RECT MASK 2 8.878 23.335 8.938 23.608 ;
      RECT MASK 2 9.21 23.335 9.27 23.608 ;
      RECT MASK 2 9.542 23.335 9.602 23.608 ;
      RECT MASK 2 11.929 23.335 11.989 23.608 ;
      RECT MASK 2 12.51 23.378 12.57 24.562 ;
      RECT MASK 2 12.842 23.378 12.902 24.562 ;
      RECT MASK 2 13.174 23.378 13.234 24.562 ;
      RECT MASK 2 2.447 23.41 2.507 24.44 ;
      RECT MASK 2 2.789 23.5 2.849 24.53 ;
      RECT MASK 2 5.662 23.523 5.722 23.909 ;
      RECT MASK 2 5.828 23.523 5.888 23.788 ;
      RECT MASK 2 15.875 23.528 15.935 25.792 ;
      RECT MASK 2 17.203 23.528 17.263 25.792 ;
      RECT MASK 2 18.531 23.528 18.591 25.792 ;
      RECT MASK 2 19.859 23.528 19.919 25.792 ;
      RECT MASK 2 6.222 23.733 6.282 24.111 ;
      RECT MASK 2 9.937 23.733 9.997 24.605 ;
      RECT MASK 2 10.933 23.733 10.993 24.106 ;
      RECT MASK 2 9.293 23.834 9.353 24.207 ;
      RECT MASK 2 11.265 23.834 11.325 24.106 ;
      RECT MASK 2 5.828 23.909 5.888 24.448 ;
      RECT MASK 2 12.215 24.137 12.275 24.605 ;
      RECT MASK 2 14.962 24.147 15.022 24.956 ;
      RECT MASK 2 15.46 24.147 15.52 24.956 ;
      RECT MASK 2 16.29 24.147 16.35 24.956 ;
      RECT MASK 2 16.788 24.147 16.848 24.956 ;
      RECT MASK 2 17.618 24.147 17.678 24.956 ;
      RECT MASK 2 18.116 24.147 18.176 24.956 ;
      RECT MASK 2 18.946 24.147 19.006 24.956 ;
      RECT MASK 2 19.444 24.147 19.504 24.956 ;
      RECT MASK 2 2.237 24.28 2.297 24.9 ;
      RECT MASK 2 9.542 24.295 9.602 24.562 ;
      RECT MASK 2 11.929 24.295 11.989 24.562 ;
      RECT MASK 2 1.184 24.319 1.224 25.08 ;
      RECT MASK 2 6.222 24.33 6.282 25.14 ;
      RECT MASK 2 6.554 24.33 6.614 25.14 ;
      RECT MASK 2 6.886 24.33 6.946 25.14 ;
      RECT MASK 2 7.218 24.33 7.278 25.14 ;
      RECT MASK 2 7.55 24.33 7.61 25.14 ;
      RECT MASK 2 7.882 24.33 7.942 25.14 ;
      RECT MASK 2 8.214 24.33 8.274 25.14 ;
      RECT MASK 2 8.546 24.33 8.606 25.14 ;
      RECT MASK 2 8.878 24.33 8.938 25.14 ;
      RECT MASK 2 9.21 24.33 9.27 25.14 ;
      RECT MASK 2 11.265 24.33 11.325 25.14 ;
      RECT MASK 2 11.597 24.33 11.657 25.14 ;
      RECT MASK 2 10.601 24.332 10.661 25.14 ;
      RECT MASK 2 2.517 24.69 2.551 24.9 ;
      RECT MASK 2 2.745 24.69 2.779 24.9 ;
      RECT MASK 2 21.344 24.81 21.404 25.05 ;
      RECT MASK 2 21.676 24.81 21.736 25.05 ;
      RECT MASK 2 22.008 24.81 22.068 25.05 ;
      RECT MASK 2 22.34 24.81 22.4 25.05 ;
      RECT MASK 2 22.672 24.81 22.732 25.05 ;
      RECT MASK 2 23.004 24.81 23.064 25.05 ;
      RECT MASK 2 23.336 24.81 23.396 25.05 ;
      RECT MASK 2 23.668 24.81 23.728 25.05 ;
      RECT MASK 2 24 24.81 24.06 25.05 ;
      RECT MASK 2 24.332 24.81 24.392 25.05 ;
      RECT MASK 2 24.664 24.81 24.724 25.05 ;
      RECT MASK 2 24.996 24.81 25.056 25.05 ;
      RECT MASK 2 25.328 24.81 25.388 25.05 ;
      RECT MASK 2 26.564 24.81 26.624 25.05 ;
      RECT MASK 2 26.896 24.81 26.956 25.05 ;
      RECT MASK 2 27.228 24.81 27.288 25.05 ;
      RECT MASK 2 27.56 24.81 27.62 25.05 ;
      RECT MASK 2 27.892 24.81 27.952 25.05 ;
      RECT MASK 2 28.224 24.81 28.284 25.05 ;
      RECT MASK 2 28.556 24.81 28.616 25.05 ;
      RECT MASK 2 28.888 24.81 28.948 25.05 ;
      RECT MASK 2 29.22 24.81 29.28 25.05 ;
      RECT MASK 2 29.552 24.81 29.612 25.05 ;
      RECT MASK 2 29.884 24.81 29.944 25.05 ;
      RECT MASK 2 30.216 24.81 30.276 25.05 ;
      RECT MASK 2 30.548 24.81 30.608 25.05 ;
      RECT MASK 2 30.88 24.81 30.94 25.05 ;
      RECT MASK 2 31.212 24.81 31.272 25.05 ;
      RECT MASK 2 31.544 24.81 31.604 25.05 ;
      RECT MASK 2 21.986 25.2 22.046 26.892 ;
      RECT MASK 2 22.26 25.2 22.32 26.892 ;
      RECT MASK 2 22.534 25.2 22.594 26.892 ;
      RECT MASK 2 22.808 25.2 22.868 26.892 ;
      RECT MASK 2 23.082 25.2 23.142 26.892 ;
      RECT MASK 2 23.356 25.2 23.416 26.892 ;
      RECT MASK 2 23.63 25.2 23.69 26.892 ;
      RECT MASK 2 23.904 25.2 23.964 26.892 ;
      RECT MASK 2 24.178 25.2 24.238 26.892 ;
      RECT MASK 2 24.452 25.2 24.512 26.892 ;
      RECT MASK 2 24.726 25.2 24.786 26.892 ;
      RECT MASK 2 21.026 25.255 21.086 26.892 ;
      RECT MASK 2 25.526 25.255 25.586 26.892 ;
      RECT MASK 2 6.911 25.26 6.971 26.924 ;
      RECT MASK 2 7.185 25.26 7.245 26.924 ;
      RECT MASK 2 7.459 25.26 7.519 26.924 ;
      RECT MASK 2 7.733 25.26 7.793 26.924 ;
      RECT MASK 2 8.007 25.26 8.067 26.924 ;
      RECT MASK 2 8.281 25.26 8.341 26.924 ;
      RECT MASK 2 8.555 25.26 8.615 26.924 ;
      RECT MASK 2 8.829 25.26 8.889 26.924 ;
      RECT MASK 2 9.103 25.26 9.163 26.924 ;
      RECT MASK 2 9.377 25.26 9.437 26.924 ;
      RECT MASK 2 9.651 25.26 9.711 26.924 ;
      RECT MASK 2 9.925 25.26 9.985 26.924 ;
      RECT MASK 2 10.199 25.26 10.259 26.924 ;
      RECT MASK 2 10.473 25.26 10.533 26.924 ;
      RECT MASK 2 10.747 25.26 10.807 26.924 ;
      RECT MASK 2 11.021 25.26 11.081 26.924 ;
      RECT MASK 2 11.295 25.26 11.355 26.924 ;
      RECT MASK 2 11.569 25.26 11.629 26.924 ;
      RECT MASK 2 11.843 25.26 11.903 26.924 ;
      RECT MASK 2 12.117 25.26 12.177 26.924 ;
      RECT MASK 2 12.391 25.26 12.451 26.924 ;
      RECT MASK 2 6.038 25.309 6.098 26.924 ;
      RECT MASK 2 13.238 25.309 13.298 26.924 ;
      RECT MASK 2 14.132 25.5425 14.192 26.46 ;
      RECT MASK 2 20.44 25.5425 20.5 26.46 ;
      RECT MASK 2 14.962 25.5885 15.022 26.46 ;
      RECT MASK 2 15.46 25.5885 15.52 26.46 ;
      RECT MASK 2 16.29 25.5885 16.35 26.46 ;
      RECT MASK 2 16.788 25.5885 16.848 26.46 ;
      RECT MASK 2 17.618 25.5885 17.678 26.46 ;
      RECT MASK 2 18.116 25.5885 18.176 26.46 ;
      RECT MASK 2 18.946 25.5885 19.006 26.46 ;
      RECT MASK 2 19.444 25.5885 19.504 26.46 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 1 29.072 0.73 32.4235 0.77 ;
      RECT MASK 1 29.072 1.05 32.4235 1.09 ;
      RECT MASK 1 30.013 1.3 31.52 1.36 ;
      RECT MASK 1 0.43 1.47 28.388 1.53 ;
      RECT MASK 1 29.072 1.66 32.4235 1.7 ;
      RECT MASK 1 0.43 2.19 28.388 2.25 ;
      RECT MASK 1 29.072 2.24 32.4235 2.28 ;
      RECT MASK 1 0.43 2.91 28.388 2.97 ;
      RECT MASK 1 0.43 3.63 28.388 3.69 ;
      RECT MASK 1 0.43 4.35 28.388 4.41 ;
      RECT MASK 1 0.43 5.07 28.388 5.13 ;
      RECT MASK 1 29.072 5.25 32.4235 5.31 ;
      RECT MASK 1 29.072 5.73 32.4235 5.79 ;
      RECT MASK 1 0.43 5.79 28.388 5.85 ;
      RECT MASK 1 29.072 6.21 32.4235 6.27 ;
      RECT MASK 1 0.43 6.51 28.388 6.57 ;
      RECT MASK 1 29.244 7.17 29.535 7.23 ;
      RECT MASK 1 29.908 7.17 30.199 7.23 ;
      RECT MASK 1 30.572 7.17 30.863 7.23 ;
      RECT MASK 1 31.236 7.17 31.527 7.23 ;
      RECT MASK 1 0.43 7.23 28.388 7.29 ;
      RECT MASK 1 29.465 7.65 29.761 7.71 ;
      RECT MASK 1 30.129 7.65 30.425 7.71 ;
      RECT MASK 1 30.793 7.65 31.089 7.71 ;
      RECT MASK 1 31.457 7.65 31.753 7.71 ;
      RECT MASK 1 0.43 7.95 28.388 8.01 ;
      RECT MASK 1 28.9785 8.13 31.859 8.19 ;
      RECT MASK 1 0.43 8.67 28.388 8.73 ;
      RECT MASK 1 28.9785 8.73 32.4235 8.79 ;
      RECT MASK 1 13.653 9.15 17.352 9.21 ;
      RECT MASK 1 30.468 9.27 31.532 9.33 ;
      RECT MASK 1 1.926 9.39 14.92 9.45 ;
      RECT MASK 1 17.242 9.51 29.646 9.57 ;
      RECT MASK 1 30.732 9.51 31.064 9.57 ;
      RECT MASK 1 1.926 9.63 14.92 9.69 ;
      RECT MASK 1 10.627 10.26 15.54 10.32 ;
      RECT MASK 1 0.684 10.32 10.254 10.5 ;
      RECT MASK 1 10.627 10.5 15.54 10.56 ;
      RECT MASK 1 2.442 11.04 5.0325 11.1 ;
      RECT MASK 1 12.408 11.206 12.767 11.246 ;
      RECT MASK 1 13.072 11.206 13.763 11.246 ;
      RECT MASK 1 14.896 11.206 30.8415 11.246 ;
      RECT MASK 1 0.774 11.28 11.081 11.34 ;
      RECT MASK 1 13.57 11.398 13.846 11.438 ;
      RECT MASK 1 14.483 11.398 15.5205 11.438 ;
      RECT MASK 1 15.728 11.398 16.502 11.438 ;
      RECT MASK 1 16.89 11.398 17.332 11.438 ;
      RECT MASK 1 24.194 11.398 31.79 11.438 ;
      RECT MASK 1 12.065 11.473 12.369 11.533 ;
      RECT MASK 1 0.774 11.52 11.081 11.58 ;
      RECT MASK 1 17.388 11.583 17.996 11.623 ;
      RECT MASK 1 20.21 11.583 27.784 11.623 ;
      RECT MASK 1 14.4 11.586 16.668 11.626 ;
      RECT MASK 1 2.448 11.76 5.0325 11.82 ;
      RECT MASK 1 5.786 11.76 8.0795 11.82 ;
      RECT MASK 1 11.55 11.806 32.4105 11.996 ;
      RECT MASK 1 4.0575 12 6.189 12.06 ;
      RECT MASK 1 11.55 12.235 32.4105 12.425 ;
      RECT MASK 1 8.764 12.6 11.247 12.66 ;
      RECT MASK 1 20.603 12.66 32.3865 12.84 ;
      RECT MASK 1 13.676 13.14 14.593 13.2 ;
      RECT MASK 1 21.49 13.63 31.0865 13.73 ;
      RECT MASK 1 3.6115 13.74 11.084 13.8 ;
      RECT MASK 1 15.89 13.8 17.1905 13.86 ;
      RECT MASK 1 3.6115 13.98 11.084 14.04 ;
      RECT MASK 1 14.224 14.04 15.745 14.1 ;
      RECT MASK 1 16.056 14.04 17.524 14.1 ;
      RECT MASK 1 3.6115 14.22 4.911 14.28 ;
      RECT MASK 1 6.034 14.22 8.0795 14.28 ;
      RECT MASK 1 2.61 14.2205 2.8765 14.2805 ;
      RECT MASK 1 20.992 14.35 32.35 14.45 ;
      RECT MASK 1 13.178 14.52 18.32 14.58 ;
      RECT MASK 1 18.815 14.52 20.178 14.58 ;
      RECT MASK 1 17.786 14.74 20.401 14.8 ;
      RECT MASK 1 13.971 14.76 15.629 14.82 ;
      RECT MASK 1 16.0505 14.76 17.3205 14.82 ;
      RECT MASK 1 14.58 15 18.023 15.06 ;
      RECT MASK 1 18.7275 15.02 20.401 15.08 ;
      RECT MASK 1 21.49 15.07 31.0865 15.17 ;
      RECT MASK 1 3.433 15.39 10.583 15.57 ;
      RECT MASK 1 18.7225 15.46 20.401 15.52 ;
      RECT MASK 1 14.58 15.48 18.023 15.54 ;
      RECT MASK 1 1.2725 15.51 3.02 15.57 ;
      RECT MASK 1 13.971 15.72 15.629 15.78 ;
      RECT MASK 1 16.0505 15.72 17.3205 15.78 ;
      RECT MASK 1 17.786 15.74 20.401 15.8 ;
      RECT MASK 1 2.088 16.095 10.583 16.275 ;
      RECT MASK 1 13.178 16.2 18.32 16.26 ;
      RECT MASK 1 18.815 16.2 20.178 16.26 ;
      RECT MASK 1 14.224 16.44 15.745 16.5 ;
      RECT MASK 1 16.056 16.44 17.524 16.5 ;
      RECT MASK 1 2.693 16.5 11.081 16.56 ;
      RECT MASK 1 21.988 16.53 22.752 16.59 ;
      RECT MASK 1 15.89 16.68 17.1905 16.74 ;
      RECT MASK 1 2.693 16.74 11.081 16.8 ;
      RECT MASK 1 21.3765 16.99 32.35 17.09 ;
      RECT MASK 1 0.635 17.07 1.7 17.13 ;
      RECT MASK 1 2.088 17.1 10.583 17.28 ;
      RECT MASK 1 21.3765 17.4 32.35 17.58 ;
      RECT MASK 1 0.635 17.67 1.7 17.73 ;
      RECT MASK 1 5.075 17.84 20.894 17.9 ;
      RECT MASK 1 1.169 18.15 1.465 18.21 ;
      RECT MASK 1 21.3765 18.19 32.35 18.29 ;
      RECT MASK 1 2.088 18.285 6.614 18.465 ;
      RECT MASK 1 7.148 18.317 20.606 18.397 ;
      RECT MASK 1 23.15 18.43 27.4345 18.53 ;
      RECT MASK 1 0.948 18.63 1.239 18.69 ;
      RECT MASK 1 20.992 18.67 32.35 18.77 ;
      RECT MASK 1 10.5435 19.127 20.1785 19.187 ;
      RECT MASK 1 5.482 19.19 6.803 19.27 ;
      RECT MASK 1 2.088 19.275 4.724 19.455 ;
      RECT MASK 1 7.148 19.474 20.636 19.664 ;
      RECT MASK 1 5.762 19.58 6.0775 19.6 ;
      RECT MASK 1 0.829 19.59 1.884 19.65 ;
      RECT MASK 1 20.992 19.63 32.35 19.73 ;
      RECT MASK 1 5.472 19.75 6.803 19.83 ;
      RECT MASK 1 7.148 19.864 20.636 20.054 ;
      RECT MASK 1 23.15 19.87 27.4345 19.97 ;
      RECT MASK 1 2.088 19.875 4.724 20.055 ;
      RECT MASK 1 0.829 20.07 1.884 20.13 ;
      RECT MASK 1 5.472 20.07 6.803 20.15 ;
      RECT MASK 1 20.988 20.11 32.35 20.21 ;
      RECT MASK 1 13.865 20.422 20.636 20.622 ;
      RECT MASK 1 3.463 20.515 6.88 20.535 ;
      RECT MASK 1 0.829 20.55 1.884 20.61 ;
      RECT MASK 1 21.656 20.76 25.076 20.94 ;
      RECT MASK 1 9.905 20.802 19.944 20.862 ;
      RECT MASK 1 17.178 21.1455 19.28 21.2055 ;
      RECT MASK 1 6.036 21.24 12.295 21.3 ;
      RECT MASK 1 12.485 21.24 15.088 21.3 ;
      RECT MASK 1 15.606 21.246 16.619 21.306 ;
      RECT MASK 1 9.522 21.48 10.349 21.54 ;
      RECT MASK 1 11.83 21.48 12.425 21.54 ;
      RECT MASK 1 2.769 21.66 5.415 21.72 ;
      RECT MASK 1 10.416 21.72 12.009 21.78 ;
      RECT MASK 1 13.315 21.75 20.837 21.81 ;
      RECT MASK 1 4.245 21.96 6.057 22.02 ;
      RECT MASK 1 9.917 21.96 12.172 22.02 ;
      RECT MASK 1 1.963 22.08 3.3865 22.14 ;
      RECT MASK 1 13.865 22.195 20.636 22.255 ;
      RECT MASK 1 3.61 22.2 13.444 22.26 ;
      RECT MASK 1 13.647 22.435 15.13 22.495 ;
      RECT MASK 1 15.5195 22.435 20.886 22.495 ;
      RECT MASK 1 6.2 22.44 10.1925 22.5 ;
      RECT MASK 1 11.909 22.44 12.452 22.5 ;
      RECT MASK 1 12.651 22.44 13.429 22.5 ;
      RECT MASK 1 13.87 22.695 20.636 22.755 ;
      RECT MASK 1 13.87 22.938 20.636 23.138 ;
      RECT MASK 1 22.46 22.965 24.26 23.145 ;
      RECT MASK 1 13.87 23.318 20.636 23.518 ;
      RECT MASK 1 6.2 23.34 10.1925 23.4 ;
      RECT MASK 1 11.909 23.34 12.452 23.4 ;
      RECT MASK 1 12.651 23.34 13.429 23.4 ;
      RECT MASK 1 0.829 23.58 1.536 23.62 ;
      RECT MASK 1 3.61 23.58 13.444 23.64 ;
      RECT MASK 1 1.963 23.62 3.3865 23.68 ;
      RECT MASK 1 15.1085 23.7025 20.753 23.7625 ;
      RECT MASK 1 4.245 23.82 6.057 23.88 ;
      RECT MASK 1 9.917 23.82 12.172 23.88 ;
      RECT MASK 1 12.485 23.82 13.752 23.88 ;
      RECT MASK 1 1.0445 23.92 1.453 23.96 ;
      RECT MASK 1 15.1085 23.9425 20.753 24.0025 ;
      RECT MASK 1 10.416 24.06 12.009 24.12 ;
      RECT MASK 1 2.769 24.12 5.415 24.18 ;
      RECT MASK 1 0.829 24.16 1.884 24.2 ;
      RECT MASK 1 14.055 24.1825 20.636 24.2425 ;
      RECT MASK 1 9.522 24.3 10.349 24.36 ;
      RECT MASK 1 11.83 24.3 12.425 24.36 ;
      RECT MASK 1 6.036 24.54 12.295 24.6 ;
      RECT MASK 1 13.87 24.63 20.636 24.69 ;
      RECT MASK 1 20.9895 24.84 32.129 25.02 ;
      RECT MASK 1 15.1085 25.2625 20.753 25.3225 ;
      RECT MASK 1 15.1085 25.5025 20.753 25.5625 ;
      RECT MASK 1 3.4385 25.818 31.308 25.998 ;
      RECT MASK 1 3.4385 26.212 31.308 26.402 ;
    LAYER M3 SPACING 0 ;
      RECT 0 0 32.604 27.36 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 2 0.608 0.66 28.388 0.84 ;
      RECT MASK 2 29.072 0.89 32.4235 0.93 ;
      RECT MASK 2 0.43 1.11 28.388 1.17 ;
      RECT MASK 2 29.349 1.18 29.895 1.24 ;
      RECT MASK 2 30.677 1.18 31.785 1.24 ;
      RECT MASK 2 30.583 1.42 31.421 1.48 ;
      RECT MASK 2 29.072 1.74 31.824 1.78 ;
      RECT MASK 2 0.43 1.83 28.388 1.89 ;
      RECT MASK 2 0.43 2.55 28.388 2.61 ;
      RECT MASK 2 29.072 2.73 32.4235 2.79 ;
      RECT MASK 2 29.072 3.21 32.4235 3.27 ;
      RECT MASK 2 0.43 3.27 28.388 3.33 ;
      RECT MASK 2 29.072 3.45 32.4235 3.51 ;
      RECT MASK 2 29.072 3.69 32.4235 3.75 ;
      RECT MASK 2 0.43 3.99 28.388 4.05 ;
      RECT MASK 2 29.072 4.41 32.4235 4.47 ;
      RECT MASK 2 29.072 4.65 32.4235 4.71 ;
      RECT MASK 2 0.43 4.71 28.388 4.77 ;
      RECT MASK 2 29.072 4.89 32.4235 4.95 ;
      RECT MASK 2 0.43 5.43 28.388 5.49 ;
      RECT MASK 2 0.43 6.15 28.388 6.21 ;
      RECT MASK 2 28.9785 6.57 32.4235 6.63 ;
      RECT MASK 2 0.43 6.87 28.388 6.93 ;
      RECT MASK 2 28.9785 7.05 32.4235 7.11 ;
      RECT MASK 2 28.9785 7.53 32.4235 7.59 ;
      RECT MASK 2 0.43 7.59 28.388 7.65 ;
      RECT MASK 2 28.9785 8.01 32.4235 8.07 ;
      RECT MASK 2 0.43 8.31 28.388 8.37 ;
      RECT MASK 2 29.46 8.91 30.863 8.97 ;
      RECT MASK 2 0.43 9.03 28.388 9.09 ;
      RECT MASK 2 29.072 9.09 32.4235 9.15 ;
      RECT MASK 2 12.657 9.27 30.31 9.33 ;
      RECT MASK 2 2.7085 9.51 4.3135 9.57 ;
      RECT MASK 2 7.958 9.51 14.835 9.57 ;
      RECT MASK 2 29.81 9.63 31.643 9.69 ;
      RECT MASK 2 29.072 9.81 32.4235 9.87 ;
      RECT MASK 2 0.608 9.9 28.388 10.08 ;
      RECT MASK 2 15.867 10.32 28.53 10.5 ;
      RECT MASK 2 10.627 10.38 15.54 10.44 ;
      RECT MASK 2 29.072 10.41 32.4235 10.47 ;
      RECT MASK 2 11.55 10.752 32.4105 10.932 ;
      RECT MASK 2 11.137 11.112 16.004 11.152 ;
      RECT MASK 2 22.111 11.112 26.2175 11.152 ;
      RECT MASK 2 4.1815 11.16 6.272 11.22 ;
      RECT MASK 2 14.227 11.3 29.899 11.34 ;
      RECT MASK 2 12.906 11.302 13.67 11.342 ;
      RECT MASK 2 6.207 11.4 11.081 11.46 ;
      RECT MASK 2 17.989 11.487 21.3495 11.527 ;
      RECT MASK 2 22.202 11.489 23.308 11.529 ;
      RECT MASK 2 13.487 11.49 14.8505 11.53 ;
      RECT MASK 2 16.06 11.494 16.9715 11.534 ;
      RECT MASK 2 11.91 11.593 12.894 11.653 ;
      RECT MASK 2 4.305 11.64 5.342 11.7 ;
      RECT MASK 2 5.786 11.64 8.305 11.7 ;
      RECT MASK 2 4.479 11.88 5.187 11.94 ;
      RECT MASK 2 5.786 11.88 8.305 11.94 ;
      RECT MASK 2 11.55 12.074 32.4105 12.154 ;
      RECT MASK 2 0.635 12.36 11.081 12.54 ;
      RECT MASK 2 0.635 12.72 10.9725 12.9 ;
      RECT MASK 2 20.782 13.0625 30.557 13.1225 ;
      RECT MASK 2 13.4045 13.26 13.6795 13.32 ;
      RECT MASK 2 20.992 13.27 32.35 13.37 ;
      RECT MASK 2 12.164 13.5 15.581 13.68 ;
      RECT MASK 2 15.885 13.5 17.285 13.68 ;
      RECT MASK 2 17.628 13.5 19.876 13.68 ;
      RECT MASK 2 3.6115 13.86 10.931 13.92 ;
      RECT MASK 2 12.164 13.92 19.876 13.98 ;
      RECT MASK 2 20.992 13.99 32.35 14.09 ;
      RECT MASK 2 0.635 14.1 10.254 14.16 ;
      RECT MASK 2 16.2205 14.16 17.635 14.22 ;
      RECT MASK 2 0.635 14.34 10.254 14.4 ;
      RECT MASK 2 16.715 14.4 17.373 14.46 ;
      RECT MASK 2 17.9105 14.4 18.5375 14.46 ;
      RECT MASK 2 16.2205 14.6395 17.6795 14.6995 ;
      RECT MASK 2 12.348 14.64 13.776 14.7 ;
      RECT MASK 2 20.992 14.71 32.35 14.81 ;
      RECT MASK 2 0.635 14.82 10.254 15 ;
      RECT MASK 2 11.975 14.88 13.607 14.94 ;
      RECT MASK 2 13.916 14.88 14.846 14.94 ;
      RECT MASK 2 15.188 14.88 20.401 14.94 ;
      RECT MASK 2 11.975 15.18 13.607 15.36 ;
      RECT MASK 2 13.911 15.18 14.851 15.36 ;
      RECT MASK 2 15.188 15.18 20.401 15.36 ;
      RECT MASK 2 0.824 15.39 1.889 15.45 ;
      RECT MASK 2 20.992 15.43 32.35 15.53 ;
      RECT MASK 2 11.975 15.6 13.607 15.66 ;
      RECT MASK 2 13.916 15.6 14.846 15.66 ;
      RECT MASK 2 15.188 15.6 20.401 15.66 ;
      RECT MASK 2 16.2205 15.8405 17.6795 15.9005 ;
      RECT MASK 2 20.992 15.91 32.35 16.01 ;
      RECT MASK 2 0.824 15.99 1.889 16.05 ;
      RECT MASK 2 12.348 16.08 13.61 16.14 ;
      RECT MASK 2 16.715 16.08 17.373 16.14 ;
      RECT MASK 2 17.9105 16.08 18.5375 16.14 ;
      RECT MASK 2 16.2205 16.32 17.635 16.38 ;
      RECT MASK 2 1.169 16.38 12.885 16.44 ;
      RECT MASK 2 20.6605 16.41 23.089 16.47 ;
      RECT MASK 2 12.278 16.56 19.876 16.62 ;
      RECT MASK 2 2.693 16.62 11.081 16.68 ;
      RECT MASK 2 0.824 16.71 1.889 16.77 ;
      RECT MASK 2 12.278 16.86 15.581 17.04 ;
      RECT MASK 2 15.885 16.86 17.285 17.04 ;
      RECT MASK 2 17.628 16.86 19.876 17.04 ;
      RECT MASK 2 2.088 17.4 6.614 17.58 ;
      RECT MASK 2 6.805 17.7 13.278 17.76 ;
      RECT MASK 2 0.837 17.79 1.571 17.85 ;
      RECT MASK 2 7.148 18.007 20.606 18.197 ;
      RECT MASK 2 0.635 18.27 1.7 18.33 ;
      RECT MASK 2 7.148 18.628 20.606 18.818 ;
      RECT MASK 2 2.088 18.67 6.614 18.85 ;
      RECT MASK 2 0.635 18.75 1.7 18.81 ;
      RECT MASK 2 7.3385 19.007 9.3445 19.067 ;
      RECT MASK 2 10.5435 19.007 20.1785 19.067 ;
      RECT MASK 2 5.472 19.03 6.803 19.11 ;
      RECT MASK 2 0.635 19.23 1.7 19.29 ;
      RECT MASK 2 9.905 19.247 18.721 19.307 ;
      RECT MASK 2 5.472 19.35 6.803 19.43 ;
      RECT MASK 2 7.148 19.724 20.636 19.804 ;
      RECT MASK 2 5.482 19.91 6.803 19.99 ;
      RECT MASK 2 7.148 20.114 20.636 20.174 ;
      RECT MASK 2 9.905 20.302 18.721 20.362 ;
      RECT MASK 2 3.048 20.44 5.671 20.46 ;
      RECT MASK 2 13.865 20.682 20.636 20.742 ;
      RECT MASK 2 0.829 20.91 1.884 20.97 ;
      RECT MASK 2 13.865 20.922 20.636 21.002 ;
      RECT MASK 2 2.202 20.94 13.6395 21.12 ;
      RECT MASK 2 15.025 21.126 15.706 21.186 ;
      RECT MASK 2 0.829 21.15 1.884 21.21 ;
      RECT MASK 2 2.217 21.36 13.7215 21.42 ;
      RECT MASK 2 0.829 21.39 1.884 21.45 ;
      RECT MASK 2 13.865 21.478 20.837 21.678 ;
      RECT MASK 2 0.829 21.6535 1.884 21.7135 ;
      RECT MASK 2 2.422 21.78 4.189 21.84 ;
      RECT MASK 2 2.015 21.84 2.287 21.9 ;
      RECT MASK 2 5.399 21.84 11.0795 21.9 ;
      RECT MASK 2 13.865 21.882 20.669 22.082 ;
      RECT MASK 2 20.975 21.885 32.129 22.065 ;
      RECT MASK 2 5.747 22.08 13.535 22.14 ;
      RECT MASK 2 0.829 22.11 1.636 22.17 ;
      RECT MASK 2 15.02 22.315 15.628 22.375 ;
      RECT MASK 2 17.178 22.315 19.197 22.375 ;
      RECT MASK 2 1.963 22.32 3.3865 22.38 ;
      RECT MASK 2 3.659 22.32 13.229 22.38 ;
      RECT MASK 2 0.829 22.35 1.636 22.41 ;
      RECT MASK 2 18.028 22.555 18.528 22.615 ;
      RECT MASK 2 19.356 22.555 19.856 22.615 ;
      RECT MASK 2 0.829 22.59 1.636 22.65 ;
      RECT MASK 2 2.1125 22.62 3.1835 22.8 ;
      RECT MASK 2 4.486 22.62 9.608 22.8 ;
      RECT MASK 2 10.058 22.62 13.602 22.8 ;
      RECT MASK 2 20.975 22.635 32.129 22.815 ;
      RECT MASK 2 13.87 22.815 20.636 22.875 ;
      RECT MASK 2 1.963 23.04 3.3865 23.22 ;
      RECT MASK 2 3.659 23.04 9.608 23.22 ;
      RECT MASK 2 10.058 23.04 13.602 23.22 ;
      RECT MASK 2 0.829 23.07 1.636 23.13 ;
      RECT MASK 2 1.963 23.46 3.3865 23.52 ;
      RECT MASK 2 3.659 23.46 13.229 23.52 ;
      RECT MASK 2 15.1085 23.5825 20.753 23.6425 ;
      RECT MASK 2 5.747 23.7 13.535 23.76 ;
      RECT MASK 2 22.46 23.715 24.26 23.895 ;
      RECT MASK 2 15.1085 23.8225 20.753 23.8825 ;
      RECT MASK 2 5.399 23.94 11.0795 24 ;
      RECT MASK 2 13.315 23.94 13.923 24 ;
      RECT MASK 2 2.422 24 4.189 24.06 ;
      RECT MASK 2 15.1085 24.0625 20.753 24.1225 ;
      RECT MASK 2 0.872 24.08 1.536 24.12 ;
      RECT MASK 2 13.87 24.358 20.837 24.558 ;
      RECT MASK 2 2.217 24.42 13.7215 24.48 ;
      RECT MASK 2 0.832 24.44 2.078 24.48 ;
      RECT MASK 2 2.202 24.72 13.6395 24.9 ;
      RECT MASK 2 13.996 24.762 20.669 24.962 ;
      RECT MASK 2 0.832 24.77 2.073 24.81 ;
      RECT MASK 2 0.832 24.93 2.073 24.97 ;
      RECT MASK 2 0.832 25.09 2.073 25.13 ;
      RECT MASK 2 15.1085 25.1425 20.753 25.2025 ;
      RECT MASK 2 15.1085 25.3825 20.753 25.4425 ;
      RECT MASK 2 3.4385 25.424 13.524 25.604 ;
      RECT MASK 2 20.9405 25.424 32.1465 25.604 ;
      RECT MASK 2 13.87 25.6225 20.636 25.6825 ;
      RECT MASK 2 13.87 26.075 20.636 26.135 ;
    LAYER M3 SPACING 0 ;
      RECT MASK 1 0.824 0.3005 0.944 27.0595 ;
      RECT MASK 1 1.58 0.3005 1.7 27.0595 ;
      RECT MASK 1 1.958 0.3005 2.078 27.0595 ;
      RECT MASK 1 2.714 0.3005 2.834 27.0595 ;
      RECT MASK 1 3.47 0.3005 3.59 27.0595 ;
      RECT MASK 1 3.848 0.3005 3.968 27.0595 ;
      RECT MASK 1 4.604 0.3005 4.724 27.0595 ;
      RECT MASK 1 5.36 0.3005 5.48 27.0595 ;
      RECT MASK 1 5.738 0.3005 5.858 27.0595 ;
      RECT MASK 1 6.494 0.3005 6.614 27.0595 ;
      RECT MASK 1 7.25 0.3005 7.37 16.6905 ;
      RECT MASK 1 7.628 0.3005 7.748 17.099 ;
      RECT MASK 1 8.384 0.3005 8.504 18.999 ;
      RECT MASK 1 9.14 0.3005 9.26 16.6905 ;
      RECT MASK 1 9.518 0.3005 9.638 17.099 ;
      RECT MASK 1 10.274 0.3005 10.394 18.999 ;
      RECT MASK 1 11.03 0.3005 11.15 16.6905 ;
      RECT MASK 1 11.408 0.3005 11.528 17.099 ;
      RECT MASK 1 12.164 0.3005 12.284 18.999 ;
      RECT MASK 1 12.92 0.3005 13.04 16.768 ;
      RECT MASK 1 13.298 0.3005 13.418 11.2805 ;
      RECT MASK 1 14.054 0.3005 14.174 18.999 ;
      RECT MASK 1 14.81 0.3005 14.93 16.6905 ;
      RECT MASK 1 15.188 0.3005 15.308 11.2805 ;
      RECT MASK 1 15.944 0.3005 16.064 18.999 ;
      RECT MASK 1 16.7 0.3005 16.82 16.6905 ;
      RECT MASK 1 17.078 0.3005 17.198 11.2805 ;
      RECT MASK 1 17.834 0.3005 17.954 18.999 ;
      RECT MASK 1 18.59 0.3005 18.71 16.6905 ;
      RECT MASK 1 18.968 0.3005 19.088 11.2805 ;
      RECT MASK 1 19.724 0.3005 19.844 18.999 ;
      RECT MASK 1 20.48 0.3005 20.6 16.6905 ;
      RECT MASK 1 20.858 0.3005 20.978 11.2805 ;
      RECT MASK 1 21.614 0.3005 21.734 27.0595 ;
      RECT MASK 1 22.37 0.3005 22.49 27.0595 ;
      RECT MASK 1 22.748 0.3005 22.868 11.2805 ;
      RECT MASK 1 23.504 0.3005 23.624 27.0595 ;
      RECT MASK 1 24.26 0.3005 24.38 27.0595 ;
      RECT MASK 1 24.638 0.3005 24.758 11.2805 ;
      RECT MASK 1 25.394 0.3005 25.514 27.0595 ;
      RECT MASK 1 26.15 0.3005 26.27 27.0595 ;
      RECT MASK 1 26.528 0.3005 26.648 11.2805 ;
      RECT MASK 1 27.284 0.3005 27.404 27.0595 ;
      RECT MASK 1 28.04 0.3005 28.16 27.0595 ;
      RECT MASK 1 28.418 0.3005 28.538 11.2805 ;
      RECT MASK 1 29.174 0.3005 29.294 27.0595 ;
      RECT MASK 1 29.93 0.3005 30.05 27.0595 ;
      RECT MASK 1 30.308 0.3005 30.428 11.2805 ;
      RECT MASK 1 31.064 0.3005 31.184 27.0595 ;
      RECT MASK 1 31.82 0.3005 31.94 27.0595 ;
      RECT MASK 1 32.198 0.3005 32.318 27.0595 ;
      RECT MASK 1 31.435 1.075 31.495 1.37 ;
      RECT MASK 1 30.608 1.41 30.668 1.7605 ;
      RECT MASK 1 23.126 8.061 23.246 11.2805 ;
      RECT MASK 1 25.016 8.061 25.136 11.2805 ;
      RECT MASK 1 29.543 8.864 29.583 15.4565 ;
      RECT MASK 1 13.678 9.14 13.738 11.2695 ;
      RECT MASK 1 30.775 9.485 30.815 11.274 ;
      RECT MASK 1 19.346 9.5975 19.466 11.1195 ;
      RECT MASK 1 20.102 9.5975 20.222 11.1195 ;
      RECT MASK 1 21.236 9.5975 21.356 11.1195 ;
      RECT MASK 1 27.6925 11.559 27.7525 12.014 ;
      RECT MASK 1 5.1035 11.6265 5.1635 17.905 ;
      RECT MASK 1 13.298 11.7555 13.418 12.7255 ;
      RECT MASK 1 13.676 11.7555 13.796 12.7255 ;
      RECT MASK 1 15.188 11.7555 15.308 12.7255 ;
      RECT MASK 1 15.566 11.7555 15.686 12.7255 ;
      RECT MASK 1 17.078 11.7555 17.198 12.7255 ;
      RECT MASK 1 17.456 11.7555 17.576 12.7255 ;
      RECT MASK 1 18.968 11.7555 19.088 12.7255 ;
      RECT MASK 1 19.346 11.7555 19.466 12.7255 ;
      RECT MASK 1 20.858 11.7555 20.978 12.7255 ;
      RECT MASK 1 21.236 11.7555 21.356 12.7255 ;
      RECT MASK 1 22.748 11.7555 22.868 12.7255 ;
      RECT MASK 1 23.126 11.7555 23.246 12.7255 ;
      RECT MASK 1 24.638 11.7555 24.758 12.7255 ;
      RECT MASK 1 25.016 11.7555 25.136 12.7255 ;
      RECT MASK 1 26.528 11.7555 26.648 12.7255 ;
      RECT MASK 1 26.906 11.7555 27.026 12.7255 ;
      RECT MASK 1 28.418 11.7555 28.538 12.7255 ;
      RECT MASK 1 28.796 11.7555 28.916 12.7255 ;
      RECT MASK 1 30.308 11.7555 30.428 12.7255 ;
      RECT MASK 1 30.686 11.7555 30.806 12.7255 ;
      RECT MASK 1 31.442 11.7555 31.562 12.7255 ;
      RECT MASK 1 8.006 13.1145 8.126 18.999 ;
      RECT MASK 1 8.762 13.1145 8.882 18.999 ;
      RECT MASK 1 9.896 13.1145 10.016 18.9055 ;
      RECT MASK 1 10.652 13.1145 10.772 18.837 ;
      RECT MASK 1 11.786 13.1145 11.906 18.999 ;
      RECT MASK 1 12.542 13.1145 12.662 18.999 ;
      RECT MASK 1 13.676 13.1145 13.796 18.818 ;
      RECT MASK 1 15.566 13.1145 15.686 18.999 ;
      RECT MASK 1 16.322 13.1145 16.442 18.8205 ;
      RECT MASK 1 17.456 13.1145 17.576 18.999 ;
      RECT MASK 1 18.212 13.1145 18.332 18.999 ;
      RECT MASK 1 19.346 13.1145 19.466 18.8205 ;
      RECT MASK 1 13.298 13.1955 13.418 17.099 ;
      RECT MASK 1 15.188 13.1955 15.308 15.2205 ;
      RECT MASK 1 17.078 13.1955 17.198 17.099 ;
      RECT MASK 1 18.968 13.1955 19.088 17.099 ;
      RECT MASK 1 20.858 13.1955 20.978 27.0595 ;
      RECT MASK 1 22.748 13.1955 22.868 27.0595 ;
      RECT MASK 1 24.638 13.1955 24.758 27.0595 ;
      RECT MASK 1 26.528 13.1955 26.648 27.0595 ;
      RECT MASK 1 28.418 13.1955 28.538 27.0595 ;
      RECT MASK 1 14.432 13.546 14.552 18.8205 ;
      RECT MASK 1 30.308 14.0705 30.428 27.0595 ;
      RECT MASK 1 20.093 14.51 20.153 15.611 ;
      RECT MASK 1 15.179 15.3605 15.239 22.4185 ;
      RECT MASK 1 20.093 16.187 20.153 17.6005 ;
      RECT MASK 1 7.25 17.1485 7.37 18.999 ;
      RECT MASK 1 9.14 17.1485 9.26 18.999 ;
      RECT MASK 1 11.03 17.1485 11.15 18.999 ;
      RECT MASK 1 14.81 17.1485 14.93 18.999 ;
      RECT MASK 1 16.7 17.1485 16.82 18.999 ;
      RECT MASK 1 18.59 17.1485 18.71 18.999 ;
      RECT MASK 1 20.48 17.1485 20.6 18.999 ;
      RECT MASK 1 7.628 17.5465 7.748 18.999 ;
      RECT MASK 1 9.518 17.5465 9.638 18.999 ;
      RECT MASK 1 11.408 17.5465 11.528 18.837 ;
      RECT MASK 1 12.92 17.5465 13.04 18.999 ;
      RECT MASK 1 13.298 17.5465 13.418 18.818 ;
      RECT MASK 1 17.078 17.5465 17.198 18.8205 ;
      RECT MASK 1 18.968 17.5465 19.088 18.8205 ;
      RECT MASK 1 20.102 17.8585 20.222 18.8205 ;
      RECT MASK 1 19.415 18.9805 19.475 20.919 ;
      RECT MASK 1 10.643 19.0195 10.703 19.333 ;
      RECT MASK 1 14.423 19.0195 14.483 19.313 ;
      RECT MASK 1 16.313 19.0195 16.373 19.313 ;
      RECT MASK 1 20.093 19.0195 20.153 19.313 ;
      RECT MASK 1 9.965 19.154 10.025 20.799 ;
      RECT MASK 1 13.745 19.194 13.805 20.799 ;
      RECT MASK 1 7.25 19.259 7.37 27.1205 ;
      RECT MASK 1 7.628 19.259 7.748 27.1205 ;
      RECT MASK 1 8.006 19.259 8.126 20.6405 ;
      RECT MASK 1 8.384 19.259 8.504 20.6405 ;
      RECT MASK 1 8.762 19.259 8.882 20.6405 ;
      RECT MASK 1 9.14 19.259 9.26 27.1205 ;
      RECT MASK 1 9.518 19.259 9.638 27.1205 ;
      RECT MASK 1 11.03 19.259 11.15 27.1205 ;
      RECT MASK 1 11.408 19.259 11.528 27.1205 ;
      RECT MASK 1 11.786 19.259 11.906 20.6405 ;
      RECT MASK 1 12.164 19.259 12.284 20.6405 ;
      RECT MASK 1 12.542 19.259 12.662 27.1205 ;
      RECT MASK 1 12.92 19.259 13.04 27.1205 ;
      RECT MASK 1 13.298 19.259 13.418 27.1205 ;
      RECT MASK 1 14.054 19.259 14.174 21.2005 ;
      RECT MASK 1 14.81 19.259 14.93 21.2005 ;
      RECT MASK 1 15.566 19.259 15.686 21.2005 ;
      RECT MASK 1 15.944 19.259 16.064 21.2005 ;
      RECT MASK 1 16.7 19.259 16.82 21.2005 ;
      RECT MASK 1 17.078 19.259 17.198 21.2005 ;
      RECT MASK 1 17.456 19.259 17.576 21.2005 ;
      RECT MASK 1 17.834 19.259 17.954 21.2005 ;
      RECT MASK 1 18.212 19.259 18.332 21.2005 ;
      RECT MASK 1 18.59 19.259 18.71 21.2005 ;
      RECT MASK 1 18.968 19.259 19.088 21.2005 ;
      RECT MASK 1 19.724 19.259 19.844 21.2005 ;
      RECT MASK 1 20.48 19.259 20.6 27.0595 ;
      RECT MASK 1 10.274 19.4685 10.394 20.6405 ;
      RECT MASK 1 10.652 19.469 10.772 27.1205 ;
      RECT MASK 1 14.432 19.469 14.552 21.2005 ;
      RECT MASK 1 16.322 19.469 16.442 21.2005 ;
      RECT MASK 1 20.102 19.469 20.222 21.2005 ;
      RECT MASK 1 3.083 19.8405 3.143 20.525 ;
      RECT MASK 1 8.006 20.995 8.126 27.0595 ;
      RECT MASK 1 8.384 20.995 8.504 27.0595 ;
      RECT MASK 1 8.762 20.995 8.882 27.0595 ;
      RECT MASK 1 10.274 20.995 10.394 27.0595 ;
      RECT MASK 1 12.164 20.995 12.284 27.0595 ;
      RECT MASK 1 9.896 21.242 10.016 27.0595 ;
      RECT MASK 1 11.786 21.242 11.906 27.0595 ;
      RECT MASK 1 14.054 21.478 14.174 22.4205 ;
      RECT MASK 1 14.432 21.478 14.552 22.4205 ;
      RECT MASK 1 14.81 21.478 14.93 22.4205 ;
      RECT MASK 1 15.566 21.478 15.686 22.4205 ;
      RECT MASK 1 15.944 21.478 16.064 22.4205 ;
      RECT MASK 1 16.322 21.478 16.442 22.4205 ;
      RECT MASK 1 16.7 21.478 16.82 22.4205 ;
      RECT MASK 1 17.078 21.478 17.198 22.4205 ;
      RECT MASK 1 17.456 21.478 17.576 22.4205 ;
      RECT MASK 1 17.834 21.478 17.954 22.4205 ;
      RECT MASK 1 18.212 21.478 18.332 22.4205 ;
      RECT MASK 1 18.59 21.478 18.71 22.4205 ;
      RECT MASK 1 18.968 21.478 19.088 22.4205 ;
      RECT MASK 1 19.346 21.478 19.466 22.4205 ;
      RECT MASK 1 19.724 21.478 19.844 22.4205 ;
      RECT MASK 1 20.102 21.478 20.222 22.4205 ;
      RECT MASK 1 19.376 22.55 19.436 25.5675 ;
      RECT MASK 1 14.054 22.685 14.174 23.88 ;
      RECT MASK 1 14.432 22.685 14.552 23.88 ;
      RECT MASK 1 14.81 22.685 14.93 23.88 ;
      RECT MASK 1 15.188 22.685 15.308 23.88 ;
      RECT MASK 1 15.566 22.685 15.686 23.88 ;
      RECT MASK 1 15.944 22.685 16.064 23.88 ;
      RECT MASK 1 16.322 22.685 16.442 23.88 ;
      RECT MASK 1 16.7 22.685 16.82 23.88 ;
      RECT MASK 1 17.078 22.685 17.198 23.88 ;
      RECT MASK 1 17.456 22.685 17.576 23.88 ;
      RECT MASK 1 17.834 22.685 17.954 23.88 ;
      RECT MASK 1 18.212 22.685 18.332 23.88 ;
      RECT MASK 1 18.59 22.685 18.71 23.88 ;
      RECT MASK 1 18.968 22.685 19.088 23.88 ;
      RECT MASK 1 19.724 22.685 19.844 23.88 ;
      RECT MASK 1 20.102 22.685 20.222 23.88 ;
      RECT MASK 1 1.359 23.436 1.419 23.987 ;
      RECT MASK 1 14.054 24.14 14.174 25.3295 ;
      RECT MASK 1 14.432 24.14 14.552 25.3295 ;
      RECT MASK 1 14.81 24.14 14.93 25.3295 ;
      RECT MASK 1 15.188 24.14 15.308 25.3295 ;
      RECT MASK 1 15.566 24.14 15.686 25.3295 ;
      RECT MASK 1 15.944 24.14 16.064 25.3295 ;
      RECT MASK 1 16.322 24.14 16.442 25.3295 ;
      RECT MASK 1 16.7 24.14 16.82 25.3295 ;
      RECT MASK 1 17.078 24.14 17.198 25.3295 ;
      RECT MASK 1 17.456 24.14 17.576 25.3295 ;
      RECT MASK 1 17.834 24.14 17.954 25.3295 ;
      RECT MASK 1 18.212 24.14 18.332 25.3295 ;
      RECT MASK 1 18.59 24.14 18.71 25.3295 ;
      RECT MASK 1 18.968 24.14 19.088 25.3295 ;
      RECT MASK 1 19.724 24.14 19.844 25.3295 ;
      RECT MASK 1 20.102 24.14 20.222 25.3295 ;
      RECT MASK 1 14.054 25.5895 14.174 27.1205 ;
      RECT MASK 1 14.432 25.5895 14.552 27.0595 ;
      RECT MASK 1 14.81 25.5895 14.93 27.0595 ;
      RECT MASK 1 15.188 25.5895 15.308 27.0595 ;
      RECT MASK 1 15.566 25.5895 15.686 27.0595 ;
      RECT MASK 1 15.944 25.5895 16.064 27.0595 ;
      RECT MASK 1 16.322 25.5895 16.442 27.0595 ;
      RECT MASK 1 16.7 25.5895 16.82 27.0595 ;
      RECT MASK 1 17.078 25.5895 17.198 27.0595 ;
      RECT MASK 1 17.456 25.5895 17.576 27.0595 ;
      RECT MASK 1 17.834 25.5895 17.954 27.0595 ;
      RECT MASK 1 18.212 25.5895 18.332 27.0595 ;
      RECT MASK 1 18.59 25.5895 18.71 27.0595 ;
      RECT MASK 1 18.968 25.5895 19.088 27.0595 ;
      RECT MASK 1 19.724 25.5895 19.844 27.0595 ;
      RECT MASK 1 20.102 25.5895 20.222 27.0595 ;
      RECT MASK 1 19.346 25.7075 19.466 27.0595 ;
    LAYER M4 SPACING 0 ;
      RECT 0 0 32.604 27.36 ;
    LAYER M3 SPACING 0 ;
      RECT MASK 2 0.635 0.3005 0.755 27.0595 ;
      RECT MASK 2 1.013 0.3005 1.133 27.0595 ;
      RECT MASK 2 1.769 0.3005 1.889 27.0595 ;
      RECT MASK 2 2.525 0.3005 2.645 27.0595 ;
      RECT MASK 2 2.903 0.3005 3.023 27.0595 ;
      RECT MASK 2 3.659 0.3005 3.779 27.0595 ;
      RECT MASK 2 4.415 0.3005 4.535 27.0595 ;
      RECT MASK 2 4.793 0.3005 4.913 27.0595 ;
      RECT MASK 2 5.549 0.3005 5.669 27.0595 ;
      RECT MASK 2 6.305 0.3005 6.425 27.0595 ;
      RECT MASK 2 6.683 0.3005 6.803 27.0595 ;
      RECT MASK 2 7.439 0.3005 7.559 18.999 ;
      RECT MASK 2 8.195 0.3005 8.315 16.6905 ;
      RECT MASK 2 8.573 0.3005 8.693 17.099 ;
      RECT MASK 2 9.329 0.3005 9.449 18.999 ;
      RECT MASK 2 10.085 0.3005 10.205 16.6905 ;
      RECT MASK 2 10.463 0.3005 10.583 17.099 ;
      RECT MASK 2 11.219 0.3005 11.339 18.999 ;
      RECT MASK 2 11.975 0.3005 12.095 16.6905 ;
      RECT MASK 2 12.353 0.3005 12.473 11.2805 ;
      RECT MASK 2 13.109 0.3005 13.229 18.999 ;
      RECT MASK 2 13.865 0.3005 13.985 16.6905 ;
      RECT MASK 2 14.243 0.3005 14.363 11.2805 ;
      RECT MASK 2 14.999 0.3005 15.119 18.999 ;
      RECT MASK 2 15.755 0.3005 15.875 16.6905 ;
      RECT MASK 2 16.133 0.3005 16.253 11.2805 ;
      RECT MASK 2 16.889 0.3005 17.009 18.999 ;
      RECT MASK 2 17.645 0.3005 17.765 16.6905 ;
      RECT MASK 2 18.023 0.3005 18.143 11.2805 ;
      RECT MASK 2 18.779 0.3005 18.899 18.999 ;
      RECT MASK 2 19.535 0.3005 19.655 16.6905 ;
      RECT MASK 2 19.913 0.3005 20.033 11.2805 ;
      RECT MASK 2 20.669 0.3005 20.789 27.0595 ;
      RECT MASK 2 21.425 0.3005 21.545 27.0595 ;
      RECT MASK 2 21.803 0.3005 21.923 11.2805 ;
      RECT MASK 2 22.559 0.3005 22.679 27.0595 ;
      RECT MASK 2 23.315 0.3005 23.435 27.0595 ;
      RECT MASK 2 23.693 0.3005 23.813 11.2805 ;
      RECT MASK 2 24.449 0.3005 24.569 27.0595 ;
      RECT MASK 2 25.205 0.3005 25.325 27.0595 ;
      RECT MASK 2 25.583 0.3005 25.703 11.2805 ;
      RECT MASK 2 26.339 0.3005 26.459 27.0595 ;
      RECT MASK 2 27.095 0.3005 27.215 27.0595 ;
      RECT MASK 2 27.473 0.3005 27.593 11.2805 ;
      RECT MASK 2 28.229 0.3005 28.349 27.0595 ;
      RECT MASK 2 28.985 0.3005 29.105 27.0595 ;
      RECT MASK 2 29.363 0.3005 29.483 11.2805 ;
      RECT MASK 2 30.119 0.3005 30.239 27.0595 ;
      RECT MASK 2 30.875 0.3005 30.995 27.0595 ;
      RECT MASK 2 31.253 0.3005 31.373 11.2805 ;
      RECT MASK 2 32.009 0.3005 32.129 27.0595 ;
      RECT MASK 2 29.81 0.3945 29.87 1.2525 ;
      RECT MASK 2 31.7 0.957 31.76 1.25 ;
      RECT MASK 2 22.181 8.061 22.301 11.2805 ;
      RECT MASK 2 24.071 8.061 24.191 11.2805 ;
      RECT MASK 2 25.961 8.061 26.081 11.2805 ;
      RECT MASK 2 17.267 9.14 17.327 9.58 ;
      RECT MASK 2 30.488 9.245 30.528 13.1655 ;
      RECT MASK 2 12.682 9.26 12.742 11.2695 ;
      RECT MASK 2 18.401 9.5975 18.521 11.1195 ;
      RECT MASK 2 27.851 9.5975 27.971 11.1195 ;
      RECT MASK 2 31.631 9.5975 31.751 11.1195 ;
      RECT MASK 2 29.83 9.605 29.87 11.3675 ;
      RECT MASK 2 14.508 11.375 14.568 13.212 ;
      RECT MASK 2 31.7 11.375 31.76 11.8625 ;
      RECT MASK 2 13.512 11.4635 13.572 13.345 ;
      RECT MASK 2 12.353 11.7555 12.473 12.7255 ;
      RECT MASK 2 12.731 11.7555 12.851 12.7255 ;
      RECT MASK 2 14.243 11.7555 14.363 12.7255 ;
      RECT MASK 2 16.133 11.7555 16.253 12.7255 ;
      RECT MASK 2 16.511 11.7555 16.631 12.7255 ;
      RECT MASK 2 18.023 11.7555 18.143 12.7255 ;
      RECT MASK 2 18.401 11.7555 18.521 12.7255 ;
      RECT MASK 2 19.913 11.7555 20.033 12.7255 ;
      RECT MASK 2 20.291 11.7555 20.411 12.7255 ;
      RECT MASK 2 21.803 11.7555 21.923 12.7255 ;
      RECT MASK 2 22.181 11.7555 22.301 12.7255 ;
      RECT MASK 2 23.693 11.7555 23.813 12.7255 ;
      RECT MASK 2 24.071 11.7555 24.191 12.7255 ;
      RECT MASK 2 25.583 11.7555 25.703 12.7255 ;
      RECT MASK 2 25.961 11.7555 26.081 12.7255 ;
      RECT MASK 2 27.473 11.7555 27.593 12.7255 ;
      RECT MASK 2 27.851 11.7555 27.971 12.7255 ;
      RECT MASK 2 29.363 11.7555 29.483 12.7255 ;
      RECT MASK 2 29.741 11.7555 29.861 12.7255 ;
      RECT MASK 2 31.253 11.7555 31.373 12.7255 ;
      RECT MASK 2 7.817 13.1145 7.937 18.999 ;
      RECT MASK 2 8.951 13.1145 9.071 18.999 ;
      RECT MASK 2 9.707 13.1145 9.827 18.999 ;
      RECT MASK 2 10.841 13.1145 10.961 18.837 ;
      RECT MASK 2 11.597 13.1145 11.717 18.837 ;
      RECT MASK 2 15.377 13.1145 15.497 18.85 ;
      RECT MASK 2 16.511 13.1145 16.631 18.8205 ;
      RECT MASK 2 17.267 13.1145 17.387 18.8205 ;
      RECT MASK 2 18.401 13.1145 18.521 18.8205 ;
      RECT MASK 2 19.157 13.1145 19.277 18.8205 ;
      RECT MASK 2 12.353 13.1955 12.473 17.099 ;
      RECT MASK 2 14.243 13.1955 14.363 17.099 ;
      RECT MASK 2 16.133 13.1955 16.253 17.099 ;
      RECT MASK 2 18.023 13.1955 18.143 17.099 ;
      RECT MASK 2 19.913 13.1955 20.033 17.104 ;
      RECT MASK 2 20.291 13.1955 20.411 17.099 ;
      RECT MASK 2 21.803 13.1955 21.923 27.0595 ;
      RECT MASK 2 23.693 13.1955 23.813 27.0595 ;
      RECT MASK 2 25.583 13.1955 25.703 27.0595 ;
      RECT MASK 2 27.473 13.1955 27.593 27.0595 ;
      RECT MASK 2 29.363 13.1955 29.483 27.0595 ;
      RECT MASK 2 31.253 13.1955 31.373 27.0595 ;
      RECT MASK 2 13.487 13.546 13.607 18.818 ;
      RECT MASK 2 14.621 13.546 14.741 18.999 ;
      RECT MASK 2 12.8 15.3575 12.86 16.45 ;
      RECT MASK 2 12.731 16.7215 12.851 18.818 ;
      RECT MASK 2 8.195 17.1485 8.315 18.999 ;
      RECT MASK 2 10.085 17.1485 10.205 18.999 ;
      RECT MASK 2 11.975 17.1485 12.095 18.999 ;
      RECT MASK 2 13.865 17.1485 13.985 18.999 ;
      RECT MASK 2 15.755 17.1485 15.875 18.85 ;
      RECT MASK 2 17.645 17.1485 17.765 18.999 ;
      RECT MASK 2 19.535 17.1485 19.655 18.999 ;
      RECT MASK 2 8.573 17.5465 8.693 18.999 ;
      RECT MASK 2 10.463 17.5465 10.583 18.837 ;
      RECT MASK 2 12.353 17.5465 12.473 18.999 ;
      RECT MASK 2 14.243 17.5465 14.363 18.8205 ;
      RECT MASK 2 16.133 17.5465 16.253 18.8205 ;
      RECT MASK 2 18.023 17.5465 18.143 18.999 ;
      RECT MASK 2 19.913 17.5465 20.033 18.8205 ;
      RECT MASK 2 20.291 17.5465 20.411 18.999 ;
      RECT MASK 2 15.437 18.9805 15.497 20.919 ;
      RECT MASK 2 10.853 18.997 10.913 20.919 ;
      RECT MASK 2 11.588 19.0195 11.648 19.333 ;
      RECT MASK 2 13.478 19.0195 13.538 19.333 ;
      RECT MASK 2 17.258 19.0195 17.318 19.313 ;
      RECT MASK 2 19.148 19.0195 19.208 19.313 ;
      RECT MASK 2 18.47 19.194 18.53 20.799 ;
      RECT MASK 2 7.439 19.259 7.559 20.6405 ;
      RECT MASK 2 7.817 19.259 7.937 20.6405 ;
      RECT MASK 2 8.195 19.259 8.315 27.1205 ;
      RECT MASK 2 8.573 19.259 8.693 27.1205 ;
      RECT MASK 2 8.951 19.259 9.071 20.6405 ;
      RECT MASK 2 9.329 19.259 9.449 20.6405 ;
      RECT MASK 2 9.707 19.259 9.827 20.6405 ;
      RECT MASK 2 10.085 19.259 10.205 27.1205 ;
      RECT MASK 2 10.463 19.259 10.583 27.1205 ;
      RECT MASK 2 11.219 19.259 11.339 20.6405 ;
      RECT MASK 2 11.975 19.259 12.095 27.1205 ;
      RECT MASK 2 12.353 19.259 12.473 27.1205 ;
      RECT MASK 2 12.731 19.259 12.851 20.6405 ;
      RECT MASK 2 13.109 19.259 13.229 20.6405 ;
      RECT MASK 2 13.865 19.259 13.985 21.2005 ;
      RECT MASK 2 14.243 19.259 14.363 21.2005 ;
      RECT MASK 2 14.621 19.259 14.741 21.2005 ;
      RECT MASK 2 14.999 19.259 15.119 21.2005 ;
      RECT MASK 2 15.755 19.259 15.875 21.2005 ;
      RECT MASK 2 16.133 19.259 16.253 21.2005 ;
      RECT MASK 2 16.511 19.259 16.631 21.2005 ;
      RECT MASK 2 16.889 19.259 17.009 21.2005 ;
      RECT MASK 2 17.645 19.259 17.765 21.2005 ;
      RECT MASK 2 18.023 19.259 18.143 21.2005 ;
      RECT MASK 2 18.779 19.259 18.899 21.2005 ;
      RECT MASK 2 19.535 19.259 19.655 21.2005 ;
      RECT MASK 2 19.913 19.259 20.033 21.2005 ;
      RECT MASK 2 20.291 19.259 20.411 21.2005 ;
      RECT MASK 2 11.597 19.469 11.717 27.1205 ;
      RECT MASK 2 13.487 19.469 13.607 27.1205 ;
      RECT MASK 2 17.267 19.469 17.387 21.2005 ;
      RECT MASK 2 19.157 19.469 19.277 21.2005 ;
      RECT MASK 2 7.439 20.995 7.559 27.0595 ;
      RECT MASK 2 7.817 20.995 7.937 27.0595 ;
      RECT MASK 2 8.951 20.995 9.071 27.0595 ;
      RECT MASK 2 9.329 20.995 9.449 27.0595 ;
      RECT MASK 2 9.707 20.995 9.827 27.0595 ;
      RECT MASK 2 11.219 20.995 11.339 27.0595 ;
      RECT MASK 2 13.109 20.995 13.229 27.0595 ;
      RECT MASK 2 10.841 21.242 10.961 27.0595 ;
      RECT MASK 2 12.731 21.242 12.851 27.0595 ;
      RECT MASK 2 13.865 21.478 13.985 22.4205 ;
      RECT MASK 2 14.243 21.478 14.363 22.4205 ;
      RECT MASK 2 14.621 21.478 14.741 22.4205 ;
      RECT MASK 2 14.999 21.478 15.119 22.4205 ;
      RECT MASK 2 15.377 21.478 15.497 22.4205 ;
      RECT MASK 2 15.755 21.478 15.875 22.4205 ;
      RECT MASK 2 16.133 21.478 16.253 22.4205 ;
      RECT MASK 2 16.511 21.478 16.631 22.4205 ;
      RECT MASK 2 16.889 21.478 17.009 22.4205 ;
      RECT MASK 2 17.267 21.478 17.387 22.4205 ;
      RECT MASK 2 17.645 21.478 17.765 22.4205 ;
      RECT MASK 2 18.023 21.478 18.143 22.4205 ;
      RECT MASK 2 18.401 21.478 18.521 22.4205 ;
      RECT MASK 2 18.779 21.478 18.899 22.4205 ;
      RECT MASK 2 19.157 21.478 19.277 22.4205 ;
      RECT MASK 2 19.535 21.478 19.655 22.4205 ;
      RECT MASK 2 19.913 21.478 20.033 22.4205 ;
      RECT MASK 2 20.291 21.478 20.411 22.4205 ;
      RECT MASK 2 2.202 21.8225 2.262 22.6435 ;
      RECT MASK 2 18.431 22.55 18.491 25.4475 ;
      RECT MASK 2 13.865 22.685 13.985 23.88 ;
      RECT MASK 2 14.243 22.685 14.363 23.88 ;
      RECT MASK 2 14.621 22.685 14.741 23.88 ;
      RECT MASK 2 14.999 22.685 15.119 23.88 ;
      RECT MASK 2 15.377 22.685 15.497 23.88 ;
      RECT MASK 2 15.755 22.685 15.875 23.88 ;
      RECT MASK 2 16.133 22.685 16.253 23.88 ;
      RECT MASK 2 16.511 22.685 16.631 23.88 ;
      RECT MASK 2 16.889 22.685 17.009 23.88 ;
      RECT MASK 2 17.267 22.685 17.387 23.4325 ;
      RECT MASK 2 17.645 22.685 17.765 23.88 ;
      RECT MASK 2 18.023 22.685 18.143 23.88 ;
      RECT MASK 2 18.779 22.685 18.899 23.88 ;
      RECT MASK 2 19.157 22.685 19.277 23.88 ;
      RECT MASK 2 19.535 22.685 19.655 23.88 ;
      RECT MASK 2 19.913 22.685 20.033 23.88 ;
      RECT MASK 2 20.291 22.685 20.411 23.88 ;
      RECT MASK 2 17.258 23.5725 17.318 24.2405 ;
      RECT MASK 2 13.865 24.14 13.985 25.3295 ;
      RECT MASK 2 14.243 24.14 14.363 25.3295 ;
      RECT MASK 2 14.621 24.14 14.741 25.3295 ;
      RECT MASK 2 14.999 24.14 15.119 25.3295 ;
      RECT MASK 2 15.377 24.14 15.497 25.3295 ;
      RECT MASK 2 15.755 24.14 15.875 25.3295 ;
      RECT MASK 2 16.133 24.14 16.253 25.3295 ;
      RECT MASK 2 16.511 24.14 16.631 25.3295 ;
      RECT MASK 2 16.889 24.14 17.009 25.3295 ;
      RECT MASK 2 17.645 24.14 17.765 25.3295 ;
      RECT MASK 2 18.023 24.14 18.143 25.3295 ;
      RECT MASK 2 18.779 24.14 18.899 25.3295 ;
      RECT MASK 2 19.157 24.14 19.277 25.3295 ;
      RECT MASK 2 19.535 24.14 19.655 25.3295 ;
      RECT MASK 2 19.913 24.14 20.033 25.3295 ;
      RECT MASK 2 20.291 24.14 20.411 25.3295 ;
      RECT MASK 2 17.267 24.3805 17.387 25.3295 ;
      RECT MASK 2 13.865 25.5895 13.985 27.1205 ;
      RECT MASK 2 14.243 25.5895 14.363 27.0595 ;
      RECT MASK 2 14.621 25.5895 14.741 27.0595 ;
      RECT MASK 2 14.999 25.5895 15.119 27.0595 ;
      RECT MASK 2 15.377 25.5895 15.497 27.0595 ;
      RECT MASK 2 15.755 25.5895 15.875 27.0595 ;
      RECT MASK 2 16.133 25.5895 16.253 27.0595 ;
      RECT MASK 2 16.511 25.5895 16.631 27.0595 ;
      RECT MASK 2 16.889 25.5895 17.009 27.0595 ;
      RECT MASK 2 17.267 25.5895 17.387 27.0595 ;
      RECT MASK 2 17.645 25.5895 17.765 27.0595 ;
      RECT MASK 2 18.023 25.5895 18.143 27.0595 ;
      RECT MASK 2 18.401 25.5895 18.521 27.0595 ;
      RECT MASK 2 18.779 25.5895 18.899 27.0595 ;
      RECT MASK 2 19.913 25.5895 20.033 27.0595 ;
      RECT MASK 2 20.291 25.5895 20.411 27.0595 ;
      RECT MASK 2 19.157 25.7075 19.277 27.0595 ;
      RECT MASK 2 19.535 25.7075 19.655 27.0595 ;
    LAYER M4 SPACING 0 ;
      RECT MASK 2 7.2315 22.7205 20.448 22.8005 ;
    LAYER M5 SPACING 0 ;
      POLYGON 27.8275 0 27.8275 0.08 27.9075 0.08 27.9075 0 29.8905 0 29.8905 0.08 29.9705 0.08 29.9705 0 32.604 0 32.604 27.36 32.1935 27.36 32.1935 27.28 32.1135 27.28 32.1135 27.36 31.6125 27.36 31.6125 27.28 31.5325 27.28 31.5325 27.36 31.4525 27.36 31.4525 27.28 31.3725 27.28 31.3725 27.36 30.8715 27.36 30.8715 27.28 30.7915 27.28 30.7915 27.36 21.0785 27.36 21.0785 27.28 20.9985 27.28 20.9985 27.36 20.4975 27.36 20.4975 27.28 20.4175 27.28 20.4175 27.36 1.0715 27.36 1.0715 27.28 0.9915 27.28 0.9915 27.36 0.4905 27.36 0.4905 27.28 0.4105 27.28 0.4105 27.36 0 27.36 0 0 ;
      RECT MASK 1 10.274 0.186 10.474 27.1805 ;
      RECT MASK 1 11.756 0.186 11.956 16.0455 ;
      RECT MASK 1 13.238 0.186 13.438 19.016 ;
      RECT MASK 1 14.72 0.186 14.92 27.1805 ;
      RECT MASK 1 16.202 0.186 16.402 16.0455 ;
      RECT MASK 1 17.684 0.186 17.884 27.1805 ;
      RECT MASK 1 19.166 0.186 19.366 16.0455 ;
      RECT MASK 1 20.648 0.186 20.848 0.3795 ;
      RECT MASK 1 22.13 0.186 22.33 0.3795 ;
      RECT MASK 1 23.612 0.186 23.812 0.3795 ;
      RECT MASK 1 25.094 0.186 25.294 0.3795 ;
      RECT MASK 1 26.576 0.186 26.776 0.3795 ;
      RECT MASK 1 28.058 0.186 28.258 0.3795 ;
      RECT MASK 1 29.54 0.186 29.74 0.3795 ;
      RECT MASK 1 31.022 0.186 31.222 0.3795 ;
      RECT MASK 1 11.015 0.4085 11.215 27.1805 ;
      RECT MASK 1 19.166 16.31 19.366 23.8775 ;
      RECT MASK 1 11.756 16.3555 11.956 22.5255 ;
      RECT MASK 1 16.202 16.3555 16.402 22.5255 ;
      RECT MASK 1 13.238 19.252 13.438 27.1805 ;
      RECT MASK 1 0.9915 22.5605 1.0715 23.2205 ;
      RECT MASK 1 11.756 22.7205 11.956 27.1805 ;
      RECT MASK 1 16.202 22.7205 16.402 27.1805 ;
      RECT MASK 1 19.166 24.2755 19.366 27.1805 ;
      RECT MASK 1 20.648 26.987 20.848 27.1805 ;
      RECT MASK 1 22.13 26.987 22.33 27.1805 ;
      RECT MASK 1 23.612 26.987 23.812 27.1805 ;
      RECT MASK 1 24.353 26.987 24.553 27.1805 ;
      RECT MASK 1 25.094 26.987 25.294 27.1805 ;
      RECT MASK 1 26.576 26.987 26.776 27.1805 ;
      RECT MASK 1 28.058 26.987 28.258 27.1805 ;
      RECT MASK 1 29.54 26.987 29.74 27.1805 ;
      RECT MASK 1 30.281 26.987 30.481 27.1805 ;
      RECT MASK 1 31.022 26.987 31.222 27.1805 ;
    LAYER M6 SPACING 0 ;
      POLYGON 32.604 0 32.604 24.3005 32.244 24.3005 32.244 24.6605 32.604 24.6605 32.604 27.36 0 27.36 0 23.2205 0.36 23.2205 0.36 22.8605 0 22.8605 0 0 ;
      RECT MASK 1 0.3 17.1005 32.304 17.4605 ;
      RECT MASK 1 0.3 18.5405 32.304 18.9005 ;
      RECT MASK 1 0.3 19.9805 32.304 20.3405 ;
      RECT MASK 1 0.3 21.4205 32.304 21.7805 ;
      RECT MASK 1 0.3 22.1405 32.304 22.5005 ;
      RECT MASK 1 1.382 22.8605 32.304 23.2205 ;
    LAYER M7 SPACING 0 ;
      POLYGON 14.877 0 14.877 0.45 15.327 0.45 15.327 0 32.604 0 32.604 27.36 0 27.36 0 0 ;
    LAYER M8 SPACING 0 ;
      POLYGON 0 0 0 27.36 32.604 27.36 32.604 27.1405 0.3 27.1405 0.3 26.6905 32.304 26.6905 32.304 27.1405 32.604 27.1405 32.604 26.3405 0.3 26.3405 0.3 25.8905 32.304 25.8905 32.304 26.3405 32.604 26.3405 32.604 25.5405 0.3 25.5405 0.3 25.0905 32.314 25.0905 32.314 25.5405 32.604 25.5405 32.604 24.7305 0.3 24.7305 0.3 24.2305 24.314 24.2305 24.314 24.7305 24.614 24.7305 24.614 24.2305 32.314 24.2305 32.314 24.7305 32.604 24.7305 32.604 23.8705 0.3 23.8705 0.3 23.4205 32.304 23.4205 32.304 23.8705 32.604 23.8705 32.604 23.0705 0.3 23.0705 0.3 22.6205 32.304 22.6205 32.304 23.0705 32.604 23.0705 32.604 22.2605 0.3 22.2605 0.3 21.6605 32.304 21.6605 32.304 22.2605 32.604 22.2605 32.604 21.3005 0.3 21.3005 0.3 20.8505 32.304 20.8505 32.304 21.3005 32.604 21.3005 32.604 20.5005 0.3 20.5005 0.3 20.0505 32.304 20.0505 32.304 20.5005 32.604 20.5005 32.604 19.6905 0.3 19.6905 0.3 19.1905 10.1235 19.1905 10.1235 19.6905 10.555 19.6905 10.555 19.1905 20.1615 19.1905 20.1615 19.6905 20.497 19.6905 20.497 19.1905 32.304 19.1905 32.304 19.6905 32.604 19.6905 32.604 18.8305 0.3 18.8305 0.3 18.3805 32.304 18.3805 32.304 18.8305 32.604 18.8305 32.604 18.0305 0.3 18.0305 0.3 17.5805 32.304 17.5805 32.304 18.0305 32.604 18.0305 32.604 17.2305 0.3 17.2305 0.3 16.7805 32.304 16.7805 32.304 17.2305 32.604 17.2305 32.604 16.4305 0.3 16.4305 0.3 15.9805 32.304 15.9805 32.304 16.4305 32.604 16.4305 32.604 15.6305 0.3 15.6305 0.3 15.1805 32.304 15.1805 32.304 15.6305 32.604 15.6305 32.604 14.8305 0.3 14.8305 0.3 14.3805 32.304 14.3805 32.304 14.8305 32.604 14.8305 32.604 14.0305 0.3 14.0305 0.3 13.5805 32.304 13.5805 32.304 14.0305 32.604 14.0305 32.604 13.2305 0.3 13.2305 0.3 12.7805 32.304 12.7805 32.304 13.2305 32.604 13.2305 32.604 12.4305 0.3 12.4305 0.3 11.9805 32.304 11.9805 32.304 12.4305 32.604 12.4305 32.604 11.6305 0.3 11.6305 0.3 11.1805 32.304 11.1805 32.304 11.6305 32.604 11.6305 32.604 10.8305 0.3 10.8305 0.3 10.3805 32.304 10.3805 32.304 10.8305 32.604 10.8305 32.604 10.0305 0.3 10.0305 0.3 9.5805 32.304 9.5805 32.304 10.0305 32.604 10.0305 32.604 9.2305 0.3 9.2305 0.3 8.7805 32.304 8.7805 32.304 9.2305 32.604 9.2305 32.604 8.4305 0.3 8.4305 0.3 7.9805 32.304 7.9805 32.304 8.4305 32.604 8.4305 32.604 7.6305 0.3 7.6305 0.3 7.1805 32.304 7.1805 32.304 7.6305 32.604 7.6305 32.604 6.8305 0.3 6.8305 0.3 6.3805 32.304 6.3805 32.304 6.8305 32.604 6.8305 32.604 6.0305 0.3 6.0305 0.3 5.5805 32.304 5.5805 32.304 6.0305 32.604 6.0305 32.604 5.2305 0.3 5.2305 0.3 4.7805 32.304 4.7805 32.304 5.2305 32.604 5.2305 32.604 4.4305 0.3 4.4305 0.3 3.9805 32.304 3.9805 32.304 4.4305 32.604 4.4305 32.604 3.6305 0.3 3.6305 0.3 3.1805 32.304 3.1805 32.304 3.6305 32.604 3.6305 32.604 2.8305 0.3 2.8305 0.3 2.3805 32.304 2.3805 32.304 2.8305 32.604 2.8305 32.604 2.0305 0.3 2.0305 0.3 1.5805 32.304 1.5805 32.304 2.0305 32.604 2.0305 32.604 1.2305 0.3 1.2305 0.3 0.7805 32.304 0.7805 32.304 1.2305 32.604 1.2305 32.604 0 ;
    LAYER M0 SPACING 0 ;
      RECT 0 0 32.604 27.36 ;
      RECT MASK 1 0.662 0.73 28.157 0.77 ;
      RECT MASK 1 29.121 0.88 31.871 0.92 ;
      RECT MASK 1 0.838 1.0235 0.918 9.7165 ;
      RECT MASK 1 28.062 1.0235 28.142 9.7165 ;
      RECT MASK 1 29.239 1.22 29.761 1.26 ;
      RECT MASK 1 29.903 1.22 30.425 1.26 ;
      RECT MASK 1 30.567 1.22 31.089 1.26 ;
      RECT MASK 1 31.231 1.22 31.753 1.26 ;
      RECT MASK 1 29.28 1.38 29.7105 1.42 ;
      RECT MASK 1 29.944 1.38 30.3745 1.42 ;
      RECT MASK 1 30.608 1.38 31.0385 1.42 ;
      RECT MASK 1 31.3 1.38 31.684 1.42 ;
      RECT MASK 1 1.632 1.449 2.836 1.589 ;
      RECT MASK 1 3.164 1.449 4.368 1.589 ;
      RECT MASK 1 4.696 1.449 5.9 1.589 ;
      RECT MASK 1 6.228 1.449 7.432 1.589 ;
      RECT MASK 1 7.76 1.449 8.964 1.589 ;
      RECT MASK 1 9.292 1.449 10.496 1.589 ;
      RECT MASK 1 10.824 1.449 12.028 1.589 ;
      RECT MASK 1 12.356 1.449 13.56 1.589 ;
      RECT MASK 1 13.888 1.449 15.092 1.589 ;
      RECT MASK 1 15.42 1.449 16.624 1.589 ;
      RECT MASK 1 16.952 1.449 18.156 1.589 ;
      RECT MASK 1 18.484 1.449 19.688 1.589 ;
      RECT MASK 1 20.016 1.449 21.22 1.589 ;
      RECT MASK 1 21.548 1.449 22.752 1.589 ;
      RECT MASK 1 23.08 1.449 24.284 1.589 ;
      RECT MASK 1 24.612 1.449 25.816 1.589 ;
      RECT MASK 1 26.144 1.449 27.348 1.589 ;
      RECT MASK 1 29.239 1.54 29.6575 1.58 ;
      RECT MASK 1 29.903 1.54 30.3215 1.58 ;
      RECT MASK 1 30.567 1.54 30.9855 1.58 ;
      RECT MASK 1 31.231 1.54 31.6495 1.58 ;
      RECT MASK 1 29.28 1.815 29.7105 1.855 ;
      RECT MASK 1 29.944 1.815 30.3745 1.855 ;
      RECT MASK 1 30.608 1.815 31.0385 1.855 ;
      RECT MASK 1 31.3 1.815 31.684 1.855 ;
      RECT MASK 1 29.2365 1.975 29.7675 2.015 ;
      RECT MASK 1 29.9005 1.975 30.4315 2.015 ;
      RECT MASK 1 30.5645 1.975 31.0955 2.015 ;
      RECT MASK 1 31.2285 1.975 31.7595 2.015 ;
      RECT MASK 1 29.121 2.35 31.871 2.39 ;
      RECT MASK 1 29.121 2.77 31.871 2.81 ;
      RECT MASK 1 29.249 3.33 29.429 3.39 ;
      RECT MASK 1 29.571 3.33 29.751 3.39 ;
      RECT MASK 1 29.913 3.33 30.093 3.39 ;
      RECT MASK 1 30.235 3.33 30.415 3.39 ;
      RECT MASK 1 30.577 3.33 30.757 3.39 ;
      RECT MASK 1 30.899 3.33 31.079 3.39 ;
      RECT MASK 1 31.241 3.33 31.421 3.39 ;
      RECT MASK 1 31.563 3.33 31.743 3.39 ;
      RECT MASK 1 29.249 3.57 29.429 3.63 ;
      RECT MASK 1 29.571 3.57 29.751 3.63 ;
      RECT MASK 1 29.913 3.57 30.093 3.63 ;
      RECT MASK 1 30.235 3.57 30.415 3.63 ;
      RECT MASK 1 30.577 3.57 30.757 3.63 ;
      RECT MASK 1 30.899 3.57 31.079 3.63 ;
      RECT MASK 1 31.241 3.57 31.421 3.63 ;
      RECT MASK 1 31.563 3.57 31.743 3.63 ;
      RECT MASK 1 29.028 3.84 29.208 3.9 ;
      RECT MASK 1 29.538 3.84 29.794 3.9 ;
      RECT MASK 1 30.202 3.84 30.458 3.9 ;
      RECT MASK 1 30.866 3.84 31.122 3.9 ;
      RECT MASK 1 31.53 3.84 31.786 3.9 ;
      RECT MASK 1 29.028 4.26 29.208 4.32 ;
      RECT MASK 1 29.538 4.26 29.794 4.32 ;
      RECT MASK 1 30.202 4.26 30.458 4.32 ;
      RECT MASK 1 30.866 4.26 31.122 4.32 ;
      RECT MASK 1 31.53 4.26 31.786 4.32 ;
      RECT MASK 1 29.249 4.53 29.429 4.59 ;
      RECT MASK 1 29.571 4.53 29.751 4.59 ;
      RECT MASK 1 29.913 4.53 30.093 4.59 ;
      RECT MASK 1 30.235 4.53 30.415 4.59 ;
      RECT MASK 1 30.577 4.53 30.757 4.59 ;
      RECT MASK 1 30.899 4.53 31.079 4.59 ;
      RECT MASK 1 31.241 4.53 31.421 4.59 ;
      RECT MASK 1 31.563 4.53 31.743 4.59 ;
      RECT MASK 1 29.249 4.77 29.429 4.83 ;
      RECT MASK 1 29.571 4.77 29.751 4.83 ;
      RECT MASK 1 29.913 4.77 30.093 4.83 ;
      RECT MASK 1 30.235 4.77 30.415 4.83 ;
      RECT MASK 1 30.577 4.77 30.757 4.83 ;
      RECT MASK 1 30.899 4.77 31.079 4.83 ;
      RECT MASK 1 31.241 4.77 31.421 4.83 ;
      RECT MASK 1 31.563 4.77 31.743 4.83 ;
      RECT MASK 1 1.632 5.089 2.07 5.699 ;
      RECT MASK 1 2.398 5.089 2.836 5.699 ;
      RECT MASK 1 3.164 5.089 3.602 5.699 ;
      RECT MASK 1 3.93 5.089 4.368 5.699 ;
      RECT MASK 1 4.696 5.089 5.134 5.699 ;
      RECT MASK 1 5.462 5.089 5.9 5.699 ;
      RECT MASK 1 6.228 5.089 6.666 5.699 ;
      RECT MASK 1 6.994 5.089 7.432 5.699 ;
      RECT MASK 1 7.76 5.089 8.198 5.699 ;
      RECT MASK 1 8.526 5.089 8.964 5.699 ;
      RECT MASK 1 9.292 5.089 9.73 5.699 ;
      RECT MASK 1 10.058 5.089 10.496 5.699 ;
      RECT MASK 1 10.824 5.089 11.262 5.699 ;
      RECT MASK 1 11.59 5.089 12.028 5.699 ;
      RECT MASK 1 12.356 5.089 12.794 5.699 ;
      RECT MASK 1 13.122 5.089 13.56 5.699 ;
      RECT MASK 1 13.888 5.089 14.326 5.699 ;
      RECT MASK 1 14.654 5.089 15.092 5.699 ;
      RECT MASK 1 15.42 5.089 15.858 5.699 ;
      RECT MASK 1 16.186 5.089 16.624 5.699 ;
      RECT MASK 1 16.952 5.089 17.39 5.699 ;
      RECT MASK 1 17.718 5.089 18.156 5.699 ;
      RECT MASK 1 18.484 5.089 18.922 5.699 ;
      RECT MASK 1 19.25 5.089 19.688 5.699 ;
      RECT MASK 1 20.016 5.089 20.454 5.699 ;
      RECT MASK 1 20.782 5.089 21.22 5.699 ;
      RECT MASK 1 21.548 5.089 21.986 5.699 ;
      RECT MASK 1 22.314 5.089 22.752 5.699 ;
      RECT MASK 1 23.08 5.089 23.518 5.699 ;
      RECT MASK 1 23.846 5.089 24.284 5.699 ;
      RECT MASK 1 24.612 5.089 25.05 5.699 ;
      RECT MASK 1 25.378 5.089 25.816 5.699 ;
      RECT MASK 1 26.144 5.089 26.582 5.699 ;
      RECT MASK 1 26.91 5.089 27.348 5.699 ;
      RECT MASK 1 29.128 5.25 31.886 5.31 ;
      RECT MASK 1 29.249 5.49 29.429 5.55 ;
      RECT MASK 1 29.571 5.49 29.751 5.55 ;
      RECT MASK 1 29.913 5.49 30.093 5.55 ;
      RECT MASK 1 30.235 5.49 30.415 5.55 ;
      RECT MASK 1 30.577 5.49 30.757 5.55 ;
      RECT MASK 1 30.899 5.49 31.079 5.55 ;
      RECT MASK 1 31.241 5.49 31.421 5.55 ;
      RECT MASK 1 31.563 5.49 31.743 5.55 ;
      RECT MASK 1 29.128 5.73 31.886 5.79 ;
      RECT MASK 1 29.121 6.19 31.871 6.23 ;
      RECT MASK 1 29.121 6.61 31.871 6.65 ;
      RECT MASK 1 29.131 6.93 29.311 6.99 ;
      RECT MASK 1 29.431 6.93 29.651 6.99 ;
      RECT MASK 1 29.795 6.93 29.975 6.99 ;
      RECT MASK 1 30.095 6.93 30.315 6.99 ;
      RECT MASK 1 30.459 6.93 30.639 6.99 ;
      RECT MASK 1 30.759 6.93 30.979 6.99 ;
      RECT MASK 1 31.123 6.93 31.303 6.99 ;
      RECT MASK 1 31.423 6.93 31.643 6.99 ;
      RECT MASK 1 29.372 7.17 29.552 7.23 ;
      RECT MASK 1 29.692 7.17 29.872 7.23 ;
      RECT MASK 1 30.036 7.17 30.216 7.23 ;
      RECT MASK 1 30.356 7.17 30.536 7.23 ;
      RECT MASK 1 30.7 7.17 30.88 7.23 ;
      RECT MASK 1 31.02 7.17 31.2 7.23 ;
      RECT MASK 1 31.364 7.17 31.544 7.23 ;
      RECT MASK 1 31.684 7.17 31.864 7.23 ;
      RECT MASK 1 29.349 7.41 29.529 7.47 ;
      RECT MASK 1 29.692 7.41 29.872 7.47 ;
      RECT MASK 1 30.013 7.41 30.193 7.47 ;
      RECT MASK 1 30.356 7.41 30.536 7.47 ;
      RECT MASK 1 30.677 7.41 30.857 7.47 ;
      RECT MASK 1 31.02 7.41 31.2 7.47 ;
      RECT MASK 1 31.341 7.41 31.521 7.47 ;
      RECT MASK 1 31.684 7.41 31.864 7.47 ;
      RECT MASK 1 29.128 7.65 29.308 7.71 ;
      RECT MASK 1 29.448 7.65 29.628 7.71 ;
      RECT MASK 1 29.792 7.65 29.972 7.71 ;
      RECT MASK 1 30.112 7.65 30.292 7.71 ;
      RECT MASK 1 30.456 7.65 30.636 7.71 ;
      RECT MASK 1 30.776 7.65 30.956 7.71 ;
      RECT MASK 1 31.12 7.65 31.3 7.71 ;
      RECT MASK 1 31.44 7.65 31.62 7.71 ;
      RECT MASK 1 29.028 7.89 31.2 7.95 ;
      RECT MASK 1 31.784 7.89 31.964 7.95 ;
      RECT MASK 1 29.123 8.13 31.886 8.19 ;
      RECT MASK 1 29.349 8.37 29.628 8.43 ;
      RECT MASK 1 30.013 8.37 30.292 8.43 ;
      RECT MASK 1 30.677 8.37 30.956 8.43 ;
      RECT MASK 1 31.341 8.37 31.62 8.43 ;
      RECT MASK 1 29.121 8.74 31.871 8.78 ;
      RECT MASK 1 29.121 9.16 31.871 9.2 ;
      RECT MASK 1 1.632 9.199 2.07 9.339 ;
      RECT MASK 1 2.398 9.199 2.836 9.339 ;
      RECT MASK 1 3.164 9.199 3.602 9.339 ;
      RECT MASK 1 3.93 9.199 5.134 9.339 ;
      RECT MASK 1 5.462 9.199 6.666 9.339 ;
      RECT MASK 1 6.994 9.199 8.198 9.339 ;
      RECT MASK 1 8.526 9.199 9.73 9.339 ;
      RECT MASK 1 10.058 9.199 11.262 9.339 ;
      RECT MASK 1 11.59 9.199 12.794 9.339 ;
      RECT MASK 1 13.122 9.199 14.326 9.339 ;
      RECT MASK 1 14.654 9.199 15.092 9.339 ;
      RECT MASK 1 15.42 9.199 15.858 9.339 ;
      RECT MASK 1 16.186 9.199 17.39 9.339 ;
      RECT MASK 1 17.718 9.199 18.922 9.339 ;
      RECT MASK 1 19.25 9.199 20.454 9.339 ;
      RECT MASK 1 20.782 9.199 21.986 9.339 ;
      RECT MASK 1 22.314 9.199 23.518 9.339 ;
      RECT MASK 1 23.846 9.199 25.05 9.339 ;
      RECT MASK 1 25.378 9.199 26.582 9.339 ;
      RECT MASK 1 26.885 9.199 27.348 9.339 ;
      RECT MASK 1 29.023 9.47 29.208 9.53 ;
      RECT MASK 1 29.128 9.69 31.2 9.75 ;
      RECT MASK 1 31.452 9.69 31.809 9.75 ;
      RECT MASK 1 29.334 9.93 29.651 9.99 ;
      RECT MASK 1 29.998 9.93 30.315 9.99 ;
      RECT MASK 1 30.662 9.93 30.979 9.99 ;
      RECT MASK 1 31.281 9.93 31.703 9.99 ;
      RECT MASK 1 0.662 9.97 28.157 10.01 ;
      RECT MASK 1 0.823 10.39 10.229 10.43 ;
      RECT MASK 1 11.4715 10.39 31.871 10.43 ;
      RECT MASK 1 24.984 10.62 25.064 11.88 ;
      RECT MASK 1 27.972 10.62 28.052 11.88 ;
      RECT MASK 1 0.838 10.6835 0.918 12.1765 ;
      RECT MASK 1 10.134 10.6835 10.214 12.1765 ;
      RECT MASK 1 25.654 10.71 25.714 11.76 ;
      RECT MASK 1 25.928 10.71 25.988 11.76 ;
      RECT MASK 1 26.202 10.71 26.262 11.76 ;
      RECT MASK 1 26.476 10.71 26.536 11.76 ;
      RECT MASK 1 26.75 10.71 26.81 11.76 ;
      RECT MASK 1 27.024 10.71 27.084 11.76 ;
      RECT MASK 1 27.298 10.71 27.358 11.76 ;
      RECT MASK 1 11.55 10.711 24.854 10.751 ;
      RECT MASK 1 11.55 10.886 24.854 10.926 ;
      RECT MASK 1 8.318 10.928 8.378 11.152 ;
      RECT MASK 1 8.65 10.928 8.71 11.152 ;
      RECT MASK 1 8.982 10.928 9.042 11.152 ;
      RECT MASK 1 9.314 10.928 9.374 11.152 ;
      RECT MASK 1 11.976 11.053 12.186 11.093 ;
      RECT MASK 1 12.474 11.053 12.684 11.093 ;
      RECT MASK 1 12.833 11.053 13.051 11.093 ;
      RECT MASK 1 13.165 11.053 13.383 11.093 ;
      RECT MASK 1 13.497 11.053 13.715 11.093 ;
      RECT MASK 1 13.829 11.053 14.012 11.093 ;
      RECT MASK 1 14.327 11.053 14.51 11.093 ;
      RECT MASK 1 14.964 11.053 15.174 11.093 ;
      RECT MASK 1 15.323 11.053 15.541 11.093 ;
      RECT MASK 1 15.655 11.053 15.873 11.093 ;
      RECT MASK 1 16.025 11.053 16.371 11.093 ;
      RECT MASK 1 16.689 11.053 17.035 11.093 ;
      RECT MASK 1 17.315 11.053 17.498 11.093 ;
      RECT MASK 1 17.813 11.053 18.235 11.093 ;
      RECT MASK 1 18.477 11.053 20.32 11.093 ;
      RECT MASK 1 20.469 11.053 22.312 11.093 ;
      RECT MASK 1 22.461 11.053 24.304 11.093 ;
      RECT MASK 1 11.709 11.237 11.889 11.277 ;
      RECT MASK 1 12.207 11.237 12.387 11.277 ;
      RECT MASK 1 12.705 11.237 12.885 11.277 ;
      RECT MASK 1 13.037 11.237 13.217 11.277 ;
      RECT MASK 1 13.369 11.237 13.549 11.277 ;
      RECT MASK 1 13.701 11.237 14.047 11.277 ;
      RECT MASK 1 14.199 11.237 14.545 11.277 ;
      RECT MASK 1 14.697 11.237 14.877 11.277 ;
      RECT MASK 1 15.195 11.237 15.375 11.277 ;
      RECT MASK 1 15.527 11.237 15.731 11.277 ;
      RECT MASK 1 15.859 11.237 16.039 11.277 ;
      RECT MASK 1 16.191 11.237 16.371 11.277 ;
      RECT MASK 1 16.689 11.237 17.035 11.277 ;
      RECT MASK 1 17.187 11.237 17.533 11.277 ;
      RECT MASK 1 17.685 11.237 17.996 11.277 ;
      RECT MASK 1 18.349 11.237 19.324 11.277 ;
      RECT MASK 1 20.341 11.237 21.316 11.277 ;
      RECT MASK 1 22.333 11.237 23.308 11.277 ;
      RECT MASK 1 1.43 11.286 2.186 11.346 ;
      RECT MASK 1 4.022 11.286 4.202 11.346 ;
      RECT MASK 1 4.598 11.286 4.778 11.346 ;
      RECT MASK 1 5.174 11.286 5.354 11.346 ;
      RECT MASK 1 5.75 11.286 5.93 11.346 ;
      RECT MASK 1 6.326 11.286 7.658 11.346 ;
      RECT MASK 1 11.709 11.463 11.889 11.503 ;
      RECT MASK 1 12.207 11.463 12.387 11.503 ;
      RECT MASK 1 12.705 11.463 12.885 11.503 ;
      RECT MASK 1 13.037 11.463 13.217 11.503 ;
      RECT MASK 1 13.369 11.463 13.549 11.503 ;
      RECT MASK 1 13.701 11.463 14.047 11.503 ;
      RECT MASK 1 14.199 11.463 14.545 11.503 ;
      RECT MASK 1 14.697 11.463 14.877 11.503 ;
      RECT MASK 1 15.195 11.463 15.375 11.503 ;
      RECT MASK 1 15.527 11.463 16.205 11.503 ;
      RECT MASK 1 16.357 11.463 16.714 11.503 ;
      RECT MASK 1 17.187 11.463 17.533 11.503 ;
      RECT MASK 1 17.685 11.463 17.996 11.503 ;
      RECT MASK 1 18.349 11.463 19.324 11.503 ;
      RECT MASK 1 20.341 11.463 21.316 11.503 ;
      RECT MASK 1 22.333 11.463 23.308 11.503 ;
      RECT MASK 1 1.43 11.514 2.186 11.574 ;
      RECT MASK 1 4.022 11.514 4.202 11.574 ;
      RECT MASK 1 4.598 11.514 4.778 11.574 ;
      RECT MASK 1 5.174 11.514 5.354 11.574 ;
      RECT MASK 1 5.75 11.514 5.93 11.574 ;
      RECT MASK 1 6.326 11.514 6.506 11.574 ;
      RECT MASK 1 6.902 11.514 7.658 11.574 ;
      RECT MASK 1 11.837 11.647 12.186 11.687 ;
      RECT MASK 1 12.335 11.647 12.684 11.687 ;
      RECT MASK 1 12.833 11.647 13.051 11.687 ;
      RECT MASK 1 13.165 11.647 13.383 11.687 ;
      RECT MASK 1 13.497 11.647 13.715 11.687 ;
      RECT MASK 1 13.829 11.647 14.012 11.687 ;
      RECT MASK 1 14.327 11.647 14.51 11.687 ;
      RECT MASK 1 14.825 11.647 15.174 11.687 ;
      RECT MASK 1 15.323 11.647 15.541 11.687 ;
      RECT MASK 1 15.655 11.647 15.873 11.687 ;
      RECT MASK 1 16.025 11.647 16.369 11.687 ;
      RECT MASK 1 16.807 11.647 17.035 11.687 ;
      RECT MASK 1 17.315 11.647 17.498 11.687 ;
      RECT MASK 1 17.813 11.647 18.235 11.687 ;
      RECT MASK 1 18.477 11.647 20.32 11.687 ;
      RECT MASK 1 20.469 11.647 22.312 11.687 ;
      RECT MASK 1 22.461 11.647 24.304 11.687 ;
      RECT MASK 1 8.318 11.708 8.378 11.932 ;
      RECT MASK 1 8.65 11.708 8.71 11.932 ;
      RECT MASK 1 8.982 11.708 9.042 11.932 ;
      RECT MASK 1 9.314 11.708 9.374 11.932 ;
      RECT MASK 1 11.55 11.814 24.498 11.854 ;
      RECT MASK 1 11.55 11.989 24.498 12.029 ;
      RECT MASK 1 24.969 12.07 28.067 12.11 ;
      RECT MASK 1 8.175 12.086 9.688 12.146 ;
      RECT MASK 1 11.4715 12.31 24.451 12.35 ;
      RECT MASK 1 0.759 12.43 10.293 12.47 ;
      RECT MASK 1 20.987 12.73 31.832 12.77 ;
      RECT MASK 1 0.759 12.85 10.293 12.89 ;
      RECT MASK 1 21.002 13.0235 21.082 24.6565 ;
      RECT MASK 1 25.65 13.0235 25.73 24.6565 ;
      RECT MASK 1 26.222 13.0235 26.302 24.6565 ;
      RECT MASK 1 31.7 13.0235 31.78 24.6565 ;
      RECT MASK 1 0.838 13.1435 0.918 14.6365 ;
      RECT MASK 1 10.134 13.1435 10.214 14.6365 ;
      RECT MASK 1 21.651 13.17 22.088 13.21 ;
      RECT MASK 1 22.647 13.17 24.085 13.21 ;
      RECT MASK 1 24.312 13.17 25.081 13.21 ;
      RECT MASK 1 7.7425 13.174 9.667 13.234 ;
      RECT MASK 1 12.343 13.36 15.579 13.4 ;
      RECT MASK 1 15.885 13.36 16.659 13.4 ;
      RECT MASK 1 22.149 13.37 24.744 13.41 ;
      RECT MASK 1 8.318 13.388 8.378 13.612 ;
      RECT MASK 1 8.65 13.388 8.71 13.612 ;
      RECT MASK 1 8.982 13.388 9.042 13.612 ;
      RECT MASK 1 9.314 13.388 9.374 13.612 ;
      RECT MASK 1 24.971 13.56 25.159 13.6 ;
      RECT MASK 1 21.573 13.57 21.761 13.61 ;
      RECT MASK 1 21.905 13.57 24.827 13.61 ;
      RECT MASK 1 3.446 13.756 5.066 13.816 ;
      RECT MASK 1 5.462 13.756 6.218 13.816 ;
      RECT MASK 1 12.534 13.838 12.594 14.088 ;
      RECT MASK 1 12.866 13.838 12.926 14.088 ;
      RECT MASK 1 14.102 13.838 14.162 14.068 ;
      RECT MASK 1 14.434 13.838 14.494 14.068 ;
      RECT MASK 1 16.242 13.838 16.302 14.0485 ;
      RECT MASK 1 21.485 13.87 23.582 13.91 ;
      RECT MASK 1 17.1785 13.942 19.876 13.966 ;
      RECT MASK 1 2.87 13.964 3.05 14.024 ;
      RECT MASK 1 3.446 13.964 5.066 14.024 ;
      RECT MASK 1 5.462 13.964 6.218 14.024 ;
      RECT MASK 1 6.614 13.964 6.794 14.024 ;
      RECT MASK 1 21.822 14.07 24.91 14.11 ;
      RECT MASK 1 13.304 14.0875 13.484 14.1275 ;
      RECT MASK 1 15.278 14.0875 15.458 14.1275 ;
      RECT MASK 1 17.1785 14.122 19.876 14.146 ;
      RECT MASK 1 8.318 14.168 8.378 14.392 ;
      RECT MASK 1 8.65 14.168 8.71 14.392 ;
      RECT MASK 1 8.982 14.168 9.042 14.392 ;
      RECT MASK 1 9.314 14.168 9.374 14.392 ;
      RECT MASK 1 21.739 14.27 24.993 14.31 ;
      RECT MASK 1 17.4665 14.298 19.655 14.322 ;
      RECT MASK 1 12.509 14.309 12.858 14.349 ;
      RECT MASK 1 14.17 14.309 14.353 14.349 ;
      RECT MASK 1 15.192 14.309 16.83 14.349 ;
      RECT MASK 1 27.2165 14.349 27.6945 14.489 ;
      RECT MASK 1 28.0225 14.349 29.3065 14.489 ;
      RECT MASK 1 29.6345 14.349 30.9185 14.489 ;
      RECT MASK 1 21.739 14.47 24.993 14.51 ;
      RECT MASK 1 12.343 14.511 12.692 14.551 ;
      RECT MASK 1 14.409 14.511 14.592 14.551 ;
      RECT MASK 1 15.147 14.511 16.9905 14.551 ;
      RECT MASK 1 7.7425 14.546 9.667 14.606 ;
      RECT MASK 1 21.822 14.67 24.91 14.71 ;
      RECT MASK 1 13.304 14.7325 13.484 14.7725 ;
      RECT MASK 1 15.278 14.7325 15.458 14.7725 ;
      RECT MASK 1 17.1915 14.748 17.5255 14.772 ;
      RECT MASK 1 17.778 14.748 19.876 14.772 ;
      RECT MASK 1 12.534 14.772 12.594 15.022 ;
      RECT MASK 1 12.866 14.772 12.926 15.022 ;
      RECT MASK 1 14.102 14.792 14.162 15.022 ;
      RECT MASK 1 14.434 14.792 14.494 15.022 ;
      RECT MASK 1 16.242 14.811 16.302 15.022 ;
      RECT MASK 1 17.1915 14.838 17.476 14.862 ;
      RECT MASK 1 17.839 14.838 19.338 14.862 ;
      RECT MASK 1 21.485 14.87 23.582 14.91 ;
      RECT MASK 1 0.823 14.89 10.293 14.93 ;
      RECT MASK 1 16.964 15.258 19.876 15.282 ;
      RECT MASK 1 21.485 15.28 23.582 15.32 ;
      RECT MASK 1 0.825 15.43 1.583 15.47 ;
      RECT MASK 1 2.123 15.46 10.518 15.5 ;
      RECT MASK 1 21.822 15.48 24.91 15.52 ;
      RECT MASK 1 12.534 15.518 12.594 15.768 ;
      RECT MASK 1 12.866 15.518 12.926 15.768 ;
      RECT MASK 1 14.102 15.518 14.162 15.748 ;
      RECT MASK 1 14.434 15.518 14.494 15.748 ;
      RECT MASK 1 16.242 15.518 16.302 15.729 ;
      RECT MASK 1 17.1915 15.678 17.476 15.702 ;
      RECT MASK 1 17.839 15.678 19.338 15.702 ;
      RECT MASK 1 21.739 15.68 24.993 15.72 ;
      RECT MASK 1 13.304 15.7675 13.484 15.8075 ;
      RECT MASK 1 15.278 15.7675 15.458 15.8075 ;
      RECT MASK 1 17.1915 15.768 17.5255 15.792 ;
      RECT MASK 1 17.778 15.768 19.876 15.792 ;
      RECT MASK 1 1.038 15.87 1.355 15.93 ;
      RECT MASK 1 2.718 15.96 2.778 17.01 ;
      RECT MASK 1 2.992 15.96 3.052 17.01 ;
      RECT MASK 1 3.266 15.96 3.326 17.01 ;
      RECT MASK 1 3.54 15.96 3.6 17.01 ;
      RECT MASK 1 3.814 15.96 3.874 17.01 ;
      RECT MASK 1 4.088 15.96 4.148 17.01 ;
      RECT MASK 1 4.362 15.96 4.422 17.01 ;
      RECT MASK 1 4.636 15.96 4.696 17.01 ;
      RECT MASK 1 4.91 15.96 4.97 17.01 ;
      RECT MASK 1 5.184 15.96 5.244 17.01 ;
      RECT MASK 1 5.458 15.96 5.518 17.01 ;
      RECT MASK 1 5.732 15.96 5.792 17.01 ;
      RECT MASK 1 6.006 15.96 6.066 17.01 ;
      RECT MASK 1 6.28 15.96 6.34 17.01 ;
      RECT MASK 1 6.554 15.96 6.614 17.01 ;
      RECT MASK 1 6.828 15.96 6.888 17.01 ;
      RECT MASK 1 7.102 15.96 7.162 17.01 ;
      RECT MASK 1 7.376 15.96 7.436 17.01 ;
      RECT MASK 1 7.65 15.96 7.71 17.01 ;
      RECT MASK 1 7.924 15.96 7.984 17.01 ;
      RECT MASK 1 8.198 15.96 8.258 17.01 ;
      RECT MASK 1 8.472 15.96 8.532 17.01 ;
      RECT MASK 1 8.746 15.96 8.806 17.01 ;
      RECT MASK 1 9.02 15.96 9.08 17.01 ;
      RECT MASK 1 9.294 15.96 9.354 17.01 ;
      RECT MASK 1 9.568 15.96 9.628 17.01 ;
      RECT MASK 1 9.842 15.96 9.902 17.01 ;
      RECT MASK 1 10.116 15.96 10.176 17.01 ;
      RECT MASK 1 10.39 15.96 10.45 17.01 ;
      RECT MASK 1 12.343 15.989 12.692 16.029 ;
      RECT MASK 1 14.409 15.989 14.592 16.029 ;
      RECT MASK 1 15.147 15.989 16.9905 16.029 ;
      RECT MASK 1 21.948 15.99 22.128 16.03 ;
      RECT MASK 1 22.28 15.99 22.46 16.03 ;
      RECT MASK 1 22.743 15.99 22.923 16.03 ;
      RECT MASK 1 23.15 15.99 24.251 16.03 ;
      RECT MASK 1 0.832 16.11 1.576 16.17 ;
      RECT MASK 1 2.118 16.145 2.238 16.225 ;
      RECT MASK 1 21.817 16.19 22.259 16.23 ;
      RECT MASK 1 22.486 16.19 23.089 16.23 ;
      RECT MASK 1 12.509 16.191 12.858 16.231 ;
      RECT MASK 1 14.17 16.191 14.353 16.231 ;
      RECT MASK 1 15.192 16.191 16.83 16.231 ;
      RECT MASK 1 17.4665 16.218 19.655 16.242 ;
      RECT MASK 1 0.727 16.33 0.912 16.39 ;
      RECT MASK 1 22.071 16.39 22.259 16.43 ;
      RECT MASK 1 22.403 16.39 22.591 16.43 ;
      RECT MASK 1 17.1785 16.394 19.876 16.418 ;
      RECT MASK 1 13.304 16.4125 13.484 16.4525 ;
      RECT MASK 1 15.278 16.4125 15.458 16.4525 ;
      RECT MASK 1 12.534 16.452 12.594 16.702 ;
      RECT MASK 1 12.866 16.452 12.926 16.702 ;
      RECT MASK 1 14.102 16.472 14.162 16.702 ;
      RECT MASK 1 14.434 16.472 14.494 16.702 ;
      RECT MASK 1 16.242 16.4915 16.302 16.702 ;
      RECT MASK 1 17.1785 16.574 19.876 16.598 ;
      RECT MASK 1 0.825 16.66 1.583 16.7 ;
      RECT MASK 1 2.118 16.745 2.238 16.825 ;
      RECT MASK 1 21.651 16.94 25.081 16.98 ;
      RECT MASK 1 0.825 17.08 1.583 17.12 ;
      RECT MASK 1 12.343 17.14 15.579 17.18 ;
      RECT MASK 1 15.885 17.14 16.659 17.18 ;
      RECT MASK 1 21.573 17.14 22.005 17.18 ;
      RECT MASK 1 22.237 17.14 22.757 17.18 ;
      RECT MASK 1 22.901 17.14 25.159 17.18 ;
      RECT MASK 1 1.053 17.43 1.332 17.49 ;
      RECT MASK 1 21.651 17.47 25.081 17.51 ;
      RECT MASK 1 2.718 17.55 2.778 18.6 ;
      RECT MASK 1 2.992 17.55 3.052 18.6 ;
      RECT MASK 1 3.266 17.55 3.326 18.6 ;
      RECT MASK 1 3.54 17.55 3.6 18.6 ;
      RECT MASK 1 3.814 17.55 3.874 18.6 ;
      RECT MASK 1 4.088 17.55 4.148 18.6 ;
      RECT MASK 1 4.362 17.55 4.422 18.6 ;
      RECT MASK 1 4.636 17.55 4.696 18.6 ;
      RECT MASK 1 4.91 17.55 4.97 18.6 ;
      RECT MASK 1 5.184 17.55 5.244 18.6 ;
      RECT MASK 1 5.458 17.55 5.518 18.6 ;
      RECT MASK 1 5.732 17.55 5.792 18.6 ;
      RECT MASK 1 6.006 17.55 6.066 18.6 ;
      RECT MASK 1 6.28 17.55 6.34 18.6 ;
      RECT MASK 1 0.827 17.67 1.598 17.73 ;
      RECT MASK 1 2.118 17.735 2.238 17.815 ;
      RECT MASK 1 23.477 17.81 23.665 17.85 ;
      RECT MASK 1 0.732 17.91 1.676 17.97 ;
      RECT MASK 1 21.651 18.11 23.587 18.15 ;
      RECT MASK 1 0.832 18.15 1.012 18.21 ;
      RECT MASK 1 1.152 18.15 1.332 18.21 ;
      RECT MASK 1 7.195 18.16 20.215 18.2 ;
      RECT MASK 1 21.573 18.31 21.839 18.35 ;
      RECT MASK 1 22.071 18.31 23.499 18.35 ;
      RECT MASK 1 2.118 18.335 2.238 18.415 ;
      RECT MASK 1 1.053 18.39 1.233 18.45 ;
      RECT MASK 1 1.396 18.39 1.576 18.45 ;
      RECT MASK 1 27.2165 18.429 28.5005 18.569 ;
      RECT MASK 1 28.8285 18.429 30.1125 18.569 ;
      RECT MASK 1 30.4405 18.429 31.135 18.569 ;
      RECT MASK 1 7.148 18.481 20.262 18.521 ;
      RECT MASK 1 21.573 18.56 21.839 18.6 ;
      RECT MASK 1 22.071 18.56 23.499 18.6 ;
      RECT MASK 1 1.076 18.63 1.256 18.69 ;
      RECT MASK 1 1.396 18.63 1.576 18.69 ;
      RECT MASK 1 7.148 18.646 20.262 18.686 ;
      RECT MASK 1 21.651 18.76 23.587 18.8 ;
      RECT MASK 1 27.2165 18.819 28.5005 18.959 ;
      RECT MASK 1 28.8285 18.819 30.1125 18.959 ;
      RECT MASK 1 30.4405 18.819 30.9185 18.959 ;
      RECT MASK 1 7.574 18.823 7.784 18.863 ;
      RECT MASK 1 8.072 18.823 8.282 18.863 ;
      RECT MASK 1 8.57 18.823 8.78 18.863 ;
      RECT MASK 1 9.095 18.823 9.313 18.863 ;
      RECT MASK 1 9.593 18.823 10.689 18.863 ;
      RECT MASK 1 10.921 18.823 12.017 18.863 ;
      RECT MASK 1 12.249 18.823 13.345 18.863 ;
      RECT MASK 1 13.577 18.823 14.673 18.863 ;
      RECT MASK 1 14.905 18.823 16.001 18.863 ;
      RECT MASK 1 16.233 18.823 17.329 18.863 ;
      RECT MASK 1 17.561 18.823 18.657 18.863 ;
      RECT MASK 1 18.889 18.823 19.985 18.863 ;
      RECT MASK 1 0.835 18.87 1.015 18.93 ;
      RECT MASK 1 1.135 18.87 1.355 18.93 ;
      RECT MASK 1 7.307 19.007 7.487 19.047 ;
      RECT MASK 1 7.805 19.007 7.985 19.047 ;
      RECT MASK 1 8.303 19.007 8.483 19.047 ;
      RECT MASK 1 8.967 19.007 9.313 19.047 ;
      RECT MASK 1 9.452 19.007 10.103 19.047 ;
      RECT MASK 1 10.78 19.007 11.431 19.047 ;
      RECT MASK 1 12.108 19.007 12.759 19.047 ;
      RECT MASK 1 13.436 19.007 14.087 19.047 ;
      RECT MASK 1 14.764 19.007 15.415 19.047 ;
      RECT MASK 1 16.092 19.007 16.743 19.047 ;
      RECT MASK 1 17.42 19.007 18.071 19.047 ;
      RECT MASK 1 18.748 19.007 19.399 19.047 ;
      RECT MASK 1 5.322 19.1 6.522 19.12 ;
      RECT MASK 1 2.718 19.14 2.778 20.19 ;
      RECT MASK 1 2.992 19.14 3.052 20.19 ;
      RECT MASK 1 3.266 19.14 3.326 20.19 ;
      RECT MASK 1 3.54 19.14 3.6 20.19 ;
      RECT MASK 1 3.814 19.14 3.874 20.19 ;
      RECT MASK 1 4.088 19.14 4.148 20.19 ;
      RECT MASK 1 4.362 19.14 4.422 20.19 ;
      RECT MASK 1 0.825 19.21 1.583 19.25 ;
      RECT MASK 1 7.307 19.233 7.487 19.273 ;
      RECT MASK 1 7.805 19.233 7.985 19.273 ;
      RECT MASK 1 8.303 19.233 8.483 19.273 ;
      RECT MASK 1 8.967 19.233 9.313 19.273 ;
      RECT MASK 1 9.452 19.233 10.103 19.273 ;
      RECT MASK 1 10.78 19.233 11.431 19.273 ;
      RECT MASK 1 12.108 19.233 12.759 19.273 ;
      RECT MASK 1 13.436 19.233 14.087 19.273 ;
      RECT MASK 1 14.764 19.233 15.415 19.273 ;
      RECT MASK 1 16.092 19.233 16.743 19.273 ;
      RECT MASK 1 17.42 19.233 18.071 19.273 ;
      RECT MASK 1 18.748 19.233 19.399 19.273 ;
      RECT MASK 1 2.118 19.325 2.238 19.405 ;
      RECT MASK 1 5.322 19.34 6.522 19.36 ;
      RECT MASK 1 7.435 19.417 7.784 19.457 ;
      RECT MASK 1 7.933 19.417 8.282 19.457 ;
      RECT MASK 1 8.431 19.417 8.78 19.457 ;
      RECT MASK 1 8.967 19.417 9.185 19.457 ;
      RECT MASK 1 9.593 19.417 10.689 19.457 ;
      RECT MASK 1 10.921 19.417 12.017 19.457 ;
      RECT MASK 1 12.249 19.417 13.345 19.457 ;
      RECT MASK 1 13.577 19.417 14.673 19.457 ;
      RECT MASK 1 14.905 19.417 16.001 19.457 ;
      RECT MASK 1 16.233 19.417 17.329 19.457 ;
      RECT MASK 1 17.561 19.417 18.657 19.457 ;
      RECT MASK 1 18.889 19.417 19.985 19.457 ;
      RECT MASK 1 5.322 19.42 6.522 19.44 ;
      RECT MASK 1 5.322 19.5 6.522 19.52 ;
      RECT MASK 1 21.651 19.54 23.919 19.58 ;
      RECT MASK 1 5.322 19.58 6.522 19.6 ;
      RECT MASK 1 7.148 19.594 20.359 19.634 ;
      RECT MASK 1 0.825 19.63 1.583 19.67 ;
      RECT MASK 1 5.322 19.66 6.522 19.68 ;
      RECT MASK 1 5.322 19.74 6.522 19.76 ;
      RECT MASK 1 21.573 19.74 21.839 19.78 ;
      RECT MASK 1 22.071 19.74 23.665 19.78 ;
      RECT MASK 1 23.809 19.74 23.997 19.78 ;
      RECT MASK 1 7.148 19.759 20.359 19.799 ;
      RECT MASK 1 5.322 19.82 6.522 19.84 ;
      RECT MASK 1 2.118 19.925 2.238 20.005 ;
      RECT MASK 1 5.322 20.06 6.522 20.08 ;
      RECT MASK 1 0.832 20.07 1.598 20.13 ;
      RECT MASK 1 7.195 20.08 20.344 20.12 ;
      RECT MASK 1 21.988 20.3 23.748 20.34 ;
      RECT MASK 1 0.953 20.31 1.133 20.37 ;
      RECT MASK 1 1.275 20.31 1.455 20.37 ;
      RECT MASK 1 13.996 20.401 20.636 20.441 ;
      RECT MASK 1 21.905 20.5 23.831 20.54 ;
      RECT MASK 1 0.832 20.55 1.598 20.61 ;
      RECT MASK 1 13.996 20.576 20.636 20.616 ;
      RECT MASK 1 14.947 20.743 15.13 20.783 ;
      RECT MASK 1 15.445 20.743 15.867 20.783 ;
      RECT MASK 1 16.109 20.743 17.288 20.783 ;
      RECT MASK 1 17.437 20.743 18.616 20.783 ;
      RECT MASK 1 18.765 20.743 19.944 20.783 ;
      RECT MASK 1 6.074 20.8 13.543 20.84 ;
      RECT MASK 1 21.651 20.83 25.081 20.87 ;
      RECT MASK 1 14.072 20.8375 14.252 20.8775 ;
      RECT MASK 1 20.38 20.8375 20.56 20.8775 ;
      RECT MASK 1 14.819 20.927 15.165 20.967 ;
      RECT MASK 1 15.317 20.927 15.628 20.967 ;
      RECT MASK 1 15.981 20.927 16.659 20.967 ;
      RECT MASK 1 17.309 20.927 17.987 20.967 ;
      RECT MASK 1 18.637 20.927 19.315 20.967 ;
      RECT MASK 1 2.108 21.01 3.2225 21.05 ;
      RECT MASK 1 3.948 21.01 4.566 21.05 ;
      RECT MASK 1 5.152 21.01 5.684 21.05 ;
      RECT MASK 1 0.953 21.03 1.133 21.09 ;
      RECT MASK 1 1.275 21.03 1.455 21.09 ;
      RECT MASK 1 14.819 21.153 15.165 21.193 ;
      RECT MASK 1 15.317 21.153 15.628 21.193 ;
      RECT MASK 1 15.981 21.153 16.659 21.193 ;
      RECT MASK 1 17.309 21.153 17.987 21.193 ;
      RECT MASK 1 18.637 21.153 19.315 21.193 ;
      RECT MASK 1 14.072 21.2425 14.252 21.2825 ;
      RECT MASK 1 20.38 21.2425 20.56 21.2825 ;
      RECT MASK 1 0.953 21.27 1.133 21.33 ;
      RECT MASK 1 1.275 21.27 1.455 21.33 ;
      RECT MASK 1 6.056 21.278 6.116 21.508 ;
      RECT MASK 1 6.388 21.278 6.448 21.508 ;
      RECT MASK 1 6.72 21.278 6.78 21.508 ;
      RECT MASK 1 7.052 21.278 7.112 21.508 ;
      RECT MASK 1 7.384 21.278 7.444 21.508 ;
      RECT MASK 1 7.716 21.278 7.776 21.508 ;
      RECT MASK 1 8.048 21.278 8.108 21.508 ;
      RECT MASK 1 8.38 21.278 8.44 21.508 ;
      RECT MASK 1 8.712 21.278 8.772 21.508 ;
      RECT MASK 1 9.044 21.278 9.104 21.508 ;
      RECT MASK 1 9.376 21.278 9.436 21.508 ;
      RECT MASK 1 10.103 21.278 10.163 21.508 ;
      RECT MASK 1 10.767 21.278 10.827 21.508 ;
      RECT MASK 1 11.099 21.278 11.159 21.508 ;
      RECT MASK 1 11.431 21.278 11.491 21.508 ;
      RECT MASK 1 11.763 21.278 11.823 21.508 ;
      RECT MASK 1 12.095 21.278 12.155 21.508 ;
      RECT MASK 1 12.676 21.278 12.736 21.508 ;
      RECT MASK 1 13.008 21.278 13.068 21.508 ;
      RECT MASK 1 13.34 21.278 13.4 21.508 ;
      RECT MASK 1 2.212 21.288 3.159 21.312 ;
      RECT MASK 1 14.947 21.337 15.13 21.377 ;
      RECT MASK 1 15.445 21.337 15.867 21.377 ;
      RECT MASK 1 16.109 21.337 17.288 21.377 ;
      RECT MASK 1 17.437 21.337 18.616 21.377 ;
      RECT MASK 1 18.765 21.337 19.944 21.377 ;
      RECT MASK 1 2.212 21.378 3.159 21.402 ;
      RECT MASK 1 3.955 21.416 5.913 21.456 ;
      RECT MASK 1 2.422 21.468 2.874 21.492 ;
      RECT MASK 1 13.996 21.504 20.636 21.544 ;
      RECT MASK 1 0.732 21.54 0.912 21.6 ;
      RECT MASK 1 1.242 21.54 1.498 21.6 ;
      RECT MASK 1 2.422 21.558 2.644 21.582 ;
      RECT MASK 1 4.27 21.602 4.33 21.832 ;
      RECT MASK 1 5.496 21.602 5.556 21.832 ;
      RECT MASK 1 13.996 21.679 20.636 21.719 ;
      RECT MASK 1 6.015 21.749 9.413 21.789 ;
      RECT MASK 1 9.746 21.749 11.63 21.789 ;
      RECT MASK 1 11.738 21.749 12.05 21.789 ;
      RECT MASK 1 12.255 21.749 13.068 21.789 ;
      RECT MASK 1 2.135 21.755 3.0545 21.795 ;
      RECT MASK 1 13.996 21.841 20.636 21.881 ;
      RECT MASK 1 2.392 21.951 2.841 21.991 ;
      RECT MASK 1 5.637 21.951 10.306 21.991 ;
      RECT MASK 1 10.741 21.951 11.116 21.991 ;
      RECT MASK 1 11.24 21.951 11.634 21.991 ;
      RECT MASK 1 11.952 21.951 12.132 21.991 ;
      RECT MASK 1 12.485 21.951 12.927 21.991 ;
      RECT MASK 1 13.061 21.951 13.425 21.991 ;
      RECT MASK 1 0.732 21.96 0.912 22.02 ;
      RECT MASK 1 1.242 21.96 1.498 22.02 ;
      RECT MASK 1 13.996 22.016 20.636 22.056 ;
      RECT MASK 1 14.781 22.183 15.203 22.223 ;
      RECT MASK 1 15.445 22.183 15.867 22.223 ;
      RECT MASK 1 16.109 22.183 17.288 22.223 ;
      RECT MASK 1 17.437 22.183 18.616 22.223 ;
      RECT MASK 1 18.765 22.183 19.944 22.223 ;
      RECT MASK 1 2.136 22.203 3.159 22.227 ;
      RECT MASK 1 23.315 22.21 23.653 22.23 ;
      RECT MASK 1 23.905 22.21 24.2605 22.23 ;
      RECT MASK 1 0.953 22.23 1.133 22.29 ;
      RECT MASK 1 1.275 22.23 1.455 22.29 ;
      RECT MASK 1 6.056 22.232 6.116 22.462 ;
      RECT MASK 1 6.388 22.232 6.448 22.462 ;
      RECT MASK 1 6.72 22.232 6.78 22.462 ;
      RECT MASK 1 7.052 22.232 7.112 22.462 ;
      RECT MASK 1 7.384 22.232 7.444 22.462 ;
      RECT MASK 1 7.716 22.232 7.776 22.462 ;
      RECT MASK 1 8.048 22.232 8.108 22.462 ;
      RECT MASK 1 8.38 22.232 8.44 22.462 ;
      RECT MASK 1 8.712 22.232 8.772 22.462 ;
      RECT MASK 1 9.044 22.232 9.104 22.462 ;
      RECT MASK 1 9.376 22.232 9.436 22.462 ;
      RECT MASK 1 10.103 22.232 10.163 22.462 ;
      RECT MASK 1 10.435 22.232 10.495 22.462 ;
      RECT MASK 1 10.767 22.232 10.827 22.462 ;
      RECT MASK 1 11.099 22.232 11.159 22.462 ;
      RECT MASK 1 11.431 22.232 11.491 22.462 ;
      RECT MASK 1 11.763 22.232 11.823 22.462 ;
      RECT MASK 1 12.095 22.232 12.155 22.462 ;
      RECT MASK 1 12.676 22.232 12.736 22.462 ;
      RECT MASK 1 13.008 22.232 13.068 22.462 ;
      RECT MASK 1 13.34 22.232 13.4 22.462 ;
      RECT MASK 1 14.072 22.2775 14.252 22.3175 ;
      RECT MASK 1 20.38 22.2775 20.56 22.3175 ;
      RECT MASK 1 22.4955 22.29 23.305 22.31 ;
      RECT MASK 1 2.422 22.293 2.874 22.317 ;
      RECT MASK 1 4.27 22.328 4.33 22.558 ;
      RECT MASK 1 5.496 22.328 5.556 22.558 ;
      RECT MASK 1 14.653 22.367 14.964 22.407 ;
      RECT MASK 1 15.317 22.367 15.628 22.407 ;
      RECT MASK 1 15.981 22.367 16.659 22.407 ;
      RECT MASK 1 17.309 22.367 17.987 22.407 ;
      RECT MASK 1 18.637 22.367 19.315 22.407 ;
      RECT MASK 1 22.698 22.37 23.305 22.39 ;
      RECT MASK 1 2.422 22.383 2.874 22.407 ;
      RECT MASK 1 4.813 22.43 4.873 22.57 ;
      RECT MASK 1 23.905 22.45 24.2605 22.47 ;
      RECT MASK 1 0.953 22.47 1.133 22.53 ;
      RECT MASK 1 1.275 22.47 1.455 22.53 ;
      RECT MASK 1 2.136 22.473 3.159 22.497 ;
      RECT MASK 1 23.265 22.53 23.6545 22.55 ;
      RECT MASK 1 14.653 22.593 14.964 22.633 ;
      RECT MASK 1 15.317 22.593 15.628 22.633 ;
      RECT MASK 1 15.981 22.593 16.659 22.633 ;
      RECT MASK 1 17.309 22.593 17.987 22.633 ;
      RECT MASK 1 18.637 22.593 19.315 22.633 ;
      RECT MASK 1 14.072 22.6825 14.252 22.7225 ;
      RECT MASK 1 20.38 22.6825 20.56 22.7225 ;
      RECT MASK 1 22.46 22.69 24.26 22.71 ;
      RECT MASK 1 22.46 22.77 24.26 22.79 ;
      RECT MASK 1 14.781 22.777 15.203 22.817 ;
      RECT MASK 1 15.445 22.777 15.867 22.817 ;
      RECT MASK 1 16.109 22.777 17.288 22.817 ;
      RECT MASK 1 17.437 22.777 18.616 22.817 ;
      RECT MASK 1 18.765 22.777 19.944 22.817 ;
      RECT MASK 1 6.046 22.9 9.626 22.94 ;
      RECT MASK 1 10.081 22.9 13.543 22.94 ;
      RECT MASK 1 13.996 22.944 20.636 22.984 ;
      RECT MASK 1 0.825 23.05 1.583 23.09 ;
      RECT MASK 1 13.996 23.119 20.636 23.159 ;
      RECT MASK 1 27.2165 23.199 27.6945 23.339 ;
      RECT MASK 1 28.0225 23.199 29.3065 23.339 ;
      RECT MASK 1 29.6345 23.199 30.9185 23.339 ;
      RECT MASK 1 4.813 23.27 4.873 23.41 ;
      RECT MASK 1 13.996 23.281 20.636 23.321 ;
      RECT MASK 1 4.27 23.282 4.33 23.512 ;
      RECT MASK 1 5.496 23.282 5.556 23.512 ;
      RECT MASK 1 23.315 23.31 23.753 23.33 ;
      RECT MASK 1 2.136 23.343 3.159 23.367 ;
      RECT MASK 1 6.056 23.378 6.116 23.608 ;
      RECT MASK 1 6.388 23.378 6.448 23.608 ;
      RECT MASK 1 6.72 23.378 6.78 23.608 ;
      RECT MASK 1 7.052 23.378 7.112 23.608 ;
      RECT MASK 1 7.384 23.378 7.444 23.608 ;
      RECT MASK 1 7.716 23.378 7.776 23.608 ;
      RECT MASK 1 8.048 23.378 8.108 23.608 ;
      RECT MASK 1 8.38 23.378 8.44 23.608 ;
      RECT MASK 1 8.712 23.378 8.772 23.608 ;
      RECT MASK 1 9.044 23.378 9.104 23.608 ;
      RECT MASK 1 9.376 23.378 9.436 23.608 ;
      RECT MASK 1 10.103 23.378 10.163 23.608 ;
      RECT MASK 1 10.435 23.378 10.495 23.608 ;
      RECT MASK 1 10.767 23.378 10.827 23.608 ;
      RECT MASK 1 11.099 23.378 11.159 23.608 ;
      RECT MASK 1 11.431 23.378 11.491 23.608 ;
      RECT MASK 1 11.763 23.378 11.823 23.608 ;
      RECT MASK 1 12.095 23.378 12.155 23.608 ;
      RECT MASK 1 12.676 23.378 12.736 23.608 ;
      RECT MASK 1 13.008 23.378 13.068 23.608 ;
      RECT MASK 1 13.34 23.378 13.4 23.608 ;
      RECT MASK 1 23.315 23.39 23.753 23.41 ;
      RECT MASK 1 2.422 23.433 2.874 23.457 ;
      RECT MASK 1 13.996 23.456 20.636 23.496 ;
      RECT MASK 1 0.825 23.47 1.583 23.51 ;
      RECT MASK 1 2.422 23.523 2.874 23.547 ;
      RECT MASK 1 22.488 23.55 23.472 23.57 ;
      RECT MASK 1 23.905 23.55 24.2605 23.57 ;
      RECT MASK 1 2.136 23.613 3.159 23.637 ;
      RECT MASK 1 14.781 23.623 15.96 23.663 ;
      RECT MASK 1 16.109 23.623 17.288 23.663 ;
      RECT MASK 1 17.437 23.623 18.616 23.663 ;
      RECT MASK 1 18.765 23.623 19.944 23.663 ;
      RECT MASK 1 14.072 23.7175 14.252 23.7575 ;
      RECT MASK 1 20.38 23.7175 20.56 23.7575 ;
      RECT MASK 1 14.653 23.807 15.331 23.847 ;
      RECT MASK 1 15.981 23.807 16.659 23.847 ;
      RECT MASK 1 17.309 23.807 17.987 23.847 ;
      RECT MASK 1 18.637 23.807 19.315 23.847 ;
      RECT MASK 1 0.9405 23.845 1.4715 23.885 ;
      RECT MASK 1 2.392 23.849 2.841 23.889 ;
      RECT MASK 1 5.637 23.849 10.306 23.889 ;
      RECT MASK 1 10.741 23.849 11.116 23.889 ;
      RECT MASK 1 11.24 23.849 11.634 23.889 ;
      RECT MASK 1 11.952 23.849 12.132 23.889 ;
      RECT MASK 1 12.485 23.849 12.927 23.889 ;
      RECT MASK 1 13.061 23.849 13.425 23.889 ;
      RECT MASK 1 0.984 24.005 1.4145 24.045 ;
      RECT MASK 1 4.27 24.008 4.33 24.238 ;
      RECT MASK 1 5.496 24.008 5.556 24.238 ;
      RECT MASK 1 14.653 24.033 15.331 24.073 ;
      RECT MASK 1 15.981 24.033 16.659 24.073 ;
      RECT MASK 1 17.309 24.033 17.987 24.073 ;
      RECT MASK 1 18.637 24.033 19.315 24.073 ;
      RECT MASK 1 2.422 24.045 3.583 24.085 ;
      RECT MASK 1 6.015 24.051 9.413 24.091 ;
      RECT MASK 1 9.746 24.051 11.63 24.091 ;
      RECT MASK 1 11.738 24.051 12.05 24.091 ;
      RECT MASK 1 12.255 24.051 13.068 24.091 ;
      RECT MASK 1 14.072 24.1225 14.252 24.1625 ;
      RECT MASK 1 20.38 24.1225 20.56 24.1625 ;
      RECT MASK 1 14.781 24.217 15.96 24.257 ;
      RECT MASK 1 16.109 24.217 17.288 24.257 ;
      RECT MASK 1 17.437 24.217 18.616 24.257 ;
      RECT MASK 1 18.765 24.217 19.944 24.257 ;
      RECT MASK 1 2.422 24.258 2.644 24.282 ;
      RECT MASK 1 0.943 24.28 1.3615 24.32 ;
      RECT MASK 1 6.056 24.332 6.116 24.562 ;
      RECT MASK 1 6.388 24.332 6.448 24.562 ;
      RECT MASK 1 6.72 24.332 6.78 24.562 ;
      RECT MASK 1 7.052 24.332 7.112 24.562 ;
      RECT MASK 1 7.384 24.332 7.444 24.562 ;
      RECT MASK 1 7.716 24.332 7.776 24.562 ;
      RECT MASK 1 8.048 24.332 8.108 24.562 ;
      RECT MASK 1 8.38 24.332 8.44 24.562 ;
      RECT MASK 1 8.712 24.332 8.772 24.562 ;
      RECT MASK 1 9.044 24.332 9.104 24.562 ;
      RECT MASK 1 9.376 24.332 9.436 24.562 ;
      RECT MASK 1 10.103 24.332 10.163 24.562 ;
      RECT MASK 1 10.767 24.332 10.827 24.562 ;
      RECT MASK 1 11.099 24.332 11.159 24.562 ;
      RECT MASK 1 11.431 24.332 11.491 24.562 ;
      RECT MASK 1 11.763 24.332 11.823 24.562 ;
      RECT MASK 1 12.095 24.332 12.155 24.562 ;
      RECT MASK 1 12.676 24.332 12.736 24.562 ;
      RECT MASK 1 13.008 24.332 13.068 24.562 ;
      RECT MASK 1 13.34 24.332 13.4 24.562 ;
      RECT MASK 1 2.422 24.348 2.874 24.372 ;
      RECT MASK 1 3.955 24.384 5.913 24.424 ;
      RECT MASK 1 13.996 24.384 20.636 24.424 ;
      RECT MASK 1 2.212 24.438 3.159 24.462 ;
      RECT MASK 1 0.984 24.44 1.4145 24.48 ;
      RECT MASK 1 2.212 24.528 3.159 24.552 ;
      RECT MASK 1 13.996 24.559 20.636 24.599 ;
      RECT MASK 1 0.943 24.6 1.465 24.64 ;
      RECT MASK 1 13.996 24.721 20.636 24.761 ;
      RECT MASK 1 2.108 24.79 3.2225 24.83 ;
      RECT MASK 1 3.948 24.79 4.566 24.83 ;
      RECT MASK 1 5.152 24.79 5.684 24.83 ;
      RECT MASK 1 13.996 24.896 20.636 24.936 ;
      RECT MASK 1 20.987 24.91 31.873 24.95 ;
      RECT MASK 1 0.825 24.94 1.583 24.98 ;
      RECT MASK 1 6.074 25 13.543 25.04 ;
      RECT MASK 1 14.781 25.063 15.96 25.103 ;
      RECT MASK 1 16.109 25.063 17.288 25.103 ;
      RECT MASK 1 17.437 25.063 18.616 25.103 ;
      RECT MASK 1 18.765 25.063 19.944 25.103 ;
      RECT MASK 1 14.072 25.1575 14.252 25.1975 ;
      RECT MASK 1 20.38 25.1575 20.56 25.1975 ;
      RECT MASK 1 14.653 25.247 15.331 25.287 ;
      RECT MASK 1 15.981 25.247 16.659 25.287 ;
      RECT MASK 1 17.309 25.247 17.987 25.287 ;
      RECT MASK 1 18.637 25.247 19.315 25.287 ;
      RECT MASK 1 6.774 25.41 6.834 26.46 ;
      RECT MASK 1 7.048 25.41 7.108 26.46 ;
      RECT MASK 1 7.322 25.41 7.382 26.46 ;
      RECT MASK 1 7.596 25.41 7.656 26.46 ;
      RECT MASK 1 7.87 25.41 7.93 26.46 ;
      RECT MASK 1 8.144 25.41 8.204 26.46 ;
      RECT MASK 1 8.418 25.41 8.478 26.46 ;
      RECT MASK 1 8.692 25.41 8.752 26.46 ;
      RECT MASK 1 8.966 25.41 9.026 26.46 ;
      RECT MASK 1 9.24 25.41 9.3 26.46 ;
      RECT MASK 1 9.514 25.41 9.574 26.46 ;
      RECT MASK 1 9.788 25.41 9.848 26.46 ;
      RECT MASK 1 10.062 25.41 10.122 26.46 ;
      RECT MASK 1 10.336 25.41 10.396 26.46 ;
      RECT MASK 1 10.61 25.41 10.67 26.46 ;
      RECT MASK 1 10.884 25.41 10.944 26.46 ;
      RECT MASK 1 11.158 25.41 11.218 26.46 ;
      RECT MASK 1 11.432 25.41 11.492 26.46 ;
      RECT MASK 1 11.706 25.41 11.766 26.46 ;
      RECT MASK 1 11.98 25.41 12.04 26.46 ;
      RECT MASK 1 12.254 25.41 12.314 26.46 ;
      RECT MASK 1 12.528 25.41 12.588 26.46 ;
      RECT MASK 1 21.849 25.41 21.909 26.46 ;
      RECT MASK 1 22.123 25.41 22.183 26.46 ;
      RECT MASK 1 22.397 25.41 22.457 26.46 ;
      RECT MASK 1 22.671 25.41 22.731 26.46 ;
      RECT MASK 1 22.945 25.41 23.005 26.46 ;
      RECT MASK 1 23.219 25.41 23.279 26.46 ;
      RECT MASK 1 23.493 25.41 23.553 26.46 ;
      RECT MASK 1 23.767 25.41 23.827 26.46 ;
      RECT MASK 1 24.041 25.41 24.101 26.46 ;
      RECT MASK 1 24.315 25.41 24.375 26.46 ;
      RECT MASK 1 24.589 25.41 24.649 26.46 ;
      RECT MASK 1 24.863 25.41 24.923 26.46 ;
      RECT MASK 1 14.653 25.473 15.331 25.513 ;
      RECT MASK 1 15.981 25.473 16.659 25.513 ;
      RECT MASK 1 17.309 25.473 17.987 25.513 ;
      RECT MASK 1 18.637 25.473 19.315 25.513 ;
      RECT MASK 1 14.072 25.5625 14.252 25.6025 ;
      RECT MASK 1 20.38 25.5625 20.56 25.6025 ;
      RECT MASK 1 14.781 25.657 15.96 25.697 ;
      RECT MASK 1 16.109 25.657 17.288 25.697 ;
      RECT MASK 1 17.437 25.657 18.616 25.697 ;
      RECT MASK 1 18.765 25.657 19.944 25.697 ;
      RECT MASK 1 13.996 25.824 20.636 25.864 ;
      RECT MASK 1 13.996 25.999 20.636 26.039 ;
      RECT MASK 1 14.107 26.32 20.525 26.36 ;
      RECT MASK 2 0.662 0.65 28.157 0.69 ;
      RECT MASK 2 29.121 0.8 31.871 0.84 ;
      RECT MASK 2 0.662 0.81 28.157 0.85 ;
      RECT MASK 2 29.121 0.96 31.871 1 ;
      RECT MASK 2 29.128 1.3 31.864 1.34 ;
      RECT MASK 2 29.128 1.46 31.864 1.5 ;
      RECT MASK 2 29.128 1.735 31.864 1.775 ;
      RECT MASK 2 29.37 1.895 29.63 1.935 ;
      RECT MASK 2 30.034 1.895 30.294 1.935 ;
      RECT MASK 2 30.698 1.895 30.958 1.935 ;
      RECT MASK 2 31.362 1.895 31.622 1.935 ;
      RECT MASK 2 29.121 2.27 31.871 2.31 ;
      RECT MASK 2 29.121 2.43 31.871 2.47 ;
      RECT MASK 2 29.121 2.69 31.871 2.73 ;
      RECT MASK 2 29.121 2.85 31.871 2.89 ;
      RECT MASK 2 29.123 3.21 31.869 3.27 ;
      RECT MASK 2 29.123 3.45 31.869 3.51 ;
      RECT MASK 2 29.123 3.69 31.869 3.75 ;
      RECT MASK 2 29.155 3.96 29.552 4.02 ;
      RECT MASK 2 29.819 3.96 30.216 4.02 ;
      RECT MASK 2 30.483 3.96 30.88 4.02 ;
      RECT MASK 2 31.147 3.96 31.505 4.02 ;
      RECT MASK 2 31.784 3.96 31.964 4.02 ;
      RECT MASK 2 29.155 4.14 29.539 4.2 ;
      RECT MASK 2 29.819 4.14 30.203 4.2 ;
      RECT MASK 2 30.483 4.14 30.867 4.2 ;
      RECT MASK 2 31.147 4.14 31.492 4.2 ;
      RECT MASK 2 31.784 4.14 31.964 4.2 ;
      RECT MASK 2 29.123 4.41 31.869 4.47 ;
      RECT MASK 2 29.123 4.65 31.869 4.71 ;
      RECT MASK 2 29.123 4.89 31.869 4.95 ;
      RECT MASK 2 29.128 5.13 31.886 5.19 ;
      RECT MASK 2 29.349 5.37 29.628 5.43 ;
      RECT MASK 2 30.013 5.37 30.292 5.43 ;
      RECT MASK 2 30.677 5.37 30.956 5.43 ;
      RECT MASK 2 31.341 5.37 31.62 5.43 ;
      RECT MASK 2 29.372 5.61 29.651 5.67 ;
      RECT MASK 2 30.036 5.61 30.315 5.67 ;
      RECT MASK 2 30.7 5.61 30.979 5.67 ;
      RECT MASK 2 31.364 5.61 31.643 5.67 ;
      RECT MASK 2 29.128 5.85 31.886 5.91 ;
      RECT MASK 2 29.121 6.11 31.871 6.15 ;
      RECT MASK 2 29.121 6.27 31.871 6.31 ;
      RECT MASK 2 29.121 6.53 31.871 6.57 ;
      RECT MASK 2 29.121 6.69 31.871 6.73 ;
      RECT MASK 2 29.128 7.05 31.864 7.11 ;
      RECT MASK 2 29.289 7.29 29.469 7.35 ;
      RECT MASK 2 29.953 7.29 30.133 7.35 ;
      RECT MASK 2 30.617 7.29 30.797 7.35 ;
      RECT MASK 2 31.281 7.29 31.461 7.35 ;
      RECT MASK 2 29.128 7.53 31.864 7.59 ;
      RECT MASK 2 29.531 7.77 29.711 7.83 ;
      RECT MASK 2 30.195 7.77 30.375 7.83 ;
      RECT MASK 2 30.859 7.77 31.039 7.83 ;
      RECT MASK 2 31.523 7.77 31.703 7.83 ;
      RECT MASK 2 29.334 8.01 29.651 8.07 ;
      RECT MASK 2 29.998 8.01 30.315 8.07 ;
      RECT MASK 2 30.662 8.01 30.979 8.07 ;
      RECT MASK 2 31.326 8.01 31.643 8.07 ;
      RECT MASK 2 29.349 8.25 29.628 8.31 ;
      RECT MASK 2 30.013 8.25 30.292 8.31 ;
      RECT MASK 2 30.677 8.25 30.956 8.31 ;
      RECT MASK 2 31.151 8.25 31.832 8.31 ;
      RECT MASK 2 29.121 8.66 31.871 8.7 ;
      RECT MASK 2 29.121 8.82 31.871 8.86 ;
      RECT MASK 2 29.121 9.08 31.871 9.12 ;
      RECT MASK 2 29.121 9.24 31.871 9.28 ;
      RECT MASK 2 29.123 9.81 31.869 9.87 ;
      RECT MASK 2 0.662 9.89 28.157 9.93 ;
      RECT MASK 2 0.662 10.05 28.157 10.09 ;
      RECT MASK 2 29.349 10.05 29.628 10.11 ;
      RECT MASK 2 30.013 10.05 30.292 10.11 ;
      RECT MASK 2 30.677 10.05 30.956 10.11 ;
      RECT MASK 2 31.198 10.05 31.454 10.11 ;
      RECT MASK 2 31.772 10.05 31.952 10.11 ;
      RECT MASK 2 0.823 10.31 10.224 10.35 ;
      RECT MASK 2 11.4715 10.31 31.871 10.35 ;
      RECT MASK 2 0.823 10.47 10.229 10.51 ;
      RECT MASK 2 11.4715 10.47 31.871 10.51 ;
      RECT MASK 2 25.791 10.71 25.851 11.76 ;
      RECT MASK 2 26.065 10.71 26.125 11.76 ;
      RECT MASK 2 26.339 10.71 26.399 11.76 ;
      RECT MASK 2 26.613 10.71 26.673 11.76 ;
      RECT MASK 2 26.887 10.71 26.947 11.76 ;
      RECT MASK 2 27.161 10.71 27.221 11.76 ;
      RECT MASK 2 8.175 10.718 9.688 10.778 ;
      RECT MASK 2 11.55 10.811 24.854 10.851 ;
      RECT MASK 2 1.634 10.928 1.694 11.152 ;
      RECT MASK 2 1.922 10.928 1.982 11.152 ;
      RECT MASK 2 2.21 10.928 2.27 11.152 ;
      RECT MASK 2 2.498 10.928 2.558 11.152 ;
      RECT MASK 2 2.786 10.928 2.846 11.152 ;
      RECT MASK 2 3.074 10.928 3.134 11.152 ;
      RECT MASK 2 3.362 10.928 3.422 11.152 ;
      RECT MASK 2 3.65 10.928 3.71 11.152 ;
      RECT MASK 2 3.938 10.928 3.998 11.152 ;
      RECT MASK 2 4.226 10.928 4.286 11.152 ;
      RECT MASK 2 4.514 10.928 4.574 11.152 ;
      RECT MASK 2 4.802 10.928 4.862 11.152 ;
      RECT MASK 2 5.09 10.928 5.15 11.152 ;
      RECT MASK 2 5.378 10.928 5.438 11.152 ;
      RECT MASK 2 5.666 10.928 5.726 11.152 ;
      RECT MASK 2 5.954 10.928 6.014 11.152 ;
      RECT MASK 2 6.242 10.928 6.302 11.152 ;
      RECT MASK 2 6.53 10.928 6.59 11.152 ;
      RECT MASK 2 6.818 10.928 6.878 11.152 ;
      RECT MASK 2 7.106 10.928 7.166 11.152 ;
      RECT MASK 2 7.394 10.928 7.454 11.152 ;
      RECT MASK 2 8.484 10.928 8.544 11.152 ;
      RECT MASK 2 8.816 10.928 8.876 11.152 ;
      RECT MASK 2 9.148 10.928 9.208 11.152 ;
      RECT MASK 2 9.48 10.928 9.54 11.152 ;
      RECT MASK 2 11.976 10.978 12.186 11.018 ;
      RECT MASK 2 12.474 10.978 12.684 11.018 ;
      RECT MASK 2 12.833 10.978 13.051 11.018 ;
      RECT MASK 2 13.165 10.978 13.383 11.018 ;
      RECT MASK 2 13.497 10.978 13.715 11.018 ;
      RECT MASK 2 13.829 10.978 14.012 11.018 ;
      RECT MASK 2 14.327 10.978 14.51 11.018 ;
      RECT MASK 2 14.964 10.978 15.174 11.018 ;
      RECT MASK 2 15.323 10.978 15.541 11.018 ;
      RECT MASK 2 15.655 10.978 15.873 11.018 ;
      RECT MASK 2 16.025 10.978 16.371 11.018 ;
      RECT MASK 2 16.689 10.978 17.035 11.018 ;
      RECT MASK 2 17.315 10.978 17.498 11.018 ;
      RECT MASK 2 17.813 10.978 18.235 11.018 ;
      RECT MASK 2 18.477 10.978 20.32 11.018 ;
      RECT MASK 2 20.469 10.978 22.312 11.018 ;
      RECT MASK 2 22.461 10.978 24.304 11.018 ;
      RECT MASK 2 11.875 11.145 12.055 11.185 ;
      RECT MASK 2 12.373 11.145 12.553 11.185 ;
      RECT MASK 2 14.863 11.145 15.043 11.185 ;
      RECT MASK 2 15.693 11.145 16.205 11.185 ;
      RECT MASK 2 16.357 11.145 16.717 11.185 ;
      RECT MASK 2 17.886 11.145 18.363 11.185 ;
      RECT MASK 2 19.214 11.145 20.355 11.185 ;
      RECT MASK 2 21.206 11.145 22.347 11.185 ;
      RECT MASK 2 23.198 11.145 24.339 11.185 ;
      RECT MASK 2 2.294 11.286 3.914 11.346 ;
      RECT MASK 2 4.31 11.286 4.49 11.346 ;
      RECT MASK 2 4.886 11.286 5.066 11.346 ;
      RECT MASK 2 5.462 11.286 5.642 11.346 ;
      RECT MASK 2 6.038 11.286 6.218 11.346 ;
      RECT MASK 2 8.597 11.29 9.427 11.35 ;
      RECT MASK 2 15.064 11.34 16.371 11.4 ;
      RECT MASK 2 11.7315 11.35 13.373 11.39 ;
      RECT MASK 2 2.294 11.514 3.914 11.574 ;
      RECT MASK 2 4.31 11.514 4.49 11.574 ;
      RECT MASK 2 4.886 11.514 5.066 11.574 ;
      RECT MASK 2 5.462 11.514 5.642 11.574 ;
      RECT MASK 2 6.038 11.514 6.218 11.574 ;
      RECT MASK 2 6.614 11.514 6.794 11.574 ;
      RECT MASK 2 8.597 11.514 9.427 11.574 ;
      RECT MASK 2 11.875 11.555 12.055 11.595 ;
      RECT MASK 2 12.373 11.555 12.553 11.595 ;
      RECT MASK 2 14.863 11.555 15.043 11.595 ;
      RECT MASK 2 15.859 11.555 16.039 11.595 ;
      RECT MASK 2 16.191 11.555 16.537 11.595 ;
      RECT MASK 2 16.689 11.555 17.035 11.595 ;
      RECT MASK 2 17.886 11.555 18.363 11.595 ;
      RECT MASK 2 19.214 11.555 20.355 11.595 ;
      RECT MASK 2 21.206 11.555 22.347 11.595 ;
      RECT MASK 2 23.198 11.555 24.339 11.595 ;
      RECT MASK 2 1.634 11.708 1.694 11.932 ;
      RECT MASK 2 1.922 11.708 1.982 11.932 ;
      RECT MASK 2 2.21 11.708 2.27 11.932 ;
      RECT MASK 2 2.498 11.708 2.558 11.932 ;
      RECT MASK 2 2.786 11.708 2.846 11.932 ;
      RECT MASK 2 3.074 11.708 3.134 11.932 ;
      RECT MASK 2 3.362 11.708 3.422 11.932 ;
      RECT MASK 2 3.65 11.708 3.71 11.932 ;
      RECT MASK 2 3.938 11.708 3.998 11.932 ;
      RECT MASK 2 4.226 11.708 4.286 11.932 ;
      RECT MASK 2 4.514 11.708 4.574 11.932 ;
      RECT MASK 2 4.802 11.708 4.862 11.932 ;
      RECT MASK 2 5.09 11.708 5.15 11.932 ;
      RECT MASK 2 5.378 11.708 5.438 11.932 ;
      RECT MASK 2 5.666 11.708 5.726 11.932 ;
      RECT MASK 2 5.954 11.708 6.014 11.932 ;
      RECT MASK 2 6.242 11.708 6.302 11.932 ;
      RECT MASK 2 6.53 11.708 6.59 11.932 ;
      RECT MASK 2 6.818 11.708 6.878 11.932 ;
      RECT MASK 2 7.106 11.708 7.166 11.932 ;
      RECT MASK 2 7.394 11.708 7.454 11.932 ;
      RECT MASK 2 8.484 11.708 8.544 11.932 ;
      RECT MASK 2 8.816 11.708 8.876 11.932 ;
      RECT MASK 2 9.148 11.708 9.208 11.932 ;
      RECT MASK 2 9.48 11.708 9.54 11.932 ;
      RECT MASK 2 11.837 11.722 12.186 11.762 ;
      RECT MASK 2 12.335 11.722 12.684 11.762 ;
      RECT MASK 2 12.833 11.722 13.051 11.762 ;
      RECT MASK 2 13.165 11.722 13.383 11.762 ;
      RECT MASK 2 13.497 11.722 13.715 11.762 ;
      RECT MASK 2 13.829 11.722 14.012 11.762 ;
      RECT MASK 2 14.327 11.722 14.51 11.762 ;
      RECT MASK 2 14.825 11.722 15.174 11.762 ;
      RECT MASK 2 15.323 11.722 15.541 11.762 ;
      RECT MASK 2 15.655 11.722 15.873 11.762 ;
      RECT MASK 2 16.025 11.722 16.369 11.762 ;
      RECT MASK 2 16.807 11.722 17.035 11.762 ;
      RECT MASK 2 17.315 11.722 17.498 11.762 ;
      RECT MASK 2 17.813 11.722 18.235 11.762 ;
      RECT MASK 2 18.477 11.722 20.32 11.762 ;
      RECT MASK 2 20.469 11.722 22.312 11.762 ;
      RECT MASK 2 22.461 11.722 24.304 11.762 ;
      RECT MASK 2 11.55 11.889 24.498 11.929 ;
      RECT MASK 2 24.969 11.99 28.067 12.03 ;
      RECT MASK 2 24.969 12.15 28.067 12.19 ;
      RECT MASK 2 11.4715 12.23 24.451 12.27 ;
      RECT MASK 2 0.759 12.35 10.293 12.39 ;
      RECT MASK 2 11.4715 12.39 24.451 12.43 ;
      RECT MASK 2 0.759 12.51 10.293 12.55 ;
      RECT MASK 2 20.987 12.65 31.832 12.69 ;
      RECT MASK 2 0.759 12.77 10.293 12.81 ;
      RECT MASK 2 20.987 12.81 31.832 12.85 ;
      RECT MASK 2 0.759 12.93 10.293 12.97 ;
      RECT MASK 2 21.739 13.07 24.993 13.11 ;
      RECT MASK 2 21.822 13.27 24.91 13.31 ;
      RECT MASK 2 12.343 13.28 15.579 13.32 ;
      RECT MASK 2 15.885 13.28 16.659 13.32 ;
      RECT MASK 2 16.964 13.368 19.743 13.392 ;
      RECT MASK 2 1.634 13.388 1.694 13.612 ;
      RECT MASK 2 1.922 13.388 1.982 13.612 ;
      RECT MASK 2 2.21 13.388 2.27 13.612 ;
      RECT MASK 2 2.498 13.388 2.558 13.612 ;
      RECT MASK 2 2.786 13.388 2.846 13.612 ;
      RECT MASK 2 3.074 13.388 3.134 13.612 ;
      RECT MASK 2 3.362 13.388 3.422 13.612 ;
      RECT MASK 2 3.65 13.388 3.71 13.612 ;
      RECT MASK 2 3.938 13.388 3.998 13.612 ;
      RECT MASK 2 4.226 13.388 4.286 13.612 ;
      RECT MASK 2 4.514 13.388 4.574 13.612 ;
      RECT MASK 2 4.802 13.388 4.862 13.612 ;
      RECT MASK 2 5.09 13.388 5.15 13.612 ;
      RECT MASK 2 5.378 13.388 5.438 13.612 ;
      RECT MASK 2 5.666 13.388 5.726 13.612 ;
      RECT MASK 2 5.954 13.388 6.014 13.612 ;
      RECT MASK 2 6.242 13.388 6.302 13.612 ;
      RECT MASK 2 6.53 13.388 6.59 13.612 ;
      RECT MASK 2 6.818 13.388 6.878 13.612 ;
      RECT MASK 2 7.106 13.388 7.166 13.612 ;
      RECT MASK 2 7.394 13.388 7.454 13.612 ;
      RECT MASK 2 8.484 13.388 8.544 13.612 ;
      RECT MASK 2 8.816 13.388 8.876 13.612 ;
      RECT MASK 2 9.148 13.388 9.208 13.612 ;
      RECT MASK 2 9.48 13.388 9.54 13.612 ;
      RECT MASK 2 12.343 13.44 15.579 13.48 ;
      RECT MASK 2 15.885 13.44 16.659 13.48 ;
      RECT MASK 2 21.485 13.47 23.582 13.51 ;
      RECT MASK 2 16.964 13.578 19.876 13.602 ;
      RECT MASK 2 12.343 13.678 15.614 13.718 ;
      RECT MASK 2 15.885 13.678 16.717 13.718 ;
      RECT MASK 2 1.43 13.756 3.338 13.816 ;
      RECT MASK 2 5.174 13.756 5.354 13.816 ;
      RECT MASK 2 6.326 13.756 7.658 13.816 ;
      RECT MASK 2 8.597 13.756 9.427 13.816 ;
      RECT MASK 2 21.573 13.77 21.761 13.81 ;
      RECT MASK 2 21.905 13.77 24.827 13.81 ;
      RECT MASK 2 24.971 13.77 25.159 13.81 ;
      RECT MASK 2 17.173 13.822 19.876 13.846 ;
      RECT MASK 2 12.7 13.838 12.76 14.088 ;
      RECT MASK 2 14.268 13.838 14.328 14.068 ;
      RECT MASK 2 14.6 13.838 14.66 14.068 ;
      RECT MASK 2 16.076 13.838 16.136 14.0485 ;
      RECT MASK 2 16.408 13.838 16.468 14.0485 ;
      RECT MASK 2 1.43 13.964 2.762 14.024 ;
      RECT MASK 2 3.158 13.964 3.338 14.024 ;
      RECT MASK 2 5.174 13.964 5.354 14.024 ;
      RECT MASK 2 6.326 13.964 6.506 14.024 ;
      RECT MASK 2 6.902 13.964 7.658 14.024 ;
      RECT MASK 2 8.597 13.964 9.427 14.024 ;
      RECT MASK 2 22.149 13.97 24.744 14.01 ;
      RECT MASK 2 17.864 13.987 19.876 14.011 ;
      RECT MASK 2 13.304 14.0125 13.484 14.0525 ;
      RECT MASK 2 15.278 14.0125 15.458 14.0525 ;
      RECT MASK 2 17.864 14.077 19.876 14.101 ;
      RECT MASK 2 1.634 14.168 1.694 14.392 ;
      RECT MASK 2 1.922 14.168 1.982 14.392 ;
      RECT MASK 2 2.21 14.168 2.27 14.392 ;
      RECT MASK 2 2.498 14.168 2.558 14.392 ;
      RECT MASK 2 2.786 14.168 2.846 14.392 ;
      RECT MASK 2 3.074 14.168 3.134 14.392 ;
      RECT MASK 2 3.362 14.168 3.422 14.392 ;
      RECT MASK 2 3.65 14.168 3.71 14.392 ;
      RECT MASK 2 3.938 14.168 3.998 14.392 ;
      RECT MASK 2 4.226 14.168 4.286 14.392 ;
      RECT MASK 2 4.514 14.168 4.574 14.392 ;
      RECT MASK 2 4.802 14.168 4.862 14.392 ;
      RECT MASK 2 5.09 14.168 5.15 14.392 ;
      RECT MASK 2 5.378 14.168 5.438 14.392 ;
      RECT MASK 2 5.666 14.168 5.726 14.392 ;
      RECT MASK 2 5.954 14.168 6.014 14.392 ;
      RECT MASK 2 6.242 14.168 6.302 14.392 ;
      RECT MASK 2 6.53 14.168 6.59 14.392 ;
      RECT MASK 2 6.818 14.168 6.878 14.392 ;
      RECT MASK 2 7.106 14.168 7.166 14.392 ;
      RECT MASK 2 7.394 14.168 7.454 14.392 ;
      RECT MASK 2 8.484 14.168 8.544 14.392 ;
      RECT MASK 2 8.816 14.168 8.876 14.392 ;
      RECT MASK 2 9.148 14.168 9.208 14.392 ;
      RECT MASK 2 9.48 14.168 9.54 14.392 ;
      RECT MASK 2 21.651 14.17 22.088 14.21 ;
      RECT MASK 2 22.647 14.17 24.085 14.21 ;
      RECT MASK 2 24.312 14.17 25.081 14.21 ;
      RECT MASK 2 12.343 14.208 12.692 14.248 ;
      RECT MASK 2 12.841 14.208 16.566 14.248 ;
      RECT MASK 2 17.864 14.253 19.876 14.277 ;
      RECT MASK 2 17.864 14.343 19.876 14.367 ;
      RECT MASK 2 14.077 14.41 14.757 14.45 ;
      RECT MASK 2 17.864 14.433 19.876 14.457 ;
      RECT MASK 2 17.188 14.523 19.876 14.547 ;
      RECT MASK 2 21.651 14.57 22.088 14.61 ;
      RECT MASK 2 22.647 14.57 24.085 14.61 ;
      RECT MASK 2 24.312 14.57 25.081 14.61 ;
      RECT MASK 2 12.509 14.612 16.566 14.652 ;
      RECT MASK 2 17.32 14.613 19.876 14.637 ;
      RECT MASK 2 17.32 14.703 19.876 14.727 ;
      RECT MASK 2 22.149 14.77 24.744 14.81 ;
      RECT MASK 2 12.7 14.772 12.76 15.022 ;
      RECT MASK 2 14.268 14.792 14.328 15.022 ;
      RECT MASK 2 14.6 14.792 14.66 15.022 ;
      RECT MASK 2 17.32 14.793 19.876 14.817 ;
      RECT MASK 2 13.304 14.8075 13.484 14.8475 ;
      RECT MASK 2 15.278 14.8075 15.458 14.8475 ;
      RECT MASK 2 0.823 14.81 10.293 14.85 ;
      RECT MASK 2 16.076 14.811 16.136 15.022 ;
      RECT MASK 2 16.408 14.811 16.468 15.022 ;
      RECT MASK 2 17.6005 14.883 19.876 14.907 ;
      RECT MASK 2 0.823 14.97 10.293 15.01 ;
      RECT MASK 2 21.573 14.97 21.761 15.01 ;
      RECT MASK 2 21.905 14.97 24.827 15.01 ;
      RECT MASK 2 24.971 14.97 25.159 15.01 ;
      RECT MASK 2 17.6005 15.056 19.876 15.08 ;
      RECT MASK 2 12.343 15.142 13.484 15.182 ;
      RECT MASK 2 13.911 15.142 14.851 15.182 ;
      RECT MASK 2 15.278 15.142 17.323 15.182 ;
      RECT MASK 2 21.573 15.18 21.761 15.22 ;
      RECT MASK 2 21.905 15.18 24.827 15.22 ;
      RECT MASK 2 24.971 15.18 25.159 15.22 ;
      RECT MASK 2 0.825 15.35 1.583 15.39 ;
      RECT MASK 2 12.343 15.358 13.484 15.398 ;
      RECT MASK 2 13.911 15.358 14.851 15.398 ;
      RECT MASK 2 15.278 15.358 17.323 15.398 ;
      RECT MASK 2 2.123 15.371 10.518 15.411 ;
      RECT MASK 2 22.149 15.38 24.744 15.42 ;
      RECT MASK 2 17.6005 15.46 19.876 15.484 ;
      RECT MASK 2 0.825 15.51 1.583 15.55 ;
      RECT MASK 2 12.7 15.518 12.76 15.768 ;
      RECT MASK 2 14.268 15.518 14.328 15.748 ;
      RECT MASK 2 14.6 15.518 14.66 15.748 ;
      RECT MASK 2 16.076 15.518 16.136 15.729 ;
      RECT MASK 2 16.408 15.518 16.468 15.729 ;
      RECT MASK 2 2.123 15.549 10.518 15.589 ;
      RECT MASK 2 21.651 15.58 22.088 15.62 ;
      RECT MASK 2 22.647 15.58 24.085 15.62 ;
      RECT MASK 2 24.312 15.58 25.081 15.62 ;
      RECT MASK 2 17.6005 15.633 19.876 15.657 ;
      RECT MASK 2 13.304 15.6925 13.484 15.7325 ;
      RECT MASK 2 15.278 15.6925 15.458 15.7325 ;
      RECT MASK 2 17.32 15.723 19.876 15.747 ;
      RECT MASK 2 1.053 15.75 1.332 15.81 ;
      RECT MASK 2 1.484 15.75 1.664 15.81 ;
      RECT MASK 2 17.32 15.813 19.876 15.837 ;
      RECT MASK 2 12.509 15.888 16.566 15.928 ;
      RECT MASK 2 21.573 15.89 22.005 15.93 ;
      RECT MASK 2 22.237 15.89 22.757 15.93 ;
      RECT MASK 2 22.901 15.89 25.159 15.93 ;
      RECT MASK 2 17.32 15.903 19.876 15.927 ;
      RECT MASK 2 2.855 15.96 2.915 17.01 ;
      RECT MASK 2 3.129 15.96 3.189 17.01 ;
      RECT MASK 2 3.403 15.96 3.463 17.01 ;
      RECT MASK 2 3.677 15.96 3.737 17.01 ;
      RECT MASK 2 3.951 15.96 4.011 17.01 ;
      RECT MASK 2 4.225 15.96 4.285 17.01 ;
      RECT MASK 2 4.499 15.96 4.559 17.01 ;
      RECT MASK 2 4.773 15.96 4.833 17.01 ;
      RECT MASK 2 5.047 15.96 5.107 17.01 ;
      RECT MASK 2 5.321 15.96 5.381 17.01 ;
      RECT MASK 2 5.595 15.96 5.655 17.01 ;
      RECT MASK 2 5.869 15.96 5.929 17.01 ;
      RECT MASK 2 6.143 15.96 6.203 17.01 ;
      RECT MASK 2 6.417 15.96 6.477 17.01 ;
      RECT MASK 2 6.691 15.96 6.751 17.01 ;
      RECT MASK 2 6.965 15.96 7.025 17.01 ;
      RECT MASK 2 7.239 15.96 7.299 17.01 ;
      RECT MASK 2 7.513 15.96 7.573 17.01 ;
      RECT MASK 2 7.787 15.96 7.847 17.01 ;
      RECT MASK 2 8.061 15.96 8.121 17.01 ;
      RECT MASK 2 8.335 15.96 8.395 17.01 ;
      RECT MASK 2 8.609 15.96 8.669 17.01 ;
      RECT MASK 2 8.883 15.96 8.943 17.01 ;
      RECT MASK 2 9.157 15.96 9.217 17.01 ;
      RECT MASK 2 9.431 15.96 9.491 17.01 ;
      RECT MASK 2 9.705 15.96 9.765 17.01 ;
      RECT MASK 2 9.979 15.96 10.039 17.01 ;
      RECT MASK 2 10.253 15.96 10.313 17.01 ;
      RECT MASK 2 0.827 15.99 1.581 16.05 ;
      RECT MASK 2 17.188 15.993 19.876 16.017 ;
      RECT MASK 2 2.118 16.025 2.238 16.105 ;
      RECT MASK 2 17.864 16.083 19.876 16.107 ;
      RECT MASK 2 14.077 16.09 14.757 16.13 ;
      RECT MASK 2 21.651 16.09 25.081 16.13 ;
      RECT MASK 2 17.864 16.173 19.876 16.197 ;
      RECT MASK 2 17.864 16.263 19.876 16.287 ;
      RECT MASK 2 2.118 16.265 2.238 16.345 ;
      RECT MASK 2 12.343 16.292 12.692 16.332 ;
      RECT MASK 2 12.841 16.292 16.566 16.332 ;
      RECT MASK 2 21.485 16.39 21.839 16.43 ;
      RECT MASK 2 22.735 16.39 22.923 16.43 ;
      RECT MASK 2 17.864 16.439 19.876 16.463 ;
      RECT MASK 2 12.7 16.452 12.76 16.702 ;
      RECT MASK 2 14.268 16.472 14.328 16.702 ;
      RECT MASK 2 14.6 16.472 14.66 16.702 ;
      RECT MASK 2 13.304 16.4875 13.484 16.5275 ;
      RECT MASK 2 15.278 16.4875 15.458 16.5275 ;
      RECT MASK 2 16.076 16.4915 16.136 16.702 ;
      RECT MASK 2 16.408 16.4915 16.468 16.702 ;
      RECT MASK 2 17.864 16.529 19.876 16.553 ;
      RECT MASK 2 0.825 16.58 1.583 16.62 ;
      RECT MASK 2 2.118 16.625 2.238 16.705 ;
      RECT MASK 2 21.485 16.64 21.839 16.68 ;
      RECT MASK 2 22.071 16.64 22.259 16.68 ;
      RECT MASK 2 22.403 16.64 22.591 16.68 ;
      RECT MASK 2 22.735 16.64 22.923 16.68 ;
      RECT MASK 2 17.173 16.694 19.876 16.718 ;
      RECT MASK 2 0.825 16.74 1.583 16.78 ;
      RECT MASK 2 12.343 16.822 15.614 16.862 ;
      RECT MASK 2 15.885 16.822 16.717 16.862 ;
      RECT MASK 2 21.817 16.84 22.259 16.88 ;
      RECT MASK 2 22.486 16.84 23.089 16.88 ;
      RECT MASK 2 2.118 16.865 2.238 16.945 ;
      RECT MASK 2 16.964 16.938 19.876 16.962 ;
      RECT MASK 2 0.825 17 1.583 17.04 ;
      RECT MASK 2 21.948 17.04 22.128 17.08 ;
      RECT MASK 2 22.28 17.04 22.46 17.08 ;
      RECT MASK 2 22.743 17.04 22.923 17.08 ;
      RECT MASK 2 23.11 17.04 23.29 17.08 ;
      RECT MASK 2 12.343 17.06 15.579 17.1 ;
      RECT MASK 2 15.885 17.06 16.659 17.1 ;
      RECT MASK 2 16.964 17.148 19.743 17.172 ;
      RECT MASK 2 0.825 17.16 1.583 17.2 ;
      RECT MASK 2 12.343 17.22 15.579 17.26 ;
      RECT MASK 2 15.885 17.22 16.659 17.26 ;
      RECT MASK 2 21.651 17.39 25.081 17.43 ;
      RECT MASK 2 1.053 17.55 1.332 17.61 ;
      RECT MASK 2 2.855 17.55 2.915 18.6 ;
      RECT MASK 2 3.129 17.55 3.189 18.6 ;
      RECT MASK 2 3.403 17.55 3.463 18.6 ;
      RECT MASK 2 3.677 17.55 3.737 18.6 ;
      RECT MASK 2 3.951 17.55 4.011 18.6 ;
      RECT MASK 2 4.225 17.55 4.285 18.6 ;
      RECT MASK 2 4.499 17.55 4.559 18.6 ;
      RECT MASK 2 4.773 17.55 4.833 18.6 ;
      RECT MASK 2 5.047 17.55 5.107 18.6 ;
      RECT MASK 2 5.321 17.55 5.381 18.6 ;
      RECT MASK 2 5.595 17.55 5.655 18.6 ;
      RECT MASK 2 5.869 17.55 5.929 18.6 ;
      RECT MASK 2 6.143 17.55 6.203 18.6 ;
      RECT MASK 2 21.651 17.55 25.081 17.59 ;
      RECT MASK 2 2.118 17.615 2.238 17.695 ;
      RECT MASK 2 1.038 17.79 1.355 17.85 ;
      RECT MASK 2 21.905 17.81 23.333 17.85 ;
      RECT MASK 2 2.118 17.855 2.238 17.935 ;
      RECT MASK 2 21.988 18.01 23.582 18.05 ;
      RECT MASK 2 1.235 18.03 1.415 18.09 ;
      RECT MASK 2 7.195 18.08 20.215 18.12 ;
      RECT MASK 2 2.118 18.215 2.238 18.295 ;
      RECT MASK 2 7.195 18.24 20.215 18.28 ;
      RECT MASK 2 0.832 18.27 1.576 18.33 ;
      RECT MASK 2 2.118 18.455 2.238 18.535 ;
      RECT MASK 2 0.993 18.51 1.173 18.57 ;
      RECT MASK 2 7.148 18.571 20.262 18.611 ;
      RECT MASK 2 9.427 18.731 20.151 18.771 ;
      RECT MASK 2 7.574 18.748 7.784 18.788 ;
      RECT MASK 2 8.072 18.748 8.282 18.788 ;
      RECT MASK 2 8.57 18.748 8.78 18.788 ;
      RECT MASK 2 9.095 18.748 9.313 18.788 ;
      RECT MASK 2 0.832 18.75 1.576 18.81 ;
      RECT MASK 2 21.988 18.86 24.251 18.9 ;
      RECT MASK 2 7.473 18.915 7.653 18.955 ;
      RECT MASK 2 7.971 18.915 8.151 18.955 ;
      RECT MASK 2 8.469 18.915 8.649 18.955 ;
      RECT MASK 2 9.915 18.915 10.817 18.955 ;
      RECT MASK 2 11.243 18.915 12.145 18.955 ;
      RECT MASK 2 12.571 18.915 13.473 18.955 ;
      RECT MASK 2 13.899 18.915 14.801 18.955 ;
      RECT MASK 2 15.227 18.915 16.129 18.955 ;
      RECT MASK 2 16.555 18.915 17.457 18.955 ;
      RECT MASK 2 17.883 18.915 18.785 18.955 ;
      RECT MASK 2 19.211 18.915 20.113 18.955 ;
      RECT MASK 2 5.322 19.06 6.522 19.08 ;
      RECT MASK 2 21.905 19.06 23.333 19.1 ;
      RECT MASK 2 23.477 19.06 23.665 19.1 ;
      RECT MASK 2 0.825 19.13 1.583 19.17 ;
      RECT MASK 2 2.855 19.14 2.915 20.19 ;
      RECT MASK 2 3.129 19.14 3.189 20.19 ;
      RECT MASK 2 3.403 19.14 3.463 20.19 ;
      RECT MASK 2 3.677 19.14 3.737 20.19 ;
      RECT MASK 2 3.951 19.14 4.011 20.19 ;
      RECT MASK 2 4.225 19.14 4.285 20.19 ;
      RECT MASK 2 2.118 19.205 2.238 19.285 ;
      RECT MASK 2 21.905 19.24 23.831 19.28 ;
      RECT MASK 2 0.825 19.29 1.583 19.33 ;
      RECT MASK 2 7.473 19.325 7.653 19.365 ;
      RECT MASK 2 7.971 19.325 8.151 19.365 ;
      RECT MASK 2 8.469 19.325 8.649 19.365 ;
      RECT MASK 2 9.915 19.325 10.817 19.365 ;
      RECT MASK 2 11.243 19.325 12.145 19.365 ;
      RECT MASK 2 12.571 19.325 13.473 19.365 ;
      RECT MASK 2 13.899 19.325 14.801 19.365 ;
      RECT MASK 2 15.227 19.325 16.129 19.365 ;
      RECT MASK 2 16.555 19.325 17.457 19.365 ;
      RECT MASK 2 17.883 19.325 18.785 19.365 ;
      RECT MASK 2 19.211 19.325 20.113 19.365 ;
      RECT MASK 2 5.322 19.38 6.522 19.4 ;
      RECT MASK 2 21.988 19.44 24.251 19.48 ;
      RECT MASK 2 2.118 19.445 2.238 19.525 ;
      RECT MASK 2 5.322 19.46 6.522 19.48 ;
      RECT MASK 2 7.435 19.492 7.784 19.532 ;
      RECT MASK 2 7.933 19.492 8.282 19.532 ;
      RECT MASK 2 8.431 19.492 8.78 19.532 ;
      RECT MASK 2 8.967 19.492 9.185 19.532 ;
      RECT MASK 2 9.427 19.509 20.151 19.549 ;
      RECT MASK 2 5.322 19.54 6.522 19.56 ;
      RECT MASK 2 0.825 19.55 1.583 19.59 ;
      RECT MASK 2 5.322 19.62 6.522 19.64 ;
      RECT MASK 2 7.148 19.669 20.359 19.709 ;
      RECT MASK 2 5.322 19.7 6.522 19.72 ;
      RECT MASK 2 0.825 19.71 1.583 19.75 ;
      RECT MASK 2 5.322 19.78 6.522 19.8 ;
      RECT MASK 2 2.118 19.805 2.238 19.885 ;
      RECT MASK 2 0.832 19.95 1.598 20.01 ;
      RECT MASK 2 7.195 20 20.359 20.04 ;
      RECT MASK 2 21.573 20 21.839 20.04 ;
      RECT MASK 2 22.071 20 23.665 20.04 ;
      RECT MASK 2 23.809 20 23.997 20.04 ;
      RECT MASK 2 2.118 20.045 2.238 20.125 ;
      RECT MASK 2 5.322 20.1 6.522 20.12 ;
      RECT MASK 2 7.195 20.16 20.359 20.2 ;
      RECT MASK 2 1.076 20.19 1.355 20.25 ;
      RECT MASK 2 21.651 20.2 23.919 20.24 ;
      RECT MASK 2 1.053 20.43 1.332 20.49 ;
      RECT MASK 2 13.996 20.501 20.636 20.541 ;
      RECT MASK 2 14.947 20.668 15.13 20.708 ;
      RECT MASK 2 15.445 20.668 15.867 20.708 ;
      RECT MASK 2 16.109 20.668 17.288 20.708 ;
      RECT MASK 2 17.437 20.668 18.616 20.708 ;
      RECT MASK 2 18.765 20.668 19.944 20.708 ;
      RECT MASK 2 0.832 20.67 1.598 20.73 ;
      RECT MASK 2 6.074 20.72 13.543 20.76 ;
      RECT MASK 2 21.651 20.75 25.081 20.79 ;
      RECT MASK 2 14.072 20.7625 14.252 20.8025 ;
      RECT MASK 2 20.38 20.7625 20.56 20.8025 ;
      RECT MASK 2 15.518 20.835 15.995 20.875 ;
      RECT MASK 2 16.479 20.835 17.323 20.875 ;
      RECT MASK 2 17.759 20.835 18.651 20.875 ;
      RECT MASK 2 19.087 20.835 19.979 20.875 ;
      RECT MASK 2 6.074 20.88 13.543 20.92 ;
      RECT MASK 2 0.827 20.91 1.581 20.97 ;
      RECT MASK 2 21.651 20.91 25.081 20.95 ;
      RECT MASK 2 3.948 20.93 4.566 20.97 ;
      RECT MASK 2 5.152 20.93 5.684 20.97 ;
      RECT MASK 2 3.948 21.09 4.566 21.13 ;
      RECT MASK 2 5.152 21.09 5.684 21.13 ;
      RECT MASK 2 5.87 21.118 13.543 21.158 ;
      RECT MASK 2 0.827 21.15 1.581 21.21 ;
      RECT MASK 2 2.212 21.243 3.159 21.267 ;
      RECT MASK 2 15.518 21.245 15.995 21.285 ;
      RECT MASK 2 16.479 21.245 17.323 21.285 ;
      RECT MASK 2 17.759 21.245 18.651 21.285 ;
      RECT MASK 2 19.087 21.245 19.979 21.285 ;
      RECT MASK 2 6.222 21.278 6.282 21.508 ;
      RECT MASK 2 6.554 21.278 6.614 21.508 ;
      RECT MASK 2 6.886 21.278 6.946 21.508 ;
      RECT MASK 2 7.218 21.278 7.278 21.508 ;
      RECT MASK 2 7.55 21.278 7.61 21.508 ;
      RECT MASK 2 7.882 21.278 7.942 21.508 ;
      RECT MASK 2 8.214 21.278 8.274 21.508 ;
      RECT MASK 2 8.546 21.278 8.606 21.508 ;
      RECT MASK 2 8.878 21.278 8.938 21.508 ;
      RECT MASK 2 9.21 21.278 9.27 21.508 ;
      RECT MASK 2 9.542 21.278 9.602 21.508 ;
      RECT MASK 2 10.269 21.278 10.329 21.508 ;
      RECT MASK 2 10.601 21.278 10.661 21.508 ;
      RECT MASK 2 11.265 21.278 11.325 21.508 ;
      RECT MASK 2 11.597 21.278 11.657 21.508 ;
      RECT MASK 2 11.929 21.278 11.989 21.508 ;
      RECT MASK 2 12.51 21.278 12.57 21.508 ;
      RECT MASK 2 12.842 21.278 12.902 21.508 ;
      RECT MASK 2 13.174 21.278 13.234 21.508 ;
      RECT MASK 2 14.072 21.3175 14.252 21.3575 ;
      RECT MASK 2 20.38 21.3175 20.56 21.3575 ;
      RECT MASK 2 3.898 21.321 5.936 21.361 ;
      RECT MASK 2 2.422 21.333 2.874 21.357 ;
      RECT MASK 2 0.827 21.39 1.581 21.45 ;
      RECT MASK 2 14.947 21.412 15.13 21.452 ;
      RECT MASK 2 15.445 21.412 15.867 21.452 ;
      RECT MASK 2 16.109 21.412 17.288 21.452 ;
      RECT MASK 2 17.437 21.412 18.616 21.452 ;
      RECT MASK 2 18.765 21.412 19.944 21.452 ;
      RECT MASK 2 2.422 21.423 2.874 21.447 ;
      RECT MASK 2 2.212 21.513 3.159 21.537 ;
      RECT MASK 2 13.996 21.579 20.636 21.619 ;
      RECT MASK 2 4.104 21.602 4.164 21.832 ;
      RECT MASK 2 5.33 21.602 5.39 21.832 ;
      RECT MASK 2 9.268 21.648 9.579 21.688 ;
      RECT MASK 2 10.126 21.648 10.804 21.688 ;
      RECT MASK 2 11.982 21.648 12.3 21.688 ;
      RECT MASK 2 12.485 21.648 12.927 21.688 ;
      RECT MASK 2 13.061 21.648 13.425 21.688 ;
      RECT MASK 2 0.859 21.66 1.243 21.72 ;
      RECT MASK 2 1.496 21.66 1.676 21.72 ;
      RECT MASK 2 0.859 21.84 1.256 21.9 ;
      RECT MASK 2 1.496 21.84 1.676 21.9 ;
      RECT MASK 2 5.761 21.85 13.508 21.89 ;
      RECT MASK 2 22.46 21.93 24.26 21.95 ;
      RECT MASK 2 13.996 21.941 20.636 21.981 ;
      RECT MASK 2 22.46 22.01 24.26 22.03 ;
      RECT MASK 2 6.079 22.052 6.307 22.092 ;
      RECT MASK 2 9.912 22.052 10.472 22.092 ;
      RECT MASK 2 10.79 22.052 11.018 22.092 ;
      RECT MASK 2 11.738 22.052 11.966 22.092 ;
      RECT MASK 2 12.319 22.052 13.068 22.092 ;
      RECT MASK 2 14.781 22.108 15.203 22.148 ;
      RECT MASK 2 15.445 22.108 15.867 22.148 ;
      RECT MASK 2 16.109 22.108 17.288 22.148 ;
      RECT MASK 2 17.437 22.108 18.616 22.148 ;
      RECT MASK 2 18.765 22.108 19.944 22.148 ;
      RECT MASK 2 0.827 22.11 1.581 22.17 ;
      RECT MASK 2 2.625 22.158 2.874 22.182 ;
      RECT MASK 2 3.955 22.168 5.936 22.208 ;
      RECT MASK 2 14.072 22.2025 14.252 22.2425 ;
      RECT MASK 2 20.38 22.2025 20.56 22.2425 ;
      RECT MASK 2 6.222 22.232 6.282 22.462 ;
      RECT MASK 2 6.554 22.232 6.614 22.462 ;
      RECT MASK 2 6.886 22.232 6.946 22.462 ;
      RECT MASK 2 7.218 22.232 7.278 22.462 ;
      RECT MASK 2 7.55 22.232 7.61 22.462 ;
      RECT MASK 2 7.882 22.232 7.942 22.462 ;
      RECT MASK 2 8.214 22.232 8.274 22.462 ;
      RECT MASK 2 8.546 22.232 8.606 22.462 ;
      RECT MASK 2 8.878 22.232 8.938 22.462 ;
      RECT MASK 2 9.21 22.232 9.27 22.462 ;
      RECT MASK 2 9.542 22.232 9.602 22.462 ;
      RECT MASK 2 10.269 22.232 10.329 22.462 ;
      RECT MASK 2 11.265 22.232 11.325 22.462 ;
      RECT MASK 2 11.597 22.232 11.657 22.462 ;
      RECT MASK 2 11.929 22.232 11.989 22.462 ;
      RECT MASK 2 12.51 22.232 12.57 22.462 ;
      RECT MASK 2 12.842 22.232 12.902 22.462 ;
      RECT MASK 2 13.174 22.232 13.234 22.462 ;
      RECT MASK 2 2.422 22.248 2.874 22.272 ;
      RECT MASK 2 14.854 22.275 15.331 22.315 ;
      RECT MASK 2 15.518 22.275 15.995 22.315 ;
      RECT MASK 2 16.479 22.275 17.323 22.315 ;
      RECT MASK 2 17.759 22.275 18.651 22.315 ;
      RECT MASK 2 19.087 22.275 19.979 22.315 ;
      RECT MASK 2 4.104 22.328 4.164 22.558 ;
      RECT MASK 2 5.33 22.328 5.39 22.558 ;
      RECT MASK 2 2.136 22.338 3.159 22.362 ;
      RECT MASK 2 0.827 22.35 1.581 22.41 ;
      RECT MASK 2 2.136 22.428 3.159 22.452 ;
      RECT MASK 2 4.647 22.43 4.707 22.57 ;
      RECT MASK 2 4.979 22.43 5.039 22.57 ;
      RECT MASK 2 22.46 22.49 23.455 22.51 ;
      RECT MASK 2 5.913 22.582 9.745 22.622 ;
      RECT MASK 2 9.944 22.582 13.543 22.622 ;
      RECT MASK 2 0.827 22.59 1.581 22.65 ;
      RECT MASK 2 14.854 22.685 15.331 22.725 ;
      RECT MASK 2 15.518 22.685 15.995 22.725 ;
      RECT MASK 2 16.479 22.685 17.323 22.725 ;
      RECT MASK 2 17.759 22.685 18.651 22.725 ;
      RECT MASK 2 19.087 22.685 19.979 22.725 ;
      RECT MASK 2 2.0735 22.69 3.2225 22.73 ;
      RECT MASK 2 14.072 22.7575 14.252 22.7975 ;
      RECT MASK 2 20.38 22.7575 20.56 22.7975 ;
      RECT MASK 2 6.046 22.82 9.626 22.86 ;
      RECT MASK 2 10.081 22.82 13.543 22.86 ;
      RECT MASK 2 14.781 22.852 15.203 22.892 ;
      RECT MASK 2 15.445 22.852 15.867 22.892 ;
      RECT MASK 2 16.109 22.852 17.288 22.892 ;
      RECT MASK 2 17.437 22.852 18.616 22.892 ;
      RECT MASK 2 18.765 22.852 19.944 22.892 ;
      RECT MASK 2 0.825 22.97 1.583 23.01 ;
      RECT MASK 2 6.046 22.98 9.626 23.02 ;
      RECT MASK 2 10.081 22.98 13.543 23.02 ;
      RECT MASK 2 13.996 23.019 20.636 23.059 ;
      RECT MASK 2 22.46 23.03 24.26 23.05 ;
      RECT MASK 2 2.0735 23.11 3.2225 23.15 ;
      RECT MASK 2 22.46 23.11 24.26 23.13 ;
      RECT MASK 2 0.825 23.13 1.583 23.17 ;
      RECT MASK 2 5.913 23.218 9.745 23.258 ;
      RECT MASK 2 9.944 23.218 13.543 23.258 ;
      RECT MASK 2 4.647 23.27 4.707 23.41 ;
      RECT MASK 2 4.979 23.27 5.039 23.41 ;
      RECT MASK 2 22.4895 23.27 23.321 23.29 ;
      RECT MASK 2 23.905 23.27 24.2605 23.29 ;
      RECT MASK 2 4.104 23.282 4.164 23.512 ;
      RECT MASK 2 5.33 23.282 5.39 23.512 ;
      RECT MASK 2 6.222 23.378 6.282 23.608 ;
      RECT MASK 2 6.554 23.378 6.614 23.608 ;
      RECT MASK 2 6.886 23.378 6.946 23.608 ;
      RECT MASK 2 7.218 23.378 7.278 23.608 ;
      RECT MASK 2 7.55 23.378 7.61 23.608 ;
      RECT MASK 2 7.882 23.378 7.942 23.608 ;
      RECT MASK 2 8.214 23.378 8.274 23.608 ;
      RECT MASK 2 8.546 23.378 8.606 23.608 ;
      RECT MASK 2 8.878 23.378 8.938 23.608 ;
      RECT MASK 2 9.21 23.378 9.27 23.608 ;
      RECT MASK 2 9.542 23.378 9.602 23.608 ;
      RECT MASK 2 10.269 23.378 10.329 23.608 ;
      RECT MASK 2 11.265 23.378 11.325 23.608 ;
      RECT MASK 2 11.597 23.378 11.657 23.608 ;
      RECT MASK 2 11.929 23.378 11.989 23.608 ;
      RECT MASK 2 12.51 23.378 12.57 23.608 ;
      RECT MASK 2 12.842 23.378 12.902 23.608 ;
      RECT MASK 2 13.174 23.378 13.234 23.608 ;
      RECT MASK 2 13.996 23.381 20.636 23.421 ;
      RECT MASK 2 2.136 23.388 3.159 23.412 ;
      RECT MASK 2 0.825 23.39 1.583 23.43 ;
      RECT MASK 2 22.865 23.43 23.317 23.45 ;
      RECT MASK 2 2.136 23.478 3.159 23.502 ;
      RECT MASK 2 14.781 23.548 15.96 23.588 ;
      RECT MASK 2 16.109 23.548 17.288 23.588 ;
      RECT MASK 2 17.437 23.548 18.616 23.588 ;
      RECT MASK 2 18.765 23.548 19.944 23.588 ;
      RECT MASK 2 0.825 23.55 1.583 23.59 ;
      RECT MASK 2 2.422 23.568 2.874 23.592 ;
      RECT MASK 2 23.232 23.59 23.653 23.61 ;
      RECT MASK 2 3.955 23.632 5.936 23.672 ;
      RECT MASK 2 14.072 23.6425 14.252 23.6825 ;
      RECT MASK 2 20.38 23.6425 20.56 23.6825 ;
      RECT MASK 2 2.625 23.658 2.874 23.682 ;
      RECT MASK 2 15.151 23.715 15.995 23.755 ;
      RECT MASK 2 16.479 23.715 17.323 23.755 ;
      RECT MASK 2 17.807 23.715 18.651 23.755 ;
      RECT MASK 2 19.135 23.715 19.979 23.755 ;
      RECT MASK 2 6.079 23.748 6.307 23.788 ;
      RECT MASK 2 9.912 23.748 10.472 23.788 ;
      RECT MASK 2 10.79 23.748 11.018 23.788 ;
      RECT MASK 2 11.738 23.748 11.966 23.788 ;
      RECT MASK 2 12.319 23.748 13.068 23.788 ;
      RECT MASK 2 22.46 23.75 24.26 23.77 ;
      RECT MASK 2 22.46 23.83 24.26 23.85 ;
      RECT MASK 2 1.074 23.925 1.334 23.965 ;
      RECT MASK 2 5.761 23.95 13.508 23.99 ;
      RECT MASK 2 4.104 24.008 4.164 24.238 ;
      RECT MASK 2 5.33 24.008 5.39 24.238 ;
      RECT MASK 2 0.832 24.085 1.576 24.125 ;
      RECT MASK 2 15.151 24.125 15.995 24.165 ;
      RECT MASK 2 16.479 24.125 17.323 24.165 ;
      RECT MASK 2 17.807 24.125 18.651 24.165 ;
      RECT MASK 2 19.135 24.125 19.979 24.165 ;
      RECT MASK 2 9.268 24.152 9.579 24.192 ;
      RECT MASK 2 10.126 24.152 10.804 24.192 ;
      RECT MASK 2 11.982 24.152 12.3 24.192 ;
      RECT MASK 2 12.485 24.152 12.927 24.192 ;
      RECT MASK 2 13.061 24.152 13.425 24.192 ;
      RECT MASK 2 14.072 24.1975 14.252 24.2375 ;
      RECT MASK 2 20.38 24.1975 20.56 24.2375 ;
      RECT MASK 2 14.781 24.292 15.96 24.332 ;
      RECT MASK 2 16.109 24.292 17.288 24.332 ;
      RECT MASK 2 17.437 24.292 18.616 24.332 ;
      RECT MASK 2 18.765 24.292 19.944 24.332 ;
      RECT MASK 2 2.212 24.303 3.159 24.327 ;
      RECT MASK 2 6.222 24.332 6.282 24.562 ;
      RECT MASK 2 6.554 24.332 6.614 24.562 ;
      RECT MASK 2 6.886 24.332 6.946 24.562 ;
      RECT MASK 2 7.218 24.332 7.278 24.562 ;
      RECT MASK 2 7.55 24.332 7.61 24.562 ;
      RECT MASK 2 7.882 24.332 7.942 24.562 ;
      RECT MASK 2 8.214 24.332 8.274 24.562 ;
      RECT MASK 2 8.546 24.332 8.606 24.562 ;
      RECT MASK 2 8.878 24.332 8.938 24.562 ;
      RECT MASK 2 9.21 24.332 9.27 24.562 ;
      RECT MASK 2 9.542 24.332 9.602 24.562 ;
      RECT MASK 2 10.269 24.332 10.329 24.562 ;
      RECT MASK 2 10.601 24.332 10.661 24.562 ;
      RECT MASK 2 11.265 24.332 11.325 24.562 ;
      RECT MASK 2 11.597 24.332 11.657 24.562 ;
      RECT MASK 2 11.929 24.332 11.989 24.562 ;
      RECT MASK 2 12.51 24.332 12.57 24.562 ;
      RECT MASK 2 12.842 24.332 12.902 24.562 ;
      RECT MASK 2 13.174 24.332 13.234 24.562 ;
      RECT MASK 2 0.832 24.36 1.576 24.4 ;
      RECT MASK 2 2.422 24.393 2.874 24.417 ;
      RECT MASK 2 13.996 24.459 20.636 24.499 ;
      RECT MASK 2 3.898 24.479 5.936 24.519 ;
      RECT MASK 2 2.422 24.483 2.874 24.507 ;
      RECT MASK 2 0.832 24.52 1.586 24.56 ;
      RECT MASK 2 2.212 24.573 3.159 24.597 ;
      RECT MASK 2 5.87 24.682 13.543 24.722 ;
      RECT MASK 2 3.948 24.71 4.566 24.75 ;
      RECT MASK 2 5.152 24.71 5.684 24.75 ;
      RECT MASK 2 13.996 24.821 20.636 24.861 ;
      RECT MASK 2 20.987 24.83 31.873 24.87 ;
      RECT MASK 2 0.825 24.86 1.583 24.9 ;
      RECT MASK 2 3.948 24.87 4.566 24.91 ;
      RECT MASK 2 5.152 24.87 5.684 24.91 ;
      RECT MASK 2 6.074 24.92 13.543 24.96 ;
      RECT MASK 2 14.781 24.988 15.96 25.028 ;
      RECT MASK 2 16.109 24.988 17.288 25.028 ;
      RECT MASK 2 17.437 24.988 18.616 25.028 ;
      RECT MASK 2 18.765 24.988 19.944 25.028 ;
      RECT MASK 2 20.987 24.99 31.873 25.03 ;
      RECT MASK 2 0.825 25.02 1.583 25.06 ;
      RECT MASK 2 6.074 25.08 13.543 25.12 ;
      RECT MASK 2 14.072 25.0825 14.252 25.1225 ;
      RECT MASK 2 20.38 25.0825 20.56 25.1225 ;
      RECT MASK 2 15.151 25.155 15.995 25.195 ;
      RECT MASK 2 16.479 25.155 17.323 25.195 ;
      RECT MASK 2 17.807 25.155 18.651 25.195 ;
      RECT MASK 2 19.135 25.155 19.979 25.195 ;
      RECT MASK 2 21.026 25.255 21.086 26.51 ;
      RECT MASK 2 25.526 25.255 25.586 26.561 ;
      RECT MASK 2 6.038 25.309 6.098 26.554 ;
      RECT MASK 2 13.238 25.309 13.298 26.513 ;
      RECT MASK 2 6.911 25.41 6.971 26.46 ;
      RECT MASK 2 7.185 25.41 7.245 26.46 ;
      RECT MASK 2 7.459 25.41 7.519 26.46 ;
      RECT MASK 2 7.733 25.41 7.793 26.46 ;
      RECT MASK 2 8.007 25.41 8.067 26.46 ;
      RECT MASK 2 8.281 25.41 8.341 26.46 ;
      RECT MASK 2 8.555 25.41 8.615 26.46 ;
      RECT MASK 2 8.829 25.41 8.889 26.46 ;
      RECT MASK 2 9.103 25.41 9.163 26.46 ;
      RECT MASK 2 9.377 25.41 9.437 26.46 ;
      RECT MASK 2 9.651 25.41 9.711 26.46 ;
      RECT MASK 2 9.925 25.41 9.985 26.46 ;
      RECT MASK 2 10.199 25.41 10.259 26.46 ;
      RECT MASK 2 10.473 25.41 10.533 26.46 ;
      RECT MASK 2 10.747 25.41 10.807 26.46 ;
      RECT MASK 2 11.021 25.41 11.081 26.46 ;
      RECT MASK 2 11.295 25.41 11.355 26.46 ;
      RECT MASK 2 11.569 25.41 11.629 26.46 ;
      RECT MASK 2 11.843 25.41 11.903 26.46 ;
      RECT MASK 2 12.117 25.41 12.177 26.46 ;
      RECT MASK 2 12.391 25.41 12.451 26.46 ;
      RECT MASK 2 21.986 25.41 22.046 26.46 ;
      RECT MASK 2 22.26 25.41 22.32 26.46 ;
      RECT MASK 2 22.534 25.41 22.594 26.46 ;
      RECT MASK 2 22.808 25.41 22.868 26.46 ;
      RECT MASK 2 23.082 25.41 23.142 26.46 ;
      RECT MASK 2 23.356 25.41 23.416 26.46 ;
      RECT MASK 2 23.63 25.41 23.69 26.46 ;
      RECT MASK 2 23.904 25.41 23.964 26.46 ;
      RECT MASK 2 24.178 25.41 24.238 26.46 ;
      RECT MASK 2 24.452 25.41 24.512 26.46 ;
      RECT MASK 2 24.726 25.41 24.786 26.46 ;
      RECT MASK 2 15.151 25.565 15.995 25.605 ;
      RECT MASK 2 16.479 25.565 17.323 25.605 ;
      RECT MASK 2 17.807 25.565 18.651 25.605 ;
      RECT MASK 2 19.135 25.565 19.979 25.605 ;
      RECT MASK 2 14.072 25.6375 14.252 25.6775 ;
      RECT MASK 2 20.38 25.6375 20.56 25.6775 ;
      RECT MASK 2 14.781 25.732 15.96 25.772 ;
      RECT MASK 2 16.109 25.732 17.288 25.772 ;
      RECT MASK 2 17.437 25.732 18.616 25.772 ;
      RECT MASK 2 18.765 25.732 19.944 25.772 ;
      RECT MASK 2 13.996 25.899 20.636 25.939 ;
      RECT MASK 2 14.107 26.24 20.525 26.28 ;
      RECT MASK 2 14.107 26.4 20.525 26.44 ;
      RECT MASK 2 5.994 26.69 13.43 26.83 ;
      RECT MASK 2 20.982 26.69 25.616 26.83 ;
  END
END dwc_ddrphy_por

END LIBRARY
