# LEF OUT API 
# Creation Date : Thu Dec 16 03:04:04 PST 2021
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_cmpana
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_cmpana 0 0 ;
  SYMMETRY X Y ;
  SIZE 100.8 BY 68.58 ;
  PIN Cmpdig_CalDac[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0955699375 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59003 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2723.8 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 4586.6 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 60.91875 100.8 61.01875 ;
    END
  END Cmpdig_CalDac[5]
  PIN Cmpdig_CalRef[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.08107 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.56393 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2647.8 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 4519.8 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 60.07875 100.8 60.17875 ;
    END
  END Cmpdig_CalRef[0]
  PIN Cmpdig_CalCmpr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7071299375 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.89082 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002808 LAYER D5 ;
      ANTENNAMAXAREACAR 1065.07 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 1828.95 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 59.41875 100.8 59.51875 ;
    END
  END Cmpdig_CalCmpr
  PIN Cmpdig_CalExt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.85112 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.15003 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2382.67 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 4137.56 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 58.93875 100.8 59.03875 ;
    END
  END Cmpdig_CalExt
  PIN InternalLoad
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 80.16 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 18.18 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.3 31.08 100.5 31.88 ;
    END
  END InternalLoad
  PIN ExternalLoad
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 272.462 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 49.5504 LAYER D8 ;
    ANTENNADIFFAREA 65.4797 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 3.841 63.20725 37.671 64.22725 ;
        RECT 3.841 60.64525 37.671 61.66525 ;
        RECT 3.841 58.08325 37.671 59.10325 ;
        RECT 3.841 55.52125 37.671 56.54125 ;
        RECT 4.309 50.48125 37.259 51.50125 ;
        RECT 4.309 47.91925 37.259 48.93925 ;
        RECT 4.309 45.35725 37.259 46.37725 ;
        RECT 4.309 42.79525 37.259 43.81525 ;
    END
  END ExternalLoad
  PIN Csr_CmprGainCurrAdj[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06692 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.53846 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002808 LAYER D5 ;
      ANTENNAMAXAREACAR 1334.25 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 2161.15 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 63.37875 100.8 63.47875 ;
    END
  END Csr_CmprGainCurrAdj[3]
  PIN PwrOk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.55512 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.81723 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 1826.94 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 2657.19 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 64.69875 100.8 64.79875 ;
    END
  END PwrOk
  PIN Csr_CmprGainCurrAdj[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77112 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.20602 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002808 LAYER D5 ;
      ANTENNAMAXAREACAR 879.197 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 1335.12 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 63.55875 100.8 63.65875 ;
    END
  END Csr_CmprGainCurrAdj[2]
  PIN Csr_CmprGainCurrAdj[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.62712 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.94683 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002808 LAYER D5 ;
      ANTENNAMAXAREACAR 845.008 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 1255.13 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 64.03875 100.8 64.13875 ;
    END
  END Csr_CmprGainCurrAdj[1]
  PIN Cmpdig_CalDac[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0952 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.58936 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2862.4 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 4686.08 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 62.71875 100.8 62.81875 ;
    END
  END Cmpdig_CalDac[0]
  PIN Cmpdig_CalDac[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0955699375 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59003 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2811.76 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 4649.94 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 62.05875 100.8 62.15875 ;
    END
  END Cmpdig_CalDac[2]
  PIN Cmpdig_CalDac[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.98712 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.59483 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 1905.55 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 3073.76 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 61.39875 100.8 61.49875 ;
    END
  END Cmpdig_CalDac[4]
  PIN Cmpdig_CalDac[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.41912 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.37242 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2187.96 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 3637.09 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 60.73875 100.8 60.83875 ;
    END
  END Cmpdig_CalDac[6]
  PIN Cmpdig_CalDac[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2755299375 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.11395 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2040.53 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 3411.27 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 60.25875 100.8 60.35875 ;
    END
  END Cmpdig_CalDac[7]
  PIN Csr_CmprGainCurrAdj[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0952 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.58936 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002808 LAYER D5 ;
      ANTENNAMAXAREACAR 1376.19 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 2202.22 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 64.21875 100.8 64.31875 ;
    END
  END Csr_CmprGainCurrAdj[0]
  PIN Cmpdig_CalRef[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0955699375 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59003 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2621.95 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 4513.27 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 59.59875 100.8 59.69875 ;
    END
  END Cmpdig_CalRef[1]
  PIN Cmpdig_CalInt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7791299375 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.02042 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2312.96 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 4027.09 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 58.75875 100.8 58.85875 ;
    END
  END Cmpdig_CalInt
  PIN Cmpdig_CalDac[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.20312 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.98362 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2086.11 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 3383.76 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 61.57875 100.8 61.67875 ;
    END
  END Cmpdig_CalDac[3]
  PIN Cmpdig_CalDac[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0955699375 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59003 LAYER D5 ;
    ANTENNADIFFAREA 0.324 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D5 ;
      ANTENNAMAXAREACAR 2825.65 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 4659.94 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 62.23875 100.8 62.33875 ;
    END
  END Cmpdig_CalDac[1]
  PIN Cmpana_Out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37682 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.51429 LAYER D5 ;
    ANTENNADIFFAREA 0.008424 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 58.355 100.8 58.455 ;
    END
  END Cmpana_Out
  PIN Csr_CmprGainCurrAdj[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087075 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.174735 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 65.17875 100.79975 65.27875 ;
    END
  END Csr_CmprGainCurrAdj[4]
  PIN Csr_CmprGainCurrAdj[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087075 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.174735 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 65.35875 100.79975 65.45875 ;
    END
  END Csr_CmprGainCurrAdj[5]
  PIN Csr_CmprGainCurrAdj[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087075 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.174735 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 65.83875 100.79975 65.93875 ;
    END
  END Csr_CmprGainCurrAdj[6]
  PIN Cmpdig_CmpanaClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2445 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2581 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D5 ;
      ANTENNAMAXAREACAR 1134.78 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 1361.48 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 57.96825 100.8 58.06825 ;
    END
  END Cmpdig_CmpanaClk
  PIN Csr_CmprGainCurrAdj[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087675 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.175815 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 66.01875 100.8 66.11875 ;
    END
  END Csr_CmprGainCurrAdj[7]
  PIN Csr_CmprBiasPowerUp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087675 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.175815 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 66.49875 100.8 66.59875 ;
    END
  END Csr_CmprBiasPowerUp
  PIN Csr_CmprBiasBypassEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087675 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.175815 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 66.67875 100.8 66.77875 ;
    END
  END Csr_CmprBiasBypassEn
  PIN Csr_CmprGainResAdj
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.087675 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.175815 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 67.15875 100.8 67.25875 ;
    END
  END Csr_CmprGainResAdj
  PIN Cmpdig_CmpanaEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.91512 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.46522 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003888 LAYER D5 ;
      ANTENNAMAXAREACAR 1278.74 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 1967.08 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 62.89875 100.8 62.99875 ;
    END
  END Cmpdig_CmpanaEn
  PIN PwrOk_VIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.625025 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.14304 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.6048 LAYER D5 ;
      ANTENNAMAXAREACAR 1.63579 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 2.5246 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 100.686 67.33875 100.8 67.43875 ;
    END
  END PwrOk_VIO
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER D8 ;
        RECT 0.3 32.48 100.5 33.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 66.08 100.5 66.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 1.68 100.5 2.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 4.48 100.5 5.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 7.28 100.5 8.08 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 10.08 100.5 10.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 26.88 100.5 27.68 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 29.68 100.5 30.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 12.88 100.5 13.68 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 15.68 100.5 16.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 18.48 100.5 19.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 21.28 100.5 22.08 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 24.08 100.5 24.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 63.28 100.5 64.08 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 60.48 100.5 61.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 57.68 100.5 58.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 36.68 100.5 37.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 40.88 100.5 41.68 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 45.08 100.5 45.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 49.28 100.5 50.08 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 53.48 100.5 54.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 3.841 64.64925 37.671 65.34925 ;
        RECT 3.841 62.08725 37.671 62.78725 ;
        RECT 3.841 59.52525 37.671 60.22525 ;
        RECT 3.841 56.96325 37.671 57.66325 ;
        RECT 3.841 54.40125 37.671 55.10125 ;
    END
  END VDDQ
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER D8 ;
        RECT 0.3 67.48 100.5 68.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 64.68 100.5 65.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 3.08 100.5 3.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 5.88 100.5 6.68 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 8.68 100.5 9.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 11.48 100.5 12.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 25.48 100.5 26.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 28.28 100.5 29.08 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 14.28 100.5 15.08 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 17.08 100.5 17.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 19.88 100.5 20.68 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 22.68 100.5 23.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 61.88 100.5 62.68 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 59.08 100.5 59.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 39.48 100.5 40.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 43.68 100.5 44.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 47.88 100.5 48.68 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 52.08 100.5 52.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 56.28 100.5 57.08 ;
    END
    PORT
      LAYER D8 ;
        RECT 4.309 51.92325 37.259 52.62325 ;
        RECT 4.309 49.36125 37.259 50.06125 ;
        RECT 4.309 46.79925 37.259 47.49925 ;
        RECT 4.309 44.23725 37.259 44.93725 ;
        RECT 4.309 41.67525 37.259 42.37525 ;
    END
    PORT
      LAYER D8 ;
        RECT 22.913 35.28 100.5 36.08 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER D8 ;
        RECT 0.3 33.88 100.5 34.68 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.3 38.08 100.5 38.88 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 42.28 100.5 43.08 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 46.48 100.5 47.28 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 50.68 100.5 51.48 ;
    END
    PORT
      LAYER D8 ;
        RECT 40.006 54.88 100.5 55.68 ;
    END
  END VDD
  OBS
    LAYER M1 SPACING 0 ;
      RECT 0 0 100.8 68.58 ;
    LAYER M2 SPACING 0 ;
      RECT 0 0 100.8 68.58 ;
    LAYER M3 SPACING 0 ;
      RECT 0 0 100.8 68.58 ;
    LAYER M4 SPACING 0 ;
      RECT 0 0 100.8 68.58 ;
    LAYER D5 SPACING 0 ;
      POLYGON 0 0 0 68.58 100.8 68.58 100.8 67.43875 100.686 67.43875 100.686 67.33875 100.8 67.33875 100.8 67.25875 100.686 67.25875 100.686 67.15875 100.8 67.15875 100.8 66.77875 100.686 66.77875 100.686 66.67875 100.8 66.67875 100.8 66.59875 100.686 66.59875 100.686 66.49875 100.8 66.49875 100.8 66.11875 100.686 66.11875 100.686 66.01875 100.8 66.01875 100.8 65.93875 100.686 65.93875 100.686 65.83875 100.79975 65.83875 100.79975 65.93875 100.8 65.93875 100.8 65.45875 100.686 65.45875 100.686 65.35875 100.79975 65.35875 100.79975 65.45875 100.8 65.45875 100.8 65.27875 100.686 65.27875 100.686 65.17875 100.79975 65.17875 100.79975 65.27875 100.8 65.27875 100.8 64.79875 100.686 64.79875 100.686 64.69875 100.8 64.69875 100.8 64.31875 100.686 64.31875 100.686 64.21875 100.8 64.21875 100.8 64.13875 100.686 64.13875 100.686 64.03875 100.8 64.03875 100.8 63.65875 100.686 63.65875 100.686 63.55875 100.8 63.55875 100.8 63.47875 100.686 63.47875 100.686 63.37875 100.8 63.37875 100.8 62.99875 100.686 62.99875 100.686 62.89875 100.8 62.89875 100.8 62.81875 100.686 62.81875 100.686 62.71875 100.8 62.71875 100.8 62.33875 100.686 62.33875 100.686 62.23875 100.8 62.23875 100.8 62.15875 100.686 62.15875 100.686 62.05875 100.8 62.05875 100.8 61.67875 100.686 61.67875 100.686 61.57875 100.8 61.57875 100.8 61.49875 100.686 61.49875 100.686 61.39875 100.8 61.39875 100.8 61.01875 100.686 61.01875 100.686 60.91875 100.8 60.91875 100.8 60.83875 100.686 60.83875 100.686 60.73875 100.8 60.73875 100.8 60.35875 100.686 60.35875 100.686 60.25875 100.8 60.25875 100.8 60.17875 100.686 60.17875 100.686 60.07875 100.8 60.07875 100.8 59.69875 100.686 59.69875 100.686 59.59875 100.8 59.59875 100.8 59.51875 100.686 59.51875 100.686 59.41875 100.8 59.41875 100.8 59.03875 100.686 59.03875 100.686 58.93875 100.8 58.93875 100.8 58.85875 100.686 58.85875 100.686 58.75875 100.8 58.75875 100.8 58.455 100.686 58.455 100.686 58.355 100.8 58.355 100.8 58.06825 100.686 58.06825 100.686 57.96825 100.8 57.96825 100.8 0 ;
    LAYER D6 SPACING 0 ;
      RECT 0 0 100.8 68.58 ;
    LAYER D7 SPACING 0 ;
      POLYGON 0 0 0 68.58 100.8 68.58 100.8 31.88 0.3 31.88 0.3 31.08 100.5 31.08 100.5 31.88 100.8 31.88 100.8 0 ;
  END
END dwc_ddrphy_cmpana

END LIBRARY
