# LEF OUT API 
# Creation Date : Tue Apr 16 16:06:36 IST 2019
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_pclk_master
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_pclk_master 0 0 ;
  SYMMETRY X Y ;
  SIZE 10.26 BY 48.96 ;
  PIN atpg_so
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05529 LAYER M4 ;
    ANTENNADIFFAREA 0.0074479375 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M4 ;
      ANTENNAMAXAREACAR 0 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 8.778 0.114 8.854 ;
    END
  END atpg_so
  PIN PclkEn_Dq0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.03705 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 441.875 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 34.846 0.114 34.922 ;
    END
  END PclkEn_Dq0
  PIN PclkEnDiv2_Dq0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.029298 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 318.368 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 34.542 0.114 34.618 ;
    END
  END PclkEnDiv2_Dq0
  PIN Pclk_Dq0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.728 LAYER M6 ;
    ANTENNADIFFAREA 0.806736 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 0 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0.3 29.02 9.96 29.42 ;
        RECT 0.3 26.32 9.96 26.72 ;
    END
  END Pclk_Dq0
  PIN PclkEn_Ca0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.03705 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 440.229 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 47.006 0.114 47.082 ;
    END
  END PclkEn_Ca0
  PIN PclkEnDiv2_Ca0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.029298 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 326.724 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 46.702 0.114 46.778 ;
    END
  END PclkEnDiv2_Ca0
  PIN Pclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.031464 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 2.13095 LAYER M5 ;
    ANTENNAPARTIALCUTAREA 0.001444 LAYER VIA4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER VIA4 ;
    ANTENNADIFFAREA 0 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M4 ;
      ANTENNAGATEAREA 0 LAYER VIA4 ;
      ANTENNAGATEAREA 0.041984 LAYER M5 ;
      ANTENNAMAXAREACAR 0 LAYER M4 ;
      ANTENNAMAXAREACAR 79.834599938 LAYER M5 ;
      ANTENNAMAXCUTCAR 0 LAYER VIA4 ;
    PORT
      LAYER M4 ;
        RECT 0 26.334 0.114 26.41 ;
    END
  END Pclk
  PIN Pclk_Ca0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.728 LAYER M6 ;
    ANTENNADIFFAREA 0.806736 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 0 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0.3 41.26 9.96 41.66 ;
        RECT 0.3 38.56 9.96 38.96 ;
    END
  END Pclk_Ca0
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.3 47.95 9.96 48.45 ;
        RECT 0.3 47.25 9.96 47.75 ;
        RECT 0.3 43.51 9.96 44.01 ;
        RECT 0.3 42.56 9.96 43.06 ;
        RECT 0.3 41.86 9.96 42.36 ;
        RECT 0.3 37.86 9.96 38.36 ;
        RECT 0.3 37.16 9.96 37.66 ;
        RECT 0.3 35.71 9.96 36.21 ;
        RECT 0.3 35.01 9.96 35.51 ;
        RECT 0.3 31.27 9.96 31.77 ;
        RECT 0.3 30.32 9.96 30.82 ;
        RECT 0.3 29.62 9.96 30.12 ;
        RECT 0.3 25.62 9.96 26.12 ;
        RECT 0.3 24.92 9.96 25.42 ;
        RECT 0.3 23.47 9.96 23.97 ;
        RECT 0.3 22.77 9.96 23.27 ;
        RECT 0.3 19.03 9.96 19.53 ;
        RECT 0.3 18.08 9.96 18.58 ;
        RECT 0.3 17.38 9.96 17.88 ;
        RECT 0.3 13.38 9.96 13.88 ;
        RECT 0.3 12.68 9.96 13.18 ;
        RECT 0.3 11.23 9.96 11.73 ;
        RECT 0.3 10.53 9.96 11.03 ;
        RECT 0.3 6.79 9.96 7.29 ;
        RECT 0.3 5.84 9.96 6.34 ;
        RECT 0.3 5.14 9.96 5.64 ;
        RECT 0.3 1.14 9.96 1.64 ;
        RECT 0.3 0.44 9.96 0.94 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M6 ;
        RECT 0.3 46.55 9.96 47.05 ;
        RECT 0.3 45.85 9.96 46.35 ;
        RECT 0.3 44.91 9.96 45.41 ;
        RECT 0.3 44.21 9.96 44.71 ;
        RECT 0.3 40.56 9.96 41.06 ;
        RECT 0.3 39.86 9.96 40.36 ;
        RECT 0.3 39.16 9.96 39.66 ;
        RECT 0.3 34.31 9.96 34.81 ;
        RECT 0.3 33.61 9.96 34.11 ;
        RECT 0.3 32.67 9.96 33.17 ;
        RECT 0.3 31.97 9.96 32.47 ;
        RECT 0.3 28.32 9.96 28.82 ;
        RECT 0.3 27.62 9.96 28.12 ;
        RECT 0.3 26.92 9.96 27.42 ;
        RECT 0.3 22.07 9.96 22.57 ;
        RECT 0.3 21.37 9.96 21.87 ;
        RECT 0.3 20.43 9.96 20.93 ;
        RECT 0.3 19.73 9.96 20.23 ;
        RECT 0.3 16.08 9.96 16.58 ;
        RECT 0.3 15.38 9.96 15.88 ;
        RECT 0.3 14.68 9.96 15.18 ;
        RECT 0.3 9.83 9.96 10.33 ;
        RECT 0.3 9.13 9.96 9.63 ;
        RECT 0.3 8.19 9.96 8.69 ;
        RECT 0.3 7.49 9.96 7.99 ;
        RECT 0.3 3.84 9.96 4.34 ;
        RECT 0.3 3.14 9.96 3.64 ;
        RECT 0.3 2.44 9.96 2.94 ;
    END
  END VSS
  PIN atpg_si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.045448 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 297.195 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 47.31 0.114 47.386 ;
    END
  END atpg_si
  PIN Reset_async
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.039482 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002432 LAYER M4 ;
      ANTENNAMAXAREACAR 47.6174 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 26.03 0.114 26.106 ;
    END
  END Reset_async
  PIN PclkEn_Ca1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.035644 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 432.737 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 22.61 0.114 22.686 ;
    END
  END PclkEn_Ca1
  PIN PclkEnDiv2_Ca1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.029298 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 316.296 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 22.306 0.114 22.382 ;
    END
  END PclkEnDiv2_Ca1
  PIN Pclk_Ca1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.728 LAYER M6 ;
    ANTENNADIFFAREA 0.806736 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 0 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0.3 16.78 9.96 17.18 ;
        RECT 0.3 14.08 9.96 14.48 ;
    END
  END Pclk_Ca1
  PIN PclkEn_Dq1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.035644 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 434.546 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 10.374 0.114 10.45 ;
    END
  END PclkEn_Dq1
  PIN PclkEnDiv2_Dq1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.029298 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.000608 LAYER M4 ;
      ANTENNAMAXAREACAR 314.817 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 10.07 0.114 10.146 ;
    END
  END PclkEnDiv2_Dq1
  PIN atpg_se
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.023864 LAYER M4 ;
    ANTENNADIFFAREA 0 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002432 LAYER M4 ;
      ANTENNAMAXAREACAR 55.3059 LAYER M4 ;
    PORT
      LAYER M4 ;
        RECT 0 26.638 0.114 26.714 ;
    END
  END atpg_se
  PIN Pclk_Dq1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.728 LAYER M6 ;
    ANTENNADIFFAREA 0.806736 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0 LAYER M6 ;
      ANTENNAMAXAREACAR 0 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0.3 1.84 9.96 2.24 ;
    END
    PORT
      LAYER M6 ;
        RECT 0.3 4.54 9.96 4.94 ;
    END
  END Pclk_Dq1
  OBS
    LAYER M1 ;
      RECT MASK 1 0 0 10.26 48.96 ;
    LAYER M1 ;
      RECT MASK 2 0 0 10.26 48.96 ;
    LAYER M2 ;
      RECT MASK 1 0 0 10.26 48.96 ;
    LAYER M2 ;
      RECT MASK 2 0 0 10.26 48.96 ;
    LAYER M3 ;
      RECT MASK 1 0 0 10.26 48.96 ;
    LAYER M4 ;
      POLYGON 10.26 0 10.26 48.96 0 48.96 0 47.462 0.19 47.462 0.19 47.234 0 47.234 0 47.158 0.19 47.158 0.19 46.93 0 46.93 0 46.854 0.19 46.854 0.19 46.626 0 46.626 0 34.998 0.19 34.998 0.19 34.77 0 34.77 0 34.694 0.19 34.694 0.19 34.466 0 34.466 0 26.79 0.19 26.79 0.19 26.562 0 26.562 0 26.486 0.19 26.486 0.19 26.258 0 26.258 0 26.182 0.19 26.182 0.19 25.954 0 25.954 0 22.762 0.19 22.762 0.19 22.534 0 22.534 0 22.458 0.19 22.458 0.19 22.23 0 22.23 0 10.526 0.19 10.526 0.19 10.298 0 10.298 0 10.222 0.19 10.222 0.19 9.994 0 9.994 0 8.93 0.19 8.93 0.19 8.702 0 8.702 0 0 ;
    LAYER M3 ;
      RECT MASK 2 0 0 10.26 48.96 ;
    LAYER M4 ;
      RECT 1.859 6.605 8.774 6.665 ;
      RECT 1.859 6.725 8.774 6.785 ;
      RECT 1.859 6.845 8.7745 6.905 ;
      RECT 1.859 6.965 8.774 7.025 ;
      RECT 1.859 7.085 8.774 7.145 ;
      RECT 1.859 7.325 8.774 7.385 ;
      RECT 1.859 7.445 8.7745 7.505 ;
      RECT 1.859 7.565 8.774 7.625 ;
      RECT 1.859 7.685 8.774 7.745 ;
      RECT 1.951 8.105 8.774 8.165 ;
      RECT 1.951 8.225 8.774 8.285 ;
      RECT 1.951 8.345 8.7745 8.405 ;
      RECT 1.951 8.465 8.774 8.525 ;
      RECT 0.19 8.778 0.7275 8.854 ;
      RECT 1.951 8.825 8.774 8.885 ;
      RECT 1.951 8.945 8.7745 9.005 ;
      RECT 1.951 9.065 8.774 9.125 ;
      RECT 1.951 9.185 8.774 9.245 ;
      RECT 2.5215 9.305 9.09 9.365 ;
      RECT 3.184 9.425 9.09 9.485 ;
      RECT 0.172 9.486 0.447 9.546 ;
      RECT 3.5765 9.791 6.243 9.871 ;
      RECT 3.5905 10.031 6.243 10.111 ;
      RECT 0.19 10.07 0.3855 10.146 ;
      RECT 3.233 10.171 6.5675 10.211 ;
      RECT 3.5765 10.271 6.243 10.351 ;
      RECT 0.19 10.374 0.469 10.45 ;
      RECT 3.3275 10.411 6.4705 10.451 ;
      RECT 3.5905 10.511 6.243 10.591 ;
      RECT 1.906 10.651 4.978 10.691 ;
      RECT 0.179 10.6675 0.5795 10.7435 ;
      RECT 3.5765 10.751 6.243 10.831 ;
      RECT 0.728 12.885 2.984 12.945 ;
      RECT 1.859 18.845 8.774 18.905 ;
      RECT 1.859 18.965 8.774 19.025 ;
      RECT 1.859 19.085 8.7745 19.145 ;
      RECT 1.859 19.205 8.774 19.265 ;
      RECT 1.859 19.325 8.774 19.385 ;
      RECT 1.859 19.565 8.774 19.625 ;
      RECT 1.859 19.685 8.7745 19.745 ;
      RECT 1.859 19.805 8.774 19.865 ;
      RECT 1.859 19.925 8.774 19.985 ;
      RECT 1.951 20.345 8.774 20.405 ;
      RECT 1.951 20.465 8.774 20.525 ;
      RECT 1.951 20.585 8.7745 20.645 ;
      RECT 1.951 20.705 8.774 20.765 ;
      RECT 1.951 21.065 8.774 21.125 ;
      RECT 1.951 21.185 8.7745 21.245 ;
      RECT 1.951 21.305 8.774 21.365 ;
      RECT 1.951 21.425 8.774 21.485 ;
      RECT 0.172 21.5415 0.447 21.6015 ;
      RECT 2.5215 21.545 9.09 21.605 ;
      RECT 0.2965 21.6615 0.6075 21.7215 ;
      RECT 3.184 21.665 9.09 21.725 ;
      RECT 3.5765 22.031 6.243 22.111 ;
      RECT 3.5905 22.271 6.243 22.351 ;
      RECT 0.19 22.306 0.3855 22.382 ;
      RECT 3.233 22.411 6.5675 22.451 ;
      RECT 3.5765 22.511 6.243 22.591 ;
      RECT 0.19 22.61 0.469 22.686 ;
      RECT 3.3275 22.651 6.4705 22.691 ;
      RECT 3.5905 22.751 6.243 22.831 ;
      RECT 1.906 22.891 4.978 22.931 ;
      RECT 0.2435 22.9065 0.5795 22.9825 ;
      RECT 3.5765 22.991 6.243 23.071 ;
      RECT 0.6135 25.725 2.8065 25.785 ;
      RECT 0.19 26.03 0.5195 26.106 ;
      RECT 0.6135 26.205 2.8065 26.265 ;
      RECT 0.19 26.334 0.414 26.41 ;
      RECT 0.19 26.638 0.314 26.714 ;
      RECT 0.6135 26.685 2.8065 26.745 ;
      RECT 1.859 31.085 8.774 31.145 ;
      RECT 1.859 31.205 8.774 31.265 ;
      RECT 1.859 31.325 8.7745 31.385 ;
      RECT 1.859 31.445 8.774 31.505 ;
      RECT 1.859 31.565 8.774 31.625 ;
      RECT 1.859 31.805 8.774 31.865 ;
      RECT 1.859 31.925 8.7745 31.985 ;
      RECT 1.859 32.045 8.774 32.105 ;
      RECT 1.859 32.165 8.774 32.225 ;
      RECT 1.951 32.585 8.774 32.645 ;
      RECT 1.951 32.705 8.774 32.765 ;
      RECT 1.951 32.825 8.7745 32.885 ;
      RECT 1.951 32.945 8.774 33.005 ;
      RECT 1.951 33.305 8.774 33.365 ;
      RECT 1.951 33.425 8.7745 33.485 ;
      RECT 1.951 33.545 8.774 33.605 ;
      RECT 1.951 33.665 8.774 33.725 ;
      RECT 0.172 33.7815 0.447 33.8415 ;
      RECT 2.5215 33.785 9.09 33.845 ;
      RECT 0.2965 33.9015 0.6075 33.9615 ;
      RECT 3.184 33.905 9.09 33.965 ;
      RECT 3.5765 34.271 6.243 34.351 ;
      RECT 3.5905 34.511 6.243 34.591 ;
      RECT 0.19 34.542 0.3855 34.618 ;
      RECT 3.213 34.651 6.5675 34.691 ;
      RECT 3.5765 34.751 6.243 34.831 ;
      RECT 0.19 34.846 0.4875 34.922 ;
      RECT 3.3275 34.891 6.4705 34.931 ;
      RECT 3.5905 34.991 6.243 35.071 ;
      RECT 1.906 35.131 4.978 35.171 ;
      RECT 3.5765 35.231 6.243 35.311 ;
      RECT 0.255 35.506 0.6045 35.582 ;
      RECT 1.859 43.325 8.774 43.385 ;
      RECT 1.859 43.445 8.774 43.505 ;
      RECT 1.859 43.565 8.7745 43.625 ;
      RECT 1.859 43.685 8.774 43.745 ;
      RECT 1.859 43.805 8.774 43.865 ;
      RECT 1.859 44.045 8.774 44.105 ;
      RECT 1.859 44.165 8.7745 44.225 ;
      RECT 1.859 44.285 8.774 44.345 ;
      RECT 1.859 44.405 8.774 44.465 ;
      RECT 1.951 44.825 8.774 44.885 ;
      RECT 1.951 44.945 8.774 45.005 ;
      RECT 1.951 45.065 8.7745 45.125 ;
      RECT 1.951 45.185 8.774 45.245 ;
      RECT 1.951 45.545 8.774 45.605 ;
      RECT 1.951 45.665 8.7745 45.725 ;
      RECT 1.951 45.785 8.774 45.845 ;
      RECT 1.951 45.905 8.774 45.965 ;
      RECT 0.172 46.0215 0.447 46.0815 ;
      RECT 2.5215 46.025 9.09 46.085 ;
      RECT 0.2965 46.1415 0.6075 46.2015 ;
      RECT 3.184 46.145 9.09 46.205 ;
      RECT 3.5765 46.511 6.243 46.591 ;
      RECT 0.19 46.702 0.3855 46.778 ;
      RECT 3.5905 46.751 6.243 46.831 ;
      RECT 3.2135 46.891 6.5675 46.931 ;
      RECT 3.5765 46.991 6.243 47.071 ;
      RECT 0.19 47.006 0.4875 47.082 ;
      RECT 3.3275 47.131 6.4705 47.171 ;
      RECT 3.5905 47.231 6.243 47.311 ;
      RECT 0.19 47.31 0.598 47.386 ;
      RECT 1.906 47.371 4.978 47.411 ;
      RECT 3.5765 47.471 6.243 47.551 ;
    LAYER M5 ;
      RECT 0 0 10.26 48.96 ;
    LAYER M4 ;
      RECT 0.704 12.645 3.009 12.705 ;
      RECT 0.7265 13.125 2.984 13.185 ;
      RECT 0.635 25.965 2.8005 26.025 ;
      RECT 1.9565 26.325 3.3785 26.385 ;
      RECT 0.635 26.445 2.8005 26.505 ;
      RECT 2.1675 26.955 3.498 27.015 ;
    LAYER M5 ;
      RECT 6.4665 0.897 6.5245 5.01 ;
      RECT 5.5545 0.985 5.6125 5.01 ;
      RECT 4.8705 1.018 4.9285 5.01 ;
      RECT 3.6165 5.1485 3.6745 5.6315 ;
      RECT 3.8445 5.1485 3.9025 5.6315 ;
      RECT 4.0725 5.1485 4.1305 5.6315 ;
      RECT 4.3005 5.1485 4.3585 5.6315 ;
      RECT 4.5285 5.1485 4.5865 5.6315 ;
      RECT 4.7565 5.1485 4.8145 5.6315 ;
      RECT 4.9845 5.1485 5.0425 5.6315 ;
      RECT 5.2125 5.1485 5.2705 5.6315 ;
      RECT 5.4405 5.1485 5.4985 5.6315 ;
      RECT 5.6685 5.1485 5.7265 5.6315 ;
      RECT 5.8965 5.1485 5.9545 5.6315 ;
      RECT 6.1245 5.1485 6.1825 5.6315 ;
      RECT 6.3525 5.1485 6.4105 5.6315 ;
      RECT 6.5805 5.1485 6.6385 5.6315 ;
      RECT 6.8085 5.1485 6.8665 5.6315 ;
      RECT 7.0365 5.1485 7.0945 5.6315 ;
      RECT 7.2645 5.1485 7.3225 5.6315 ;
      RECT 7.4925 5.1485 7.5505 5.6315 ;
      RECT 7.7205 5.1485 7.7785 5.6315 ;
      RECT 1.9065 5.8485 1.9645 7.784 ;
      RECT 2.0205 5.8485 2.0785 7.311 ;
      RECT 2.1345 5.8485 2.1925 7.784 ;
      RECT 2.3625 5.8485 2.4205 7.6685 ;
      RECT 2.5905 5.8485 2.6485 7.6685 ;
      RECT 2.8185 5.8485 2.8765 7.784 ;
      RECT 3.0465 5.8485 3.1045 7.784 ;
      RECT 3.5025 5.8485 3.5605 7.784 ;
      RECT 3.9585 6.203 4.0165 7.784 ;
      RECT 4.1865 6.203 4.2445 7.784 ;
      RECT 4.4145 6.203 4.4725 7.784 ;
      RECT 4.6425 6.203 4.7005 7.784 ;
      RECT 5.0985 6.203 5.1565 7.784 ;
      RECT 5.3265 6.203 5.3845 7.784 ;
      RECT 5.7825 6.203 5.8405 7.784 ;
      RECT 6.0105 6.203 6.0685 7.784 ;
      RECT 6.2385 6.203 6.2965 7.784 ;
      RECT 3.7305 6.238 3.7885 7.784 ;
      RECT 4.8705 6.238 4.9285 7.784 ;
      RECT 5.5545 6.238 5.6125 7.784 ;
      RECT 6.4665 6.238 6.5245 7.784 ;
      RECT 3.6165 6.326 3.6745 6.584 ;
      RECT 3.8445 6.326 3.9025 7.311 ;
      RECT 4.0725 6.326 4.1305 6.584 ;
      RECT 4.3005 6.326 4.3585 6.584 ;
      RECT 4.5285 6.326 4.5865 6.584 ;
      RECT 4.7565 6.326 4.8145 6.584 ;
      RECT 4.9845 6.326 5.0425 6.584 ;
      RECT 5.2125 6.326 5.2705 6.584 ;
      RECT 5.4405 6.326 5.4985 6.584 ;
      RECT 5.6685 6.326 5.7265 6.584 ;
      RECT 5.8965 6.326 5.9545 6.584 ;
      RECT 6.1245 6.326 6.1825 6.584 ;
      RECT 6.3525 6.326 6.4105 6.584 ;
      RECT 6.5805 6.326 6.6385 6.584 ;
      RECT 6.8085 6.326 6.8665 6.584 ;
      RECT 7.0365 6.326 7.0945 6.584 ;
      RECT 7.2645 6.326 7.3225 6.584 ;
      RECT 7.4925 6.326 7.5505 6.584 ;
      RECT 7.7205 6.326 7.7785 6.584 ;
      RECT 8.8605 7.4885 8.9185 10.3345 ;
      RECT 9.0885 7.4885 9.1465 10.3345 ;
      RECT 9.3165 7.4885 9.3745 10.3345 ;
      RECT 2.0205 7.4925 2.0785 9.284 ;
      RECT 2.2485 7.4925 2.3065 9.284 ;
      RECT 2.4765 7.4925 2.5345 9.284 ;
      RECT 2.7045 7.4925 2.7625 9.284 ;
      RECT 2.9325 7.4925 2.9905 9.284 ;
      RECT 3.6165 7.4925 3.6745 10.9475 ;
      RECT 3.8445 7.4925 3.9025 10.95 ;
      RECT 4.0725 7.4925 4.1305 10.95 ;
      RECT 4.3005 7.4925 4.3585 10.95 ;
      RECT 4.5285 7.4925 4.5865 10.95 ;
      RECT 4.7565 7.4925 4.8145 10.95 ;
      RECT 4.9845 7.4925 5.0425 10.95 ;
      RECT 5.2125 7.4925 5.2705 10.95 ;
      RECT 5.4405 7.4925 5.4985 10.95 ;
      RECT 5.6685 7.4925 5.7265 10.95 ;
      RECT 5.8965 7.4925 5.9545 10.95 ;
      RECT 6.1245 7.4925 6.1825 10.95 ;
      RECT 6.3525 7.4925 6.4105 9.284 ;
      RECT 6.5805 7.4925 6.6385 9.284 ;
      RECT 2.3625 7.856 2.4205 9.936 ;
      RECT 2.5905 7.856 2.6485 9.936 ;
      RECT 3.0465 8.0605 3.1045 9.284 ;
      RECT 3.5025 8.0605 3.5605 9.284 ;
      RECT 6.8085 8.864 6.8665 10.3355 ;
      RECT 7.0365 8.864 7.0945 10.3355 ;
      RECT 7.2645 8.864 7.3225 10.3355 ;
      RECT 7.4925 8.864 7.5505 10.3355 ;
      RECT 7.7205 8.864 7.7785 10.3355 ;
      RECT 7.9485 8.864 8.0065 10.3345 ;
      RECT 8.1765 8.864 8.2345 10.3345 ;
      RECT 8.4045 8.864 8.4625 10.3345 ;
      RECT 8.6325 8.864 8.6905 10.3345 ;
      RECT 0.3105 9.417 0.3685 46.1575 ;
      RECT 3.2745 10.119 3.3325 46.984 ;
      RECT 3.3885 10.346 3.4465 47.2295 ;
      RECT 6.9225 10.441 6.9805 11.75 ;
      RECT 0.4245 10.627 0.4825 21.805 ;
      RECT 0.7665 12.5735 0.8245 13.226 ;
      RECT 0.8805 12.5735 0.9385 15.176 ;
      RECT 0.9945 12.5735 1.0525 13.226 ;
      RECT 1.1085 12.5735 1.1665 15.176 ;
      RECT 1.2225 12.5735 1.2805 13.226 ;
      RECT 1.3365 12.5735 1.3945 15.176 ;
      RECT 1.4505 12.5735 1.5085 13.226 ;
      RECT 1.5645 12.5735 1.6225 15.176 ;
      RECT 1.6785 12.5735 1.7365 13.226 ;
      RECT 1.7925 12.5735 1.8505 15.179 ;
      RECT 1.9065 12.5735 1.9645 13.226 ;
      RECT 2.0205 12.5735 2.0785 15.179 ;
      RECT 2.1345 12.5735 2.1925 13.226 ;
      RECT 2.2485 12.5735 2.3065 15.179 ;
      RECT 2.3625 12.5735 2.4205 13.226 ;
      RECT 2.4765 12.5735 2.5345 15.179 ;
      RECT 2.5905 12.5735 2.6485 13.226 ;
      RECT 2.7045 12.5735 2.7625 15.179 ;
      RECT 2.8185 12.5735 2.8765 13.226 ;
      RECT 6.4665 13.137 6.5245 17.25 ;
      RECT 5.5545 13.225 5.6125 17.25 ;
      RECT 4.8705 13.258 4.9285 17.25 ;
      RECT 3.6165 17.3885 3.6745 17.8715 ;
      RECT 3.8445 17.3885 3.9025 17.8715 ;
      RECT 4.0725 17.3885 4.1305 17.8715 ;
      RECT 4.3005 17.3885 4.3585 17.8715 ;
      RECT 4.5285 17.3885 4.5865 17.8715 ;
      RECT 4.7565 17.3885 4.8145 17.8715 ;
      RECT 4.9845 17.3885 5.0425 17.8715 ;
      RECT 5.2125 17.3885 5.2705 17.8715 ;
      RECT 5.4405 17.3885 5.4985 17.8715 ;
      RECT 5.6685 17.3885 5.7265 17.8715 ;
      RECT 5.8965 17.3885 5.9545 17.8715 ;
      RECT 6.1245 17.3885 6.1825 17.8715 ;
      RECT 6.3525 17.3885 6.4105 17.8715 ;
      RECT 6.5805 17.3885 6.6385 17.8715 ;
      RECT 6.8085 17.3885 6.8665 17.8715 ;
      RECT 7.0365 17.3885 7.0945 17.8715 ;
      RECT 7.2645 17.3885 7.3225 17.8715 ;
      RECT 7.4925 17.3885 7.5505 17.8715 ;
      RECT 7.7205 17.3885 7.7785 17.8715 ;
      RECT 1.9065 18.0885 1.9645 20.024 ;
      RECT 2.0205 18.0885 2.0785 19.551 ;
      RECT 2.1345 18.0885 2.1925 20.024 ;
      RECT 2.3625 18.0885 2.4205 19.9085 ;
      RECT 2.5905 18.0885 2.6485 19.9085 ;
      RECT 2.8185 18.0885 2.8765 20.024 ;
      RECT 3.0465 18.0885 3.1045 20.024 ;
      RECT 3.5025 18.0885 3.5605 20.024 ;
      RECT 3.9585 18.443 4.0165 20.024 ;
      RECT 4.1865 18.443 4.2445 20.024 ;
      RECT 4.4145 18.443 4.4725 20.024 ;
      RECT 4.6425 18.443 4.7005 20.024 ;
      RECT 5.0985 18.443 5.1565 20.024 ;
      RECT 5.3265 18.443 5.3845 20.024 ;
      RECT 5.7825 18.443 5.8405 20.024 ;
      RECT 6.0105 18.443 6.0685 20.024 ;
      RECT 6.2385 18.443 6.2965 20.024 ;
      RECT 3.7305 18.478 3.7885 20.024 ;
      RECT 4.8705 18.478 4.9285 20.024 ;
      RECT 5.5545 18.478 5.6125 20.024 ;
      RECT 6.4665 18.478 6.5245 20.024 ;
      RECT 3.6165 18.566 3.6745 18.824 ;
      RECT 3.8445 18.566 3.9025 19.551 ;
      RECT 4.0725 18.566 4.1305 18.824 ;
      RECT 4.3005 18.566 4.3585 18.824 ;
      RECT 4.5285 18.566 4.5865 18.824 ;
      RECT 4.7565 18.566 4.8145 18.824 ;
      RECT 4.9845 18.566 5.0425 18.824 ;
      RECT 5.2125 18.566 5.2705 18.824 ;
      RECT 5.4405 18.566 5.4985 18.824 ;
      RECT 5.6685 18.566 5.7265 18.824 ;
      RECT 5.8965 18.566 5.9545 18.824 ;
      RECT 6.1245 18.566 6.1825 18.824 ;
      RECT 6.3525 18.566 6.4105 18.824 ;
      RECT 6.5805 18.566 6.6385 18.824 ;
      RECT 6.8085 18.566 6.8665 18.824 ;
      RECT 7.0365 18.566 7.0945 18.824 ;
      RECT 7.2645 18.566 7.3225 18.824 ;
      RECT 7.4925 18.566 7.5505 18.824 ;
      RECT 7.7205 18.566 7.7785 18.824 ;
      RECT 8.8605 19.7285 8.9185 22.5745 ;
      RECT 9.0885 19.7285 9.1465 22.5745 ;
      RECT 9.3165 19.7285 9.3745 22.5745 ;
      RECT 2.0205 19.7325 2.0785 21.524 ;
      RECT 2.2485 19.7325 2.3065 21.524 ;
      RECT 2.4765 19.7325 2.5345 21.524 ;
      RECT 2.7045 19.7325 2.7625 21.524 ;
      RECT 2.9325 19.7325 2.9905 21.524 ;
      RECT 3.6165 19.7325 3.6745 23.1875 ;
      RECT 3.8445 19.7325 3.9025 23.19 ;
      RECT 4.0725 19.7325 4.1305 23.19 ;
      RECT 4.3005 19.7325 4.3585 23.19 ;
      RECT 4.5285 19.7325 4.5865 23.19 ;
      RECT 4.7565 19.7325 4.8145 23.19 ;
      RECT 4.9845 19.7325 5.0425 23.19 ;
      RECT 5.2125 19.7325 5.2705 23.19 ;
      RECT 5.4405 19.7325 5.4985 23.19 ;
      RECT 5.6685 19.7325 5.7265 23.19 ;
      RECT 5.8965 19.7325 5.9545 23.19 ;
      RECT 6.1245 19.7325 6.1825 23.19 ;
      RECT 6.3525 19.7325 6.4105 21.524 ;
      RECT 6.5805 19.7325 6.6385 21.524 ;
      RECT 2.3625 20.096 2.4205 22.176 ;
      RECT 2.5905 20.096 2.6485 22.176 ;
      RECT 3.0465 20.3005 3.1045 21.524 ;
      RECT 3.5025 20.3005 3.5605 21.524 ;
      RECT 6.8085 21.104 6.8665 22.5755 ;
      RECT 7.0365 21.104 7.0945 22.5755 ;
      RECT 7.2645 21.104 7.3225 22.5755 ;
      RECT 7.4925 21.104 7.5505 22.5755 ;
      RECT 7.7205 21.104 7.7785 22.5755 ;
      RECT 7.9485 21.104 8.0065 22.5745 ;
      RECT 8.1765 21.104 8.2345 22.5745 ;
      RECT 8.4045 21.104 8.4625 22.5745 ;
      RECT 8.6325 21.104 8.6905 22.5745 ;
      RECT 6.9225 22.681 6.9805 23.99 ;
      RECT 0.4245 22.8345 0.4825 34.0585 ;
      RECT 0.768 24.9165 0.826 26.571 ;
      RECT 0.996 24.9165 1.054 26.571 ;
      RECT 1.224 24.9165 1.282 26.571 ;
      RECT 1.452 24.9165 1.51 26.571 ;
      RECT 1.68 24.9165 1.738 26.571 ;
      RECT 1.908 24.92 1.966 26.568 ;
      RECT 2.136 24.92 2.194 26.568 ;
      RECT 2.364 24.92 2.422 26.568 ;
      RECT 2.592 24.92 2.65 26.568 ;
      RECT 6.4665 25.377 6.5245 29.49 ;
      RECT 5.5545 25.465 5.6125 29.49 ;
      RECT 4.8705 25.498 4.9285 29.49 ;
      RECT 0.654 25.65 0.712 28.82 ;
      RECT 0.882 25.65 0.94 28.82 ;
      RECT 1.11 25.65 1.168 28.82 ;
      RECT 1.338 25.65 1.396 28.82 ;
      RECT 1.566 25.65 1.624 28.82 ;
      RECT 1.794 25.65 1.852 28.82 ;
      RECT 2.022 25.65 2.08 28.82 ;
      RECT 2.25 25.65 2.308 28.82 ;
      RECT 2.478 25.65 2.536 28.82 ;
      RECT 2.706 25.65 2.764 28.82 ;
      RECT 3.6165 29.6285 3.6745 30.1115 ;
      RECT 3.8445 29.6285 3.9025 30.1115 ;
      RECT 4.0725 29.6285 4.1305 30.1115 ;
      RECT 4.3005 29.6285 4.3585 30.1115 ;
      RECT 4.5285 29.6285 4.5865 30.1115 ;
      RECT 4.7565 29.6285 4.8145 30.1115 ;
      RECT 4.9845 29.6285 5.0425 30.1115 ;
      RECT 5.2125 29.6285 5.2705 30.1115 ;
      RECT 5.4405 29.6285 5.4985 30.1115 ;
      RECT 5.6685 29.6285 5.7265 30.1115 ;
      RECT 5.8965 29.6285 5.9545 30.1115 ;
      RECT 6.1245 29.6285 6.1825 30.1115 ;
      RECT 6.3525 29.6285 6.4105 30.1115 ;
      RECT 6.5805 29.6285 6.6385 30.1115 ;
      RECT 6.8085 29.6285 6.8665 30.1115 ;
      RECT 7.0365 29.6285 7.0945 30.1115 ;
      RECT 7.2645 29.6285 7.3225 30.1115 ;
      RECT 7.4925 29.6285 7.5505 30.1115 ;
      RECT 7.7205 29.6285 7.7785 30.1115 ;
      RECT 1.9065 30.3285 1.9645 32.264 ;
      RECT 2.0205 30.3285 2.0785 31.791 ;
      RECT 2.1345 30.3285 2.1925 32.264 ;
      RECT 2.3625 30.3285 2.4205 32.1485 ;
      RECT 2.5905 30.3285 2.6485 32.1485 ;
      RECT 2.8185 30.3285 2.8765 32.264 ;
      RECT 3.0465 30.3285 3.1045 32.264 ;
      RECT 3.5025 30.3285 3.5605 32.264 ;
      RECT 3.9585 30.683 4.0165 32.264 ;
      RECT 4.1865 30.683 4.2445 32.264 ;
      RECT 4.4145 30.683 4.4725 32.264 ;
      RECT 4.6425 30.683 4.7005 32.264 ;
      RECT 5.0985 30.683 5.1565 32.264 ;
      RECT 5.3265 30.683 5.3845 32.264 ;
      RECT 5.7825 30.683 5.8405 32.264 ;
      RECT 6.0105 30.683 6.0685 32.264 ;
      RECT 6.2385 30.683 6.2965 32.264 ;
      RECT 3.7305 30.718 3.7885 32.264 ;
      RECT 4.8705 30.718 4.9285 32.264 ;
      RECT 5.5545 30.718 5.6125 32.264 ;
      RECT 6.4665 30.718 6.5245 32.264 ;
      RECT 3.6165 30.806 3.6745 31.064 ;
      RECT 3.8445 30.806 3.9025 31.791 ;
      RECT 4.0725 30.806 4.1305 31.064 ;
      RECT 4.3005 30.806 4.3585 31.064 ;
      RECT 4.5285 30.806 4.5865 31.064 ;
      RECT 4.7565 30.806 4.8145 31.064 ;
      RECT 4.9845 30.806 5.0425 31.064 ;
      RECT 5.2125 30.806 5.2705 31.064 ;
      RECT 5.4405 30.806 5.4985 31.064 ;
      RECT 5.6685 30.806 5.7265 31.064 ;
      RECT 5.8965 30.806 5.9545 31.064 ;
      RECT 6.1245 30.806 6.1825 31.064 ;
      RECT 6.3525 30.806 6.4105 31.064 ;
      RECT 6.5805 30.806 6.6385 31.064 ;
      RECT 6.8085 30.806 6.8665 31.064 ;
      RECT 7.0365 30.806 7.0945 31.064 ;
      RECT 7.2645 30.806 7.3225 31.064 ;
      RECT 7.4925 30.806 7.5505 31.064 ;
      RECT 7.7205 30.806 7.7785 31.064 ;
      RECT 8.8605 31.9685 8.9185 34.8145 ;
      RECT 9.0885 31.9685 9.1465 34.8145 ;
      RECT 9.3165 31.9685 9.3745 34.8145 ;
      RECT 2.0205 31.9725 2.0785 33.764 ;
      RECT 2.2485 31.9725 2.3065 33.764 ;
      RECT 2.4765 31.9725 2.5345 33.764 ;
      RECT 2.7045 31.9725 2.7625 33.764 ;
      RECT 2.9325 31.9725 2.9905 33.764 ;
      RECT 3.6165 31.9725 3.6745 35.4275 ;
      RECT 3.8445 31.9725 3.9025 35.43 ;
      RECT 4.0725 31.9725 4.1305 35.43 ;
      RECT 4.3005 31.9725 4.3585 35.43 ;
      RECT 4.5285 31.9725 4.5865 35.43 ;
      RECT 4.7565 31.9725 4.8145 35.43 ;
      RECT 4.9845 31.9725 5.0425 35.43 ;
      RECT 5.2125 31.9725 5.2705 35.43 ;
      RECT 5.4405 31.9725 5.4985 35.43 ;
      RECT 5.6685 31.9725 5.7265 35.43 ;
      RECT 5.8965 31.9725 5.9545 35.43 ;
      RECT 6.1245 31.9725 6.1825 35.43 ;
      RECT 6.3525 31.9725 6.4105 33.764 ;
      RECT 6.5805 31.9725 6.6385 33.764 ;
      RECT 2.3625 32.336 2.4205 34.416 ;
      RECT 2.5905 32.336 2.6485 34.416 ;
      RECT 3.0465 32.5405 3.1045 33.764 ;
      RECT 3.5025 32.5405 3.5605 33.764 ;
      RECT 6.8085 33.344 6.8665 34.8155 ;
      RECT 7.0365 33.344 7.0945 34.8155 ;
      RECT 7.2645 33.344 7.3225 34.8155 ;
      RECT 7.4925 33.344 7.5505 34.8155 ;
      RECT 7.7205 33.344 7.7785 34.8155 ;
      RECT 7.9485 33.344 8.0065 34.8145 ;
      RECT 8.1765 33.344 8.2345 34.8145 ;
      RECT 8.4045 33.344 8.4625 34.8145 ;
      RECT 8.6325 33.344 8.6905 34.8145 ;
      RECT 6.9225 34.921 6.9805 36.23 ;
      RECT 0.4245 35.072 0.4825 46.259 ;
      RECT 6.4665 37.617 6.5245 41.73 ;
      RECT 5.5545 37.705 5.6125 41.73 ;
      RECT 4.8705 37.738 4.9285 41.73 ;
      RECT 3.6165 41.8685 3.6745 42.3515 ;
      RECT 3.8445 41.8685 3.9025 42.3515 ;
      RECT 4.0725 41.8685 4.1305 42.3515 ;
      RECT 4.3005 41.8685 4.3585 42.3515 ;
      RECT 4.5285 41.8685 4.5865 42.3515 ;
      RECT 4.7565 41.8685 4.8145 42.3515 ;
      RECT 4.9845 41.8685 5.0425 42.3515 ;
      RECT 5.2125 41.8685 5.2705 42.3515 ;
      RECT 5.4405 41.8685 5.4985 42.3515 ;
      RECT 5.6685 41.8685 5.7265 42.3515 ;
      RECT 5.8965 41.8685 5.9545 42.3515 ;
      RECT 6.1245 41.8685 6.1825 42.3515 ;
      RECT 6.3525 41.8685 6.4105 42.3515 ;
      RECT 6.5805 41.8685 6.6385 42.3515 ;
      RECT 6.8085 41.8685 6.8665 42.3515 ;
      RECT 7.0365 41.8685 7.0945 42.3515 ;
      RECT 7.2645 41.8685 7.3225 42.3515 ;
      RECT 7.4925 41.8685 7.5505 42.3515 ;
      RECT 7.7205 41.8685 7.7785 42.3515 ;
      RECT 1.9065 42.5685 1.9645 44.504 ;
      RECT 2.0205 42.5685 2.0785 44.031 ;
      RECT 2.1345 42.5685 2.1925 44.504 ;
      RECT 2.3625 42.5685 2.4205 44.3885 ;
      RECT 2.5905 42.5685 2.6485 44.3885 ;
      RECT 2.8185 42.5685 2.8765 44.504 ;
      RECT 3.0465 42.5685 3.1045 44.504 ;
      RECT 3.5025 42.5685 3.5605 44.504 ;
      RECT 3.9585 42.923 4.0165 44.504 ;
      RECT 4.1865 42.923 4.2445 44.504 ;
      RECT 4.4145 42.923 4.4725 44.504 ;
      RECT 4.6425 42.923 4.7005 44.504 ;
      RECT 5.0985 42.923 5.1565 44.504 ;
      RECT 5.3265 42.923 5.3845 44.504 ;
      RECT 5.7825 42.923 5.8405 44.504 ;
      RECT 6.0105 42.923 6.0685 44.504 ;
      RECT 6.2385 42.923 6.2965 44.504 ;
      RECT 3.7305 42.958 3.7885 44.504 ;
      RECT 4.8705 42.958 4.9285 44.504 ;
      RECT 5.5545 42.958 5.6125 44.504 ;
      RECT 6.4665 42.958 6.5245 44.504 ;
      RECT 3.6165 43.046 3.6745 43.304 ;
      RECT 3.8445 43.046 3.9025 44.031 ;
      RECT 4.0725 43.046 4.1305 43.304 ;
      RECT 4.3005 43.046 4.3585 43.304 ;
      RECT 4.5285 43.046 4.5865 43.304 ;
      RECT 4.7565 43.046 4.8145 43.304 ;
      RECT 4.9845 43.046 5.0425 43.304 ;
      RECT 5.2125 43.046 5.2705 43.304 ;
      RECT 5.4405 43.046 5.4985 43.304 ;
      RECT 5.6685 43.046 5.7265 43.304 ;
      RECT 5.8965 43.046 5.9545 43.304 ;
      RECT 6.1245 43.046 6.1825 43.304 ;
      RECT 6.3525 43.046 6.4105 43.304 ;
      RECT 6.5805 43.046 6.6385 43.304 ;
      RECT 6.8085 43.046 6.8665 43.304 ;
      RECT 7.0365 43.046 7.0945 43.304 ;
      RECT 7.2645 43.046 7.3225 43.304 ;
      RECT 7.4925 43.046 7.5505 43.304 ;
      RECT 7.7205 43.046 7.7785 43.304 ;
      RECT 8.8605 44.2085 8.9185 47.0545 ;
      RECT 9.0885 44.2085 9.1465 47.0545 ;
      RECT 9.3165 44.2085 9.3745 47.0545 ;
      RECT 2.0205 44.2125 2.0785 46.004 ;
      RECT 2.2485 44.2125 2.3065 46.004 ;
      RECT 2.4765 44.2125 2.5345 46.004 ;
      RECT 2.7045 44.2125 2.7625 46.004 ;
      RECT 2.9325 44.2125 2.9905 46.004 ;
      RECT 3.6165 44.2125 3.6745 47.6675 ;
      RECT 3.8445 44.2125 3.9025 47.67 ;
      RECT 4.0725 44.2125 4.1305 47.67 ;
      RECT 4.3005 44.2125 4.3585 47.67 ;
      RECT 4.5285 44.2125 4.5865 47.67 ;
      RECT 4.7565 44.2125 4.8145 47.67 ;
      RECT 4.9845 44.2125 5.0425 47.67 ;
      RECT 5.2125 44.2125 5.2705 47.67 ;
      RECT 5.4405 44.2125 5.4985 47.67 ;
      RECT 5.6685 44.2125 5.7265 47.67 ;
      RECT 5.8965 44.2125 5.9545 47.67 ;
      RECT 6.1245 44.2125 6.1825 47.67 ;
      RECT 6.3525 44.2125 6.4105 46.004 ;
      RECT 6.5805 44.2125 6.6385 46.004 ;
      RECT 2.3625 44.576 2.4205 46.656 ;
      RECT 2.5905 44.576 2.6485 46.656 ;
      RECT 3.0465 44.7805 3.1045 46.004 ;
      RECT 3.5025 44.7805 3.5605 46.004 ;
      RECT 6.8085 45.584 6.8665 47.0555 ;
      RECT 7.0365 45.584 7.0945 47.0555 ;
      RECT 7.2645 45.584 7.3225 47.0555 ;
      RECT 7.4925 45.584 7.5505 47.0555 ;
      RECT 7.7205 45.584 7.7785 47.0555 ;
      RECT 7.9485 45.584 8.0065 47.0545 ;
      RECT 8.1765 45.584 8.2345 47.0545 ;
      RECT 8.4045 45.584 8.4625 47.0545 ;
      RECT 8.6325 45.584 8.6905 47.0545 ;
      RECT 6.9225 47.161 6.9805 48.47 ;
    LAYER M0 ;
      RECT MASK 1 0 0 10.26 48.96 ;
      RECT MASK 2 0 0 10.26 48.96 ;
  END
END dwc_ddrphy_pclk_master

END LIBRARY
