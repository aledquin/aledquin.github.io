# LEF OUT API 
# Creation Date : Mon Aug 23 12:52:49 PDT 2021
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_por
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_por 0 0 ;
  SYMMETRY X Y ;
  SIZE 37.32 BY 31.32 ;
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER D8 ;
        RECT 0.5 2.7125 36.69075 3.4125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 25.5125 36.69075 26.2125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 21.9125 36.69075 22.6125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 9.9125 36.69075 10.6125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 18.3125 36.69075 19.0125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 14.7125 36.69075 15.4125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 7.5125 36.69075 8.2125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 5.1125 36.69075 5.8125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 29.1125 36.69075 29.8125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 12.3125 36.69075 13.0125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 0.3125 36.69075 1.0125 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER D8 ;
        RECT 0.5 27.9125 36.69075 28.6125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 17.1125 36.69075 17.8125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 20.7125 36.69075 21.4125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 13.5125 36.69075 14.2125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 11.1125 36.69075 11.8125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 8.7125 36.69075 9.4125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 6.3125 36.69075 7.0125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 3.9125 36.69075 4.6125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 24.3125 36.69075 25.0125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 1.5125 36.69075 2.2125 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER D8 ;
        RECT 0.5 19.5125 36.69075 20.2125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 23.1125 36.69075 23.8125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5 15.9125 36.69075 16.6125 ;
    END
  END VDD
  PIN Reset_X
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11744 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.27864 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 367.049 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 525.889 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 36.06325 31.24 36.14325 31.32 ;
    END
  END Reset_X
  PIN SetDCTSanePulse
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11744 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.27864 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 370.429 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 529.487 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 35.52325 31.24 35.60325 31.32 ;
    END
  END SetDCTSanePulse
  PIN DFTDatSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11418 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.271305 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 368.284 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 523.604 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 34.56325 31.24 34.64325 31.32 ;
    END
  END DFTDatSel
  PIN DCTMemReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11396 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.27081 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002808 LAYER D6 ;
      ANTENNAMAXAREACAR 170.601 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 242.058 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.98325 31.24 34.06325 31.32 ;
    END
  END DCTMemReset
  PIN ClrPORMemReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11236 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26721 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 366.556 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 519.265 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.20325 31.24 33.28325 31.32 ;
    END
  END ClrPORMemReset
  PIN PwrOkDlyd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.49438 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.76317 LAYER D5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001944 LAYER D5 ;
      ANTENNAMAXAREACAR 2065.07 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 2473.42 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 0 27.13625 0.12 27.25625 ;
    END
  END PwrOkDlyd
  PIN PORMemReset
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3432 LAYER D5 ;
    ANTENNADIFFAREA 0.012636 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 37.2 27.741 37.32 27.861 ;
    END
  END PORMemReset
  PIN DCTSane
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.79328 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.29928 LAYER D5 ;
    ANTENNADIFFAREA 0.012636 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 37.24 28.39625 37.32 28.47625 ;
    END
  END DCTSane
  PIN PwrOkDlyd_VIO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7715 LAYER D6 ;
    ANTENNAPARTIALMETALAREA 1.76137 LAYER D7 ;
    ANTENNAPARTIALMETALAREA 19.1168 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.419175 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.578925 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 5.04176 LAYER D8 ;
    ANTENNAPARTIALCUTAREA 0.0512 LAYER S6 ;
    ANTENNAPARTIALCUTAREA 0.384 LAYER S7 ;
    ANTENNADIFFAREA 2.58048 LAYER D6 ;
    ANTENNADIFFAREA 2.58048 LAYER S6 ;
    ANTENNADIFFAREA 2.58048 LAYER D7 ;
    ANTENNADIFFAREA 2.58048 LAYER S7 ;
    ANTENNADIFFAREA 2.58048 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 6.02 30.3125 33.32975 31.0125 ;
    END
    PORT
      LAYER D6 ;
        RECT 18.9 31.02 19.3 31.32 ;
    END
  END PwrOkDlyd_VIO
  PIN MemResetLPullDown_VIO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61814 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.40521 LAYER D5 ;
    ANTENNADIFFAREA 0.48384 LAYER D5 ;
    PORT
      LAYER D5 ;
        RECT 37.24 22.37375 37.32 22.45375 ;
    END
  END MemResetLPullDown_VIO
  PIN MemResetLPullUp_VIO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.69685 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 4.06687 LAYER D6 ;
    ANTENNADIFFAREA 0.32256 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 24.71975 0 24.83975 0.12 ;
    END
  END MemResetLPullUp_VIO
  PIN PwrOk_VIO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.50782 LAYER D5 ;
    ANTENNAPARTIALMETALAREA 1.14979 LAYER D6 ;
    ANTENNAPARTIALMETALAREA 4.746 LAYER D7 ;
    ANTENNAPARTIALMETALAREA 19.1168 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1587 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8908199375 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3464 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 5.04176 LAYER D8 ;
    ANTENNAPARTIALCUTAREA 0.0384 LAYER S5 ;
    ANTENNAPARTIALCUTAREA 0.1536 LAYER S6 ;
    ANTENNAPARTIALCUTAREA 1.0752 LAYER S7 ;
    ANTENNADIFFAREA 2.58048 LAYER D5 ;
    ANTENNADIFFAREA 2.58048 LAYER S5 ;
    ANTENNADIFFAREA 2.58048 LAYER D6 ;
    ANTENNADIFFAREA 2.58048 LAYER S6 ;
    ANTENNADIFFAREA 2.58048 LAYER D7 ;
    ANTENNADIFFAREA 2.58048 LAYER S7 ;
    ANTENNADIFFAREA 2.58048 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 6.02 26.7125 33.32975 27.4125 ;
    END
    PORT
      LAYER D5 ;
        RECT 37.02 26.48525 37.32 26.78525 ;
    END
  END PwrOk_VIO
  PIN PwrOk_VMEMP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0966999375 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.231975 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 129.82499994 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 282.764 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 1.844 31.24 1.924 31.32 ;
    END
  END PwrOk_VMEMP
  OBS
    LAYER M1 SPACING 0 ;
      RECT 0 0 37.32 31.32 ;
    LAYER M2 SPACING 0 ;
      RECT 0 0 37.32 31.32 ;
    LAYER M3 SPACING 0 ;
      RECT 0 0 37.32 31.32 ;
    LAYER M4 SPACING 0 ;
      RECT 0 0 37.32 31.32 ;
    LAYER D5 SPACING 0 ;
      POLYGON 37.32 0 37.32 22.37375 37.24 22.37375 37.24 22.45375 37.32 22.45375 37.32 26.48525 37.02 26.48525 37.02 26.78525 37.32 26.78525 37.32 27.741 37.2 27.741 37.2 27.861 37.32 27.861 37.32 28.39625 37.24 28.39625 37.24 28.47625 37.32 28.47625 37.32 31.32 0 31.32 0 27.25625 0.12 27.25625 0.12 27.13625 0 27.13625 0 0 ;
    LAYER D6 SPACING 0 ;
      POLYGON 24.71975 0 24.71975 0.12 24.83975 0.12 24.83975 0 37.32 0 37.32 31.32 36.14325 31.32 36.14325 31.24 36.06325 31.24 36.06325 31.32 35.60325 31.32 35.60325 31.24 35.52325 31.24 35.52325 31.32 34.64325 31.32 34.64325 31.24 34.56325 31.24 34.56325 31.32 34.06325 31.32 34.06325 31.24 33.98325 31.24 33.98325 31.32 33.28325 31.32 33.28325 31.24 33.20325 31.24 33.20325 31.32 19.3 31.32 19.3 31.02 18.9 31.02 18.9 31.32 1.924 31.32 1.924 31.24 1.844 31.24 1.844 31.32 0 31.32 0 0 ;
    LAYER D7 SPACING 0 ;
      RECT 0 0 37.32 31.32 ;
  END
END dwc_ddrphy_por

END LIBRARY
