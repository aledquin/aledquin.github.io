# LEF OUT API 
# Creation Date : Wed Jul 15 16:43:29 PDT 2020
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_vrefglobal
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_vrefglobal 0 0 ;
  SYMMETRY X Y ;
  SIZE 130.416 BY 109.44 ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 0.2 10 130.199 10.45 ;
        RECT 0.2 5.2 130.199 5.65 ;
        RECT 0.2 0.4 130.199 0.85 ;
    END
  END VDD
  PIN VAA
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 0.2 108.03 130.216 108.48 ;
        RECT 0.2 106.43 130.216 106.88 ;
        RECT 0.2 104.83 130.216 105.28 ;
        RECT 0.2 103.23 130.216 103.68 ;
        RECT 0.2 101.63 130.216 102.08 ;
        RECT 0.2 100.03 130.216 100.48 ;
        RECT 0.2 98.43 130.216 98.88 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.2 83.6 130.199 84.05 ;
        RECT 0.2 80.4 130.199 80.85 ;
        RECT 0.2 77.2 130.199 77.65 ;
        RECT 0.2 74 130.199 74.45 ;
        RECT 0.2 70.8 130.199 71.25 ;
        RECT 0.2 67.6 130.199 68.05 ;
        RECT 0.2 64.4 130.199 64.85 ;
        RECT 0.2 61.2 130.199 61.65 ;
        RECT 0.2 58 130.199 58.45 ;
        RECT 0.2 54.8 130.199 55.25 ;
        RECT 0.2 51.6 130.199 52.05 ;
        RECT 0.2 48.4 130.199 48.85 ;
        RECT 0.2 45.2 130.199 45.65 ;
        RECT 0.2 42 130.199 42.45 ;
        RECT 0.2 38.8 130.199 39.25 ;
        RECT 0.2 35.6 130.199 36.05 ;
        RECT 0.2 32.4 130.199 32.85 ;
        RECT 0.2 29.2 130.199 29.65 ;
        RECT 0.2 26 130.199 26.45 ;
        RECT 0.2 22.8 130.199 23.25 ;
        RECT 0.2 19.6 130.199 20.05 ;
        RECT 0.2 16.4 130.199 16.85 ;
        RECT 0.2 13.2 130.199 13.65 ;
        RECT 0.2 8.4 130.199 8.85 ;
        RECT 0.2 3.6 130.199 4.05 ;
    END
  END VAA
  PIN Csr_VrefDAC[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5632 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0412 LAYER M5 ;
      ANTENNAMAXAREACAR 425.115 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 0.9915 109.36 1.0715 109.44 ;
    END
  END Csr_VrefDAC[6]
  PIN Csr_VrefDAC[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5055999375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0412 LAYER M5 ;
      ANTENNAMAXAREACAR 408.598 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.1515 109.36 1.2315 109.44 ;
    END
  END Csr_VrefDAC[5]
  PIN Csr_VrefDAC[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5504 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0412 LAYER M5 ;
      ANTENNAMAXAREACAR 421.124 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.7325 109.36 1.8125 109.44 ;
    END
  END Csr_VrefDAC[4]
  PIN AnalogIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.308 LAYER M5 ;
    ANTENNADIFFAREA 1.62582 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 5.4375 109.36 5.5175 109.44 ;
    END
  END AnalogIn
  PIN Csr_VrefDAC[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4928 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0412 LAYER M5 ;
      ANTENNAMAXAREACAR 422.496 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 2.4735 109.36 2.5535 109.44 ;
    END
  END Csr_VrefDAC[2]
  PIN Csr_VrefDAC[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.448 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0412 LAYER M5 ;
      ANTENNAMAXAREACAR 416.458 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 2.6335 109.36 2.7135 109.44 ;
    END
  END Csr_VrefDAC[1]
  PIN Csr_VrefDAC[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.608 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0412 LAYER M5 ;
      ANTENNAMAXAREACAR 415.331 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 3.2145 109.36 3.2945 109.44 ;
    END
  END Csr_VrefDAC[0]
  PIN Csr_VrefDAC[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4352 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0412 LAYER M5 ;
      ANTENNAMAXAREACAR 406.733 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 1.8925 109.36 1.9725 109.44 ;
    END
  END Csr_VrefDAC[3]
  PIN Csr_VrefMode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6208 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.014112 LAYER M5 ;
      ANTENNAMAXAREACAR 897.482 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 3.3745 109.36 3.4545 109.44 ;
    END
  END Csr_VrefMode[2]
  PIN Csr_VrefMode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6656 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.014112 LAYER M5 ;
      ANTENNAMAXAREACAR 892.541 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 3.9555 109.36 4.0355 109.44 ;
    END
  END Csr_VrefMode[1]
  PIN Csr_VrefMode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6784 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.014112 LAYER M5 ;
      ANTENNAMAXAREACAR 891.19 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 4.1155 109.36 4.1955 109.44 ;
    END
  END Csr_VrefMode[0]
  PIN PwrOk_VIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3775999375 LAYER M5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.040032 LAYER M5 ;
      ANTENNAMAXAREACAR 297.493 LAYER M5 ;
    PORT
      LAYER M5 ;
        RECT 4.6965 109.36 4.7765 109.44 ;
    END
  END PwrOk_VIO
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M8 ;
        RECT 107.51 94.455 130.199 94.905 ;
        RECT 0.2 94.455 23.817 94.905 ;
        RECT 107.51 92.9 130.199 93.35 ;
        RECT 0.2 92.9 23.817 93.35 ;
        RECT 107.51 91.345 130.199 91.795 ;
        RECT 0.2 91.345 23.817 91.795 ;
        RECT 107.51 89.79 130.199 90.24 ;
        RECT 0.2 89.79 23.817 90.24 ;
        RECT 107.51 88.26 130.199 88.71 ;
        RECT 0.2 88.26 8.997 88.71 ;
        RECT 107.51 86.79 130.199 87.24 ;
        RECT 0.2 86.79 23.817 87.24 ;
        RECT 0.2 84.4 130.199 84.85 ;
        RECT 0.2 82.8 130.199 83.25 ;
        RECT 0.2 81.2 130.199 81.65 ;
        RECT 0.2 79.6 130.199 80.05 ;
        RECT 0.2 78 130.199 78.45 ;
        RECT 0.2 76.4 130.199 76.85 ;
        RECT 0.2 74.8 130.199 75.25 ;
        RECT 0.2 73.2 130.199 73.65 ;
        RECT 0.2 71.6 130.199 72.05 ;
        RECT 0.2 70 130.199 70.45 ;
        RECT 0.2 68.4 130.199 68.85 ;
        RECT 0.2 66.8 130.199 67.25 ;
        RECT 0.2 65.2 130.199 65.65 ;
        RECT 0.2 63.6 130.199 64.05 ;
        RECT 0.2 62 130.199 62.45 ;
        RECT 0.2 60.4 130.199 60.85 ;
        RECT 0.2 58.8 130.199 59.25 ;
        RECT 0.2 57.2 130.199 57.65 ;
        RECT 0.2 55.6 130.199 56.05 ;
        RECT 0.2 54 130.199 54.45 ;
        RECT 0.2 52.4 130.199 52.85 ;
        RECT 0.2 50.8 130.199 51.25 ;
        RECT 0.2 49.2 130.199 49.65 ;
        RECT 0.2 47.6 130.199 48.05 ;
        RECT 0.2 46 130.199 46.45 ;
        RECT 0.2 44.4 130.199 44.85 ;
        RECT 0.2 42.8 130.199 43.25 ;
        RECT 0.2 41.2 130.199 41.65 ;
        RECT 0.2 39.6 130.199 40.05 ;
        RECT 0.2 38 130.199 38.45 ;
        RECT 0.2 36.4 130.199 36.85 ;
        RECT 0.2 34.8 130.199 35.25 ;
        RECT 0.2 33.2 130.199 33.65 ;
        RECT 0.2 31.6 130.199 32.05 ;
        RECT 0.2 30 130.199 30.45 ;
        RECT 0.2 28.4 130.199 28.85 ;
        RECT 0.2 26.8 130.199 27.25 ;
        RECT 0.2 25.2 130.199 25.65 ;
        RECT 0.2 23.6 130.199 24.05 ;
        RECT 0.2 22 130.199 22.45 ;
        RECT 0.2 20.4 130.199 20.85 ;
        RECT 0.2 18.8 130.199 19.25 ;
        RECT 0.2 17.2 130.199 17.65 ;
        RECT 0.2 15.6 130.199 16.05 ;
        RECT 0.2 14 130.199 14.45 ;
        RECT 0.2 12.4 130.199 12.85 ;
        RECT 0.2 10.8 130.199 11.25 ;
        RECT 0.2 9.2 130.199 9.65 ;
        RECT 0.2 7.6 130.199 8.05 ;
        RECT 0.2 6 130.199 6.45 ;
        RECT 0.2 4.4 130.199 4.85 ;
        RECT 0.2 2.8 130.199 3.25 ;
        RECT 0.2 1.2 130.199 1.65 ;
    END
    PORT
      LAYER M8 ;
        RECT 69.796 94.19 107.057 94.69 ;
        RECT 69.796 92.39 107.057 92.89 ;
        RECT 69.796 90.59 107.057 91.09 ;
        RECT 69.796 88.79 107.057 89.29 ;
        RECT 69.796 86.99 107.057 87.49 ;
    END
    PORT
      LAYER M8 ;
        RECT 0.2 108.83 130.216 109.28 ;
        RECT 0.2 107.23 130.216 107.68 ;
        RECT 0.2 105.63 130.216 106.08 ;
        RECT 0.2 104.03 130.216 104.48 ;
        RECT 0.2 102.43 130.216 102.88 ;
        RECT 0.2 100.83 130.216 101.28 ;
        RECT 0.2 99.23 130.216 99.68 ;
        RECT 0.2 97.63 130.216 98.08 ;
        RECT 0.2 96.03 130.216 96.48 ;
    END
  END VSS
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M8 ;
        RECT 0.2 96.83 130.199 97.28 ;
        RECT 107.51 95.255 130.199 95.705 ;
        RECT 0.2 95.255 23.817 95.705 ;
        RECT 107.51 93.655 130.199 94.105 ;
        RECT 0.2 93.655 23.817 94.105 ;
        RECT 107.51 92.1 130.199 92.55 ;
        RECT 0.2 92.1 23.817 92.55 ;
        RECT 107.51 90.545 130.199 90.995 ;
        RECT 0.2 90.545 23.817 90.995 ;
        RECT 107.51 89.07 130.199 89.52 ;
        RECT 0.2 89.07 8.997 89.52 ;
        RECT 107.51 87.54 130.199 87.99 ;
        RECT 0.2 87.54 23.817 87.99 ;
        RECT 107.51 86.075 130.199 86.525 ;
        RECT 0.2 86.075 8.997 86.525 ;
        RECT 0.2 85.2 130.199 85.65 ;
        RECT 0.2 82 130.199 82.45 ;
        RECT 0.2 78.8 130.199 79.25 ;
        RECT 0.2 75.6 130.199 76.05 ;
        RECT 0.2 72.4 130.199 72.85 ;
        RECT 0.2 69.2 130.199 69.65 ;
        RECT 0.2 66 130.199 66.45 ;
        RECT 0.2 62.8 130.199 63.25 ;
        RECT 0.2 59.6 130.199 60.05 ;
        RECT 0.2 56.4 130.199 56.85 ;
        RECT 0.2 53.2 130.199 53.65 ;
        RECT 0.2 50 130.199 50.45 ;
        RECT 0.2 46.8 130.199 47.25 ;
        RECT 0.2 43.6 130.199 44.05 ;
        RECT 0.2 40.4 130.199 40.85 ;
        RECT 0.2 37.2 130.199 37.65 ;
        RECT 0.2 34 130.199 34.45 ;
        RECT 0.2 30.8 130.199 31.25 ;
        RECT 0.2 27.6 130.199 28.05 ;
        RECT 0.2 24.4 130.199 24.85 ;
        RECT 0.2 21.2 130.199 21.65 ;
        RECT 0.2 18 130.199 18.45 ;
        RECT 0.2 14.8 130.199 15.25 ;
        RECT 0.2 11.6 130.199 12.05 ;
        RECT 0.2 6.8 130.199 7.25 ;
        RECT 0.2 2 130.199 2.45 ;
    END
    PORT
      LAYER M8 ;
        RECT 24.017 94.19 69.396 94.69 ;
        RECT 24.017 92.39 69.396 92.89 ;
        RECT 103.27 91.49 107.057 91.99 ;
        RECT 24.017 90.59 69.396 91.09 ;
        RECT 103.27 89.69 107.057 90.19 ;
        RECT 24.017 88.79 69.396 89.29 ;
        RECT 103.27 87.89 107.057 88.39 ;
    END
    PORT
      LAYER M8 ;
        RECT 103.27 93.29 107.057 93.79 ;
    END
    PORT
      LAYER M8 ;
        RECT 24.017 86.99 69.396 87.49 ;
    END
  END VDDQ
  PIN VrefPAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 157.706 LAYER M8 ;
    ANTENNADIFFAREA 54.7621 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 50.4166 LAYER M8 ;
      ANTENNAMAXAREACAR 19.171 LAYER M8 ;
    PORT
      LAYER M8 ;
        RECT 24.017 91.49 102.87 91.99 ;
        RECT 24.017 89.69 102.87 90.19 ;
        RECT 24.017 87.89 102.87 88.39 ;
    END
    PORT
      LAYER M8 ;
        RECT 24.017 93.29 102.87 93.79 ;
    END
  END VrefPAD
  PIN VrefOut
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9945 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 21.693 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.5472 LAYER VIA7 ;
    ANTENNADIFFAREA 66.1865 LAYER M7 ;
    ANTENNADIFFAREA 66.1865 LAYER VIA7 ;
    ANTENNADIFFAREA 66.1865 LAYER M8 ;
    PORT
      LAYER M8 ;
        RECT 9.355 89.07 23.817 89.57 ;
        RECT 9.355 88.21 23.817 88.71 ;
        RECT 9.355 86.05 23.817 86.55 ;
    END
    PORT
      LAYER M7 ;
        RECT 15.403 108.99 15.853 109.44 ;
    END
  END VrefOut
  OBS
    LAYER M1 SPACING 0 ;
      RECT 0 0 130.416 109.44 ;
      RECT MASK 1 58.765 0.6 58.825 1.378 ;
      RECT MASK 1 59.223 0.6 59.283 1.378 ;
      RECT MASK 1 59.681 0.6 59.741 1.378 ;
      RECT MASK 1 60.2275 0.6 60.2875 2.2375 ;
      RECT MASK 1 63.803 0.6 63.863 1.378 ;
      RECT MASK 1 64.261 0.6 64.321 1.378 ;
      RECT MASK 1 64.719 0.6 64.779 1.378 ;
      RECT MASK 1 65.635 0.6 65.695 1.5175 ;
      RECT MASK 1 65.864 0.6 65.924 1.5175 ;
      RECT MASK 1 58.307 0.605 58.367 0.835 ;
      RECT MASK 1 58.994 0.605 59.054 0.835 ;
      RECT MASK 1 59.452 0.605 59.512 0.835 ;
      RECT MASK 1 59.91 0.605 59.97 0.835 ;
      RECT MASK 1 60.826 0.605 60.886 0.835 ;
      RECT MASK 1 61.284 0.605 61.344 0.835 ;
      RECT MASK 1 61.513 0.605 61.573 0.835 ;
      RECT MASK 1 61.742 0.605 61.802 0.835 ;
      RECT MASK 1 61.971 0.605 62.031 0.835 ;
      RECT MASK 1 62.2 0.605 62.26 0.835 ;
      RECT MASK 1 62.429 0.605 62.489 0.835 ;
      RECT MASK 1 62.658 0.605 62.718 0.835 ;
      RECT MASK 1 62.887 0.605 62.947 0.835 ;
      RECT MASK 1 63.116 0.605 63.176 0.835 ;
      RECT MASK 1 63.345 0.605 63.405 0.835 ;
      RECT MASK 1 64.49 0.605 64.55 0.835 ;
      RECT MASK 1 64.948 0.605 65.008 0.835 ;
      RECT MASK 1 65.177 0.605 65.237 0.835 ;
      RECT MASK 1 65.406 0.605 65.466 0.835 ;
      RECT MASK 1 46.2405 0.684 46.2805 3.061 ;
      RECT MASK 1 45.8405 0.984 45.8805 3.2295 ;
      RECT MASK 1 50.4095 1.005 50.4495 1.426 ;
      RECT MASK 1 51.0735 1.005 51.1135 1.426 ;
      RECT MASK 1 51.7375 1.005 51.7775 1.426 ;
      RECT MASK 1 52.4015 1.005 52.4415 1.426 ;
      RECT MASK 1 49.9665 1.02 50.0065 1.76 ;
      RECT MASK 1 50.6305 1.02 50.6705 1.76 ;
      RECT MASK 1 51.2945 1.02 51.3345 1.76 ;
      RECT MASK 1 51.9585 1.02 51.9985 1.76 ;
      RECT MASK 1 52.6225 1.02 52.6625 1.76 ;
      RECT MASK 1 52.1795 1.1 52.2195 1.426 ;
      RECT MASK 1 60.826 1.16 60.886 2.315 ;
      RECT MASK 1 61.284 1.16 61.344 1.378 ;
      RECT MASK 1 61.742 1.16 61.802 1.378 ;
      RECT MASK 1 62.2 1.16 62.26 1.378 ;
      RECT MASK 1 62.658 1.16 62.718 1.378 ;
      RECT MASK 1 63.116 1.16 63.176 2.315 ;
      RECT MASK 1 115.44 1.31 115.54 24.01 ;
      RECT MASK 1 128.886 1.31 128.986 24.01 ;
      RECT MASK 1 61.284 1.498 61.344 1.881 ;
      RECT MASK 1 61.742 1.498 61.802 1.881 ;
      RECT MASK 1 3.0905 1.53 3.1505 2.046 ;
      RECT MASK 1 3.3195 1.53 3.3795 2.308 ;
      RECT MASK 1 3.7775 1.53 3.8375 2.308 ;
      RECT MASK 1 4.2355 1.53 4.2955 2.308 ;
      RECT MASK 1 4.6935 1.53 4.7535 2.308 ;
      RECT MASK 1 5.1515 1.53 5.2115 2.309 ;
      RECT MASK 1 5.3805 1.53 5.4405 2.046 ;
      RECT MASK 1 5.6095 1.53 5.6695 2.308 ;
      RECT MASK 1 6.5255 1.53 6.5855 2.308 ;
      RECT MASK 1 7.4415 1.53 7.5015 2.308 ;
      RECT MASK 1 8.3575 1.53 8.4175 2.3075 ;
      RECT MASK 1 8.5865 1.53 8.6465 2.046 ;
      RECT MASK 1 9.9605 1.53 10.0205 2.046 ;
      RECT MASK 1 14.3445 1.53 14.4045 7.89 ;
      RECT MASK 1 14.5735 1.53 14.6335 2.308 ;
      RECT MASK 1 15.0315 1.53 15.0915 2.308 ;
      RECT MASK 1 15.4895 1.53 15.5495 2.308 ;
      RECT MASK 1 15.9475 1.53 16.0075 2.308 ;
      RECT MASK 1 16.4055 1.53 16.4655 2.308 ;
      RECT MASK 1 16.8635 1.53 16.9235 2.308 ;
      RECT MASK 1 17.3215 1.53 17.3815 2.308 ;
      RECT MASK 1 17.7795 1.53 17.8395 2.308 ;
      RECT MASK 1 18.2375 1.53 18.2975 2.308 ;
      RECT MASK 1 18.6955 1.53 18.7555 2.308 ;
      RECT MASK 1 19.1535 1.53 19.2135 2.308 ;
      RECT MASK 1 19.6115 1.53 19.6715 2.308 ;
      RECT MASK 1 20.0695 1.53 20.1295 2.308 ;
      RECT MASK 1 20.5275 1.53 20.5875 2.308 ;
      RECT MASK 1 20.9855 1.53 21.0455 2.308 ;
      RECT MASK 1 21.4435 1.53 21.5035 2.308 ;
      RECT MASK 1 21.6725 1.53 21.7325 7.89 ;
      RECT MASK 1 25.2045 1.53 25.2645 7.89 ;
      RECT MASK 1 25.4335 1.53 25.4935 2.308 ;
      RECT MASK 1 25.8915 1.53 25.9515 2.308 ;
      RECT MASK 1 26.3495 1.53 26.4095 2.308 ;
      RECT MASK 1 26.8075 1.53 26.8675 2.308 ;
      RECT MASK 1 27.2655 1.53 27.3255 2.308 ;
      RECT MASK 1 27.7235 1.53 27.7835 2.308 ;
      RECT MASK 1 28.1815 1.53 28.2415 2.308 ;
      RECT MASK 1 28.6395 1.53 28.6995 2.308 ;
      RECT MASK 1 29.0975 1.53 29.1575 2.308 ;
      RECT MASK 1 29.5555 1.53 29.6155 2.308 ;
      RECT MASK 1 30.0135 1.53 30.0735 2.308 ;
      RECT MASK 1 30.4715 1.53 30.5315 2.308 ;
      RECT MASK 1 30.9295 1.53 30.9895 2.308 ;
      RECT MASK 1 31.3875 1.53 31.4475 2.308 ;
      RECT MASK 1 31.8455 1.53 31.9055 2.308 ;
      RECT MASK 1 32.3035 1.53 32.3635 2.308 ;
      RECT MASK 1 32.5325 1.53 32.5925 7.89 ;
      RECT MASK 1 36.9165 1.53 36.9765 2.046 ;
      RECT MASK 1 38.2905 1.53 38.3505 2.046 ;
      RECT MASK 1 38.5195 1.53 38.5795 2.3075 ;
      RECT MASK 1 39.4355 1.53 39.4955 2.308 ;
      RECT MASK 1 40.3515 1.53 40.4115 2.308 ;
      RECT MASK 1 41.2675 1.53 41.3275 2.308 ;
      RECT MASK 1 41.4965 1.53 41.5565 2.046 ;
      RECT MASK 1 41.7255 1.53 41.7855 2.309 ;
      RECT MASK 1 42.1835 1.53 42.2435 2.308 ;
      RECT MASK 1 42.6415 1.53 42.7015 2.308 ;
      RECT MASK 1 43.0995 1.53 43.1595 2.308 ;
      RECT MASK 1 43.5575 1.53 43.6175 2.308 ;
      RECT MASK 1 43.7865 1.53 43.8465 2.046 ;
      RECT MASK 1 50.4095 1.5925 50.4495 2.155 ;
      RECT MASK 1 51.0735 1.5925 51.1135 2.155 ;
      RECT MASK 1 51.7375 1.5925 51.7775 2.155 ;
      RECT MASK 1 52.4015 1.5925 52.4415 2.155 ;
      RECT MASK 1 50.1905 1.5945 50.2245 2.115 ;
      RECT MASK 1 50.8545 1.5945 50.8885 2.115 ;
      RECT MASK 1 51.5185 1.5945 51.5525 2.115 ;
      RECT MASK 1 52.1825 1.5945 52.2165 2.115 ;
      RECT MASK 1 58.765 1.599 58.825 1.881 ;
      RECT MASK 1 59.223 1.599 59.283 1.881 ;
      RECT MASK 1 59.681 1.599 59.741 1.881 ;
      RECT MASK 1 62.2 1.599 62.26 1.982 ;
      RECT MASK 1 62.658 1.599 62.718 1.982 ;
      RECT MASK 1 63.803 1.599 63.863 1.881 ;
      RECT MASK 1 64.261 1.599 64.321 1.881 ;
      RECT MASK 1 64.719 1.599 64.779 1.881 ;
      RECT MASK 1 116.154 1.66 116.214 23.64 ;
      RECT MASK 1 128.21 1.66 128.27 23.64 ;
      RECT MASK 1 116.428 1.68 116.488 23.64 ;
      RECT MASK 1 116.702 1.68 116.762 23.64 ;
      RECT MASK 1 116.976 1.68 117.036 23.64 ;
      RECT MASK 1 117.25 1.68 117.31 23.64 ;
      RECT MASK 1 117.524 1.68 117.584 23.64 ;
      RECT MASK 1 117.798 1.68 117.858 23.64 ;
      RECT MASK 1 118.072 1.68 118.132 23.64 ;
      RECT MASK 1 118.346 1.68 118.406 23.64 ;
      RECT MASK 1 118.62 1.68 118.68 23.64 ;
      RECT MASK 1 118.894 1.68 118.954 23.64 ;
      RECT MASK 1 119.168 1.68 119.228 23.64 ;
      RECT MASK 1 119.442 1.68 119.502 23.64 ;
      RECT MASK 1 119.716 1.68 119.776 23.64 ;
      RECT MASK 1 119.99 1.68 120.05 23.64 ;
      RECT MASK 1 120.264 1.68 120.324 23.64 ;
      RECT MASK 1 120.538 1.68 120.598 23.64 ;
      RECT MASK 1 120.812 1.68 120.872 23.64 ;
      RECT MASK 1 121.086 1.68 121.146 23.64 ;
      RECT MASK 1 121.36 1.68 121.42 23.64 ;
      RECT MASK 1 121.634 1.68 121.694 23.64 ;
      RECT MASK 1 121.908 1.68 121.968 23.64 ;
      RECT MASK 1 122.182 1.68 122.242 23.64 ;
      RECT MASK 1 122.456 1.68 122.516 23.64 ;
      RECT MASK 1 122.73 1.68 122.79 23.64 ;
      RECT MASK 1 123.004 1.68 123.064 23.64 ;
      RECT MASK 1 123.278 1.68 123.338 23.64 ;
      RECT MASK 1 123.552 1.68 123.612 23.64 ;
      RECT MASK 1 123.826 1.68 123.886 23.64 ;
      RECT MASK 1 124.1 1.68 124.16 23.64 ;
      RECT MASK 1 124.374 1.68 124.434 23.64 ;
      RECT MASK 1 124.648 1.68 124.708 23.64 ;
      RECT MASK 1 124.922 1.68 124.982 23.64 ;
      RECT MASK 1 125.196 1.68 125.256 23.64 ;
      RECT MASK 1 125.47 1.68 125.53 23.64 ;
      RECT MASK 1 125.744 1.68 125.804 23.64 ;
      RECT MASK 1 126.018 1.68 126.078 23.64 ;
      RECT MASK 1 126.292 1.68 126.352 23.64 ;
      RECT MASK 1 126.566 1.68 126.626 23.64 ;
      RECT MASK 1 126.84 1.68 126.9 23.64 ;
      RECT MASK 1 127.114 1.68 127.174 23.64 ;
      RECT MASK 1 127.388 1.68 127.448 23.64 ;
      RECT MASK 1 127.662 1.68 127.722 23.64 ;
      RECT MASK 1 127.936 1.68 127.996 23.64 ;
      RECT MASK 1 49.3445 1.805 49.4045 3.725 ;
      RECT MASK 1 22.3385 1.815 22.3985 2.349 ;
      RECT MASK 1 22.5385 1.815 22.5985 2.44 ;
      RECT MASK 1 22.7385 1.815 22.7985 2.44 ;
      RECT MASK 1 22.9385 1.815 22.9985 2.44 ;
      RECT MASK 1 23.1385 1.815 23.1985 2.349 ;
      RECT MASK 1 23.7385 1.815 23.7985 2.349 ;
      RECT MASK 1 23.9385 1.815 23.9985 2.44 ;
      RECT MASK 1 24.1385 1.815 24.1985 2.44 ;
      RECT MASK 1 24.3385 1.815 24.3985 2.44 ;
      RECT MASK 1 24.5385 1.815 24.5985 2.349 ;
      RECT MASK 1 46.8405 1.955 46.8805 2.21 ;
      RECT MASK 1 47.0405 1.955 47.0805 2.202 ;
      RECT MASK 1 47.2405 1.955 47.2805 2.21 ;
      RECT MASK 1 47.4405 1.955 47.4805 2.21 ;
      RECT MASK 1 47.6405 1.955 47.6805 2.202 ;
      RECT MASK 1 47.8405 1.955 47.8805 2.21 ;
      RECT MASK 1 48.0405 1.955 48.0805 2.21 ;
      RECT MASK 1 48.2405 1.955 48.2805 2.21 ;
      RECT MASK 1 48.4405 1.955 48.4805 2.21 ;
      RECT MASK 1 48.6405 1.955 48.6805 2.33 ;
      RECT MASK 1 48.8405 1.955 48.8805 2.21 ;
      RECT MASK 1 49.0405 1.955 49.0805 2.21 ;
      RECT MASK 1 49.9665 1.955 50.0065 6.57 ;
      RECT MASK 1 50.6305 1.955 50.6705 6.57 ;
      RECT MASK 1 51.2945 1.955 51.3345 6.57 ;
      RECT MASK 1 51.9585 1.955 51.9985 6.57 ;
      RECT MASK 1 52.6225 1.955 52.6625 6.57 ;
      RECT MASK 1 65.635 2.0825 65.695 3.138 ;
      RECT MASK 1 9.5025 2.09 9.5625 2.308 ;
      RECT MASK 1 37.3745 2.09 37.4345 2.308 ;
      RECT MASK 1 6.2965 2.095 6.3565 2.912 ;
      RECT MASK 1 40.5805 2.095 40.6405 2.912 ;
      RECT MASK 1 58.765 2.102 58.825 2.602 ;
      RECT MASK 1 59.223 2.102 59.283 2.602 ;
      RECT MASK 1 59.681 2.102 59.741 2.602 ;
      RECT MASK 1 61.284 2.102 61.344 2.315 ;
      RECT MASK 1 61.742 2.102 61.802 2.315 ;
      RECT MASK 1 62.2 2.102 62.26 2.315 ;
      RECT MASK 1 62.658 2.102 62.718 2.315 ;
      RECT MASK 1 63.803 2.102 63.863 2.602 ;
      RECT MASK 1 64.261 2.102 64.321 2.602 ;
      RECT MASK 1 64.719 2.102 64.779 2.602 ;
      RECT MASK 1 2.4035 2.128 2.4635 3.212 ;
      RECT MASK 1 2.8615 2.128 2.9215 3.212 ;
      RECT MASK 1 3.5485 2.128 3.6085 3.212 ;
      RECT MASK 1 4.0065 2.128 4.0665 2.405 ;
      RECT MASK 1 4.4645 2.128 4.5245 3.212 ;
      RECT MASK 1 4.9225 2.128 4.9825 3.212 ;
      RECT MASK 1 6.0675 2.128 6.1275 3.212 ;
      RECT MASK 1 6.9835 2.128 7.0435 3.212 ;
      RECT MASK 1 7.8995 2.128 7.9595 3.212 ;
      RECT MASK 1 8.8155 2.128 8.8755 2.65 ;
      RECT MASK 1 9.0445 2.128 9.1045 2.405 ;
      RECT MASK 1 9.2735 2.128 9.3335 2.65 ;
      RECT MASK 1 9.7315 2.128 9.7915 2.645 ;
      RECT MASK 1 11.3455 2.128 11.4055 3.212 ;
      RECT MASK 1 11.8035 2.128 11.8635 3.212 ;
      RECT MASK 1 12.2615 2.128 12.3215 3.212 ;
      RECT MASK 1 12.7195 2.128 12.7795 3.212 ;
      RECT MASK 1 34.1575 2.128 34.2175 3.212 ;
      RECT MASK 1 34.6155 2.128 34.6755 3.212 ;
      RECT MASK 1 35.0735 2.128 35.1335 3.212 ;
      RECT MASK 1 35.5315 2.128 35.5915 3.212 ;
      RECT MASK 1 37.1455 2.128 37.2055 2.645 ;
      RECT MASK 1 37.6035 2.128 37.6635 2.65 ;
      RECT MASK 1 37.8325 2.128 37.8925 2.405 ;
      RECT MASK 1 38.0615 2.128 38.1215 2.65 ;
      RECT MASK 1 38.9775 2.128 39.0375 3.212 ;
      RECT MASK 1 39.8935 2.128 39.9535 3.212 ;
      RECT MASK 1 40.8095 2.128 40.8695 3.212 ;
      RECT MASK 1 41.9545 2.128 42.0145 3.212 ;
      RECT MASK 1 42.4125 2.128 42.4725 3.212 ;
      RECT MASK 1 42.8705 2.128 42.9305 2.405 ;
      RECT MASK 1 43.3285 2.128 43.3885 3.212 ;
      RECT MASK 1 44.0155 2.128 44.0755 3.212 ;
      RECT MASK 1 44.4735 2.128 44.5335 3.212 ;
      RECT MASK 1 47.0405 2.24 47.0805 2.5 ;
      RECT MASK 1 47.6405 2.24 47.6805 2.5 ;
      RECT MASK 1 5.3805 2.33 5.4405 2.912 ;
      RECT MASK 1 41.4965 2.33 41.5565 2.912 ;
      RECT MASK 1 8.5865 2.335 8.6465 3.005 ;
      RECT MASK 1 10.8455 2.335 10.9055 3.01 ;
      RECT MASK 1 36.0315 2.335 36.0915 3.01 ;
      RECT MASK 1 38.2905 2.335 38.3505 3.005 ;
      RECT MASK 1 48.4405 2.41 48.4805 2.93 ;
      RECT MASK 1 7.2125 2.428 7.2725 2.912 ;
      RECT MASK 1 39.6645 2.428 39.7245 2.912 ;
      RECT MASK 1 61.971 2.43 62.031 2.9575 ;
      RECT MASK 1 61.055 2.435 61.115 3.6775 ;
      RECT MASK 1 58.536 2.438 58.596 2.938 ;
      RECT MASK 1 58.994 2.438 59.054 2.938 ;
      RECT MASK 1 59.452 2.438 59.512 2.938 ;
      RECT MASK 1 59.91 2.438 59.97 2.938 ;
      RECT MASK 1 60.368 2.438 60.428 2.938 ;
      RECT MASK 1 50.4095 2.457 50.4495 3.166 ;
      RECT MASK 1 51.0735 2.457 51.1135 3.166 ;
      RECT MASK 1 51.7375 2.457 51.7775 3.166 ;
      RECT MASK 1 52.4015 2.457 52.4415 3.166 ;
      RECT MASK 1 23.7385 2.469 23.7985 2.667 ;
      RECT MASK 1 12.9915 2.47 13.0515 2.65 ;
      RECT MASK 1 14.688 2.47 14.748 2.65 ;
      RECT MASK 1 15.146 2.47 15.206 2.65 ;
      RECT MASK 1 15.604 2.47 15.664 2.65 ;
      RECT MASK 1 16.062 2.47 16.122 2.65 ;
      RECT MASK 1 16.52 2.47 16.58 2.65 ;
      RECT MASK 1 16.978 2.47 17.038 2.65 ;
      RECT MASK 1 17.436 2.47 17.496 2.65 ;
      RECT MASK 1 18.352 2.47 18.412 2.65 ;
      RECT MASK 1 18.81 2.47 18.87 2.65 ;
      RECT MASK 1 19.726 2.47 19.786 2.65 ;
      RECT MASK 1 20.642 2.47 20.702 2.65 ;
      RECT MASK 1 21.1 2.47 21.16 2.65 ;
      RECT MASK 1 25.777 2.47 25.837 2.65 ;
      RECT MASK 1 26.235 2.47 26.295 2.65 ;
      RECT MASK 1 27.151 2.47 27.211 2.65 ;
      RECT MASK 1 28.067 2.47 28.127 2.65 ;
      RECT MASK 1 28.525 2.47 28.585 2.65 ;
      RECT MASK 1 29.441 2.47 29.501 2.65 ;
      RECT MASK 1 29.899 2.47 29.959 2.65 ;
      RECT MASK 1 30.357 2.47 30.417 2.65 ;
      RECT MASK 1 30.815 2.47 30.875 2.65 ;
      RECT MASK 1 31.273 2.47 31.333 2.65 ;
      RECT MASK 1 31.731 2.47 31.791 2.65 ;
      RECT MASK 1 32.189 2.47 32.249 2.65 ;
      RECT MASK 1 33.8855 2.47 33.9455 2.65 ;
      RECT MASK 1 23.1385 2.484 23.1985 2.6895 ;
      RECT MASK 1 9.9815 2.529 10.0415 2.765 ;
      RECT MASK 1 11.0955 2.529 11.1555 2.77 ;
      RECT MASK 1 35.7815 2.529 35.8415 2.77 ;
      RECT MASK 1 36.8955 2.529 36.9555 2.765 ;
      RECT MASK 1 46.8405 2.53 46.8805 2.93 ;
      RECT MASK 1 47.2405 2.53 47.2805 2.93 ;
      RECT MASK 1 47.4405 2.53 47.4805 2.93 ;
      RECT MASK 1 47.8405 2.53 47.8805 2.93 ;
      RECT MASK 1 48.0405 2.53 48.0805 2.93 ;
      RECT MASK 1 48.2405 2.53 48.2805 2.93 ;
      RECT MASK 1 48.6405 2.53 48.6805 2.93 ;
      RECT MASK 1 48.8405 2.53 48.8805 2.93 ;
      RECT MASK 1 49.0405 2.53 49.0805 2.93 ;
      RECT MASK 1 47.0405 2.538 47.0805 2.922 ;
      RECT MASK 1 47.6405 2.538 47.6805 2.922 ;
      RECT MASK 1 4.0065 2.575 4.0665 3.212 ;
      RECT MASK 1 42.8705 2.575 42.9305 3.212 ;
      RECT MASK 1 9.0445 2.631 9.1045 2.811 ;
      RECT MASK 1 9.5025 2.631 9.5625 2.811 ;
      RECT MASK 1 37.3745 2.631 37.4345 2.811 ;
      RECT MASK 1 37.8325 2.631 37.8925 2.811 ;
      RECT MASK 1 14.917 2.69 14.977 2.87 ;
      RECT MASK 1 15.375 2.69 15.435 2.87 ;
      RECT MASK 1 15.833 2.69 15.893 2.87 ;
      RECT MASK 1 16.291 2.69 16.351 2.87 ;
      RECT MASK 1 16.749 2.69 16.809 2.87 ;
      RECT MASK 1 17.665 2.69 17.725 2.87 ;
      RECT MASK 1 18.123 2.69 18.183 2.87 ;
      RECT MASK 1 19.039 2.69 19.099 2.87 ;
      RECT MASK 1 19.497 2.69 19.557 2.87 ;
      RECT MASK 1 19.955 2.69 20.015 2.87 ;
      RECT MASK 1 20.413 2.69 20.473 2.87 ;
      RECT MASK 1 20.871 2.69 20.931 2.87 ;
      RECT MASK 1 21.329 2.69 21.389 2.87 ;
      RECT MASK 1 25.548 2.69 25.608 2.87 ;
      RECT MASK 1 26.006 2.69 26.066 2.87 ;
      RECT MASK 1 26.464 2.69 26.524 2.87 ;
      RECT MASK 1 26.922 2.69 26.982 2.87 ;
      RECT MASK 1 27.38 2.69 27.44 2.87 ;
      RECT MASK 1 27.838 2.69 27.898 2.87 ;
      RECT MASK 1 28.754 2.69 28.814 2.87 ;
      RECT MASK 1 29.212 2.69 29.272 2.87 ;
      RECT MASK 1 30.128 2.69 30.188 2.87 ;
      RECT MASK 1 30.586 2.69 30.646 2.87 ;
      RECT MASK 1 31.044 2.69 31.104 2.87 ;
      RECT MASK 1 31.502 2.69 31.562 2.87 ;
      RECT MASK 1 31.96 2.69 32.02 2.87 ;
      RECT MASK 1 63.803 2.725 63.863 2.938 ;
      RECT MASK 1 64.261 2.725 64.321 2.938 ;
      RECT MASK 1 64.719 2.725 64.779 2.938 ;
      RECT MASK 1 62.887 2.758 62.947 3.842 ;
      RECT MASK 1 63.345 2.758 63.405 3.842 ;
      RECT MASK 1 65.177 2.758 65.237 3.515 ;
      RECT MASK 1 22.3385 2.855 22.3985 3.54 ;
      RECT MASK 1 22.5385 2.855 22.5985 3.54 ;
      RECT MASK 1 22.7385 2.855 22.7985 3.54 ;
      RECT MASK 1 22.9385 2.855 22.9985 3.54 ;
      RECT MASK 1 23.1385 2.855 23.1985 3.54 ;
      RECT MASK 1 23.7385 2.855 23.7985 3.54 ;
      RECT MASK 1 23.9385 2.855 23.9985 3.54 ;
      RECT MASK 1 24.1385 2.855 24.1985 3.54 ;
      RECT MASK 1 24.3385 2.855 24.3985 3.54 ;
      RECT MASK 1 24.5385 2.855 24.5985 3.54 ;
      RECT MASK 1 10.1875 2.8975 10.2475 4.4915 ;
      RECT MASK 1 10.6305 2.8975 10.6905 4.4915 ;
      RECT MASK 1 47.0405 2.96 47.0805 3.22 ;
      RECT MASK 1 47.6405 2.96 47.6805 3.22 ;
      RECT MASK 1 3.3195 3.032 3.3795 4.348 ;
      RECT MASK 1 3.7775 3.032 3.8375 4.348 ;
      RECT MASK 1 4.2355 3.032 4.2955 4.348 ;
      RECT MASK 1 4.6935 3.032 4.7535 4.348 ;
      RECT MASK 1 5.1515 3.032 5.2115 4.348 ;
      RECT MASK 1 5.6095 3.032 5.6695 4.348 ;
      RECT MASK 1 6.5255 3.032 6.5855 4.348 ;
      RECT MASK 1 7.4415 3.032 7.5015 4.348 ;
      RECT MASK 1 8.3575 3.032 8.4175 4.348 ;
      RECT MASK 1 8.8155 3.032 8.8755 3.245 ;
      RECT MASK 1 9.0445 3.032 9.1045 4.348 ;
      RECT MASK 1 9.2735 3.032 9.3335 3.25 ;
      RECT MASK 1 9.5025 3.032 9.5625 4.348 ;
      RECT MASK 1 9.7315 3.032 9.7915 3.25 ;
      RECT MASK 1 14.5735 3.032 14.6335 4.348 ;
      RECT MASK 1 15.0315 3.032 15.0915 4.348 ;
      RECT MASK 1 15.4895 3.032 15.5495 4.348 ;
      RECT MASK 1 15.9475 3.032 16.0075 4.348 ;
      RECT MASK 1 16.4055 3.032 16.4655 4.348 ;
      RECT MASK 1 16.8635 3.032 16.9235 4.348 ;
      RECT MASK 1 17.3215 3.032 17.3815 4.348 ;
      RECT MASK 1 17.7795 3.032 17.8395 4.348 ;
      RECT MASK 1 18.2375 3.032 18.2975 4.348 ;
      RECT MASK 1 18.6955 3.032 18.7555 4.348 ;
      RECT MASK 1 19.1535 3.032 19.2135 4.348 ;
      RECT MASK 1 19.6115 3.032 19.6715 4.348 ;
      RECT MASK 1 20.0695 3.032 20.1295 4.348 ;
      RECT MASK 1 20.5275 3.032 20.5875 4.348 ;
      RECT MASK 1 20.9855 3.032 21.0455 4.348 ;
      RECT MASK 1 21.4435 3.032 21.5035 4.348 ;
      RECT MASK 1 25.4335 3.032 25.4935 4.348 ;
      RECT MASK 1 25.8915 3.032 25.9515 4.348 ;
      RECT MASK 1 26.3495 3.032 26.4095 4.348 ;
      RECT MASK 1 26.8075 3.032 26.8675 4.348 ;
      RECT MASK 1 27.2655 3.032 27.3255 4.348 ;
      RECT MASK 1 27.7235 3.032 27.7835 4.348 ;
      RECT MASK 1 28.1815 3.032 28.2415 4.348 ;
      RECT MASK 1 28.6395 3.032 28.6995 4.348 ;
      RECT MASK 1 29.0975 3.032 29.1575 4.348 ;
      RECT MASK 1 29.5555 3.032 29.6155 4.348 ;
      RECT MASK 1 30.0135 3.032 30.0735 4.348 ;
      RECT MASK 1 30.4715 3.032 30.5315 4.348 ;
      RECT MASK 1 30.9295 3.032 30.9895 4.348 ;
      RECT MASK 1 31.3875 3.032 31.4475 4.348 ;
      RECT MASK 1 31.8455 3.032 31.9055 4.348 ;
      RECT MASK 1 32.3035 3.032 32.3635 4.348 ;
      RECT MASK 1 37.1455 3.032 37.2055 3.25 ;
      RECT MASK 1 37.3745 3.032 37.4345 4.348 ;
      RECT MASK 1 37.6035 3.032 37.6635 3.25 ;
      RECT MASK 1 37.8325 3.032 37.8925 4.348 ;
      RECT MASK 1 38.0615 3.032 38.1215 3.245 ;
      RECT MASK 1 38.5195 3.032 38.5795 4.348 ;
      RECT MASK 1 39.4355 3.032 39.4955 4.353 ;
      RECT MASK 1 40.3515 3.032 40.4115 4.353 ;
      RECT MASK 1 41.2675 3.032 41.3275 4.353 ;
      RECT MASK 1 41.7255 3.032 41.7855 4.353 ;
      RECT MASK 1 42.1835 3.032 42.2435 4.353 ;
      RECT MASK 1 42.6415 3.032 42.7015 4.353 ;
      RECT MASK 1 43.0995 3.032 43.1595 4.353 ;
      RECT MASK 1 43.5575 3.032 43.6175 4.353 ;
      RECT MASK 1 43.7865 3.032 43.8465 4.353 ;
      RECT MASK 1 64.49 3.058 64.55 3.542 ;
      RECT MASK 1 41.4965 3.1325 41.5565 4.2315 ;
      RECT MASK 1 59.5665 3.159 59.6265 3.441 ;
      RECT MASK 1 63.574 3.205 63.634 3.542 ;
      RECT MASK 1 46.8405 3.25 46.8805 3.65 ;
      RECT MASK 1 47.2405 3.25 47.2805 3.65 ;
      RECT MASK 1 47.4405 3.25 47.4805 3.65 ;
      RECT MASK 1 47.8405 3.25 47.8805 3.65 ;
      RECT MASK 1 48.0405 3.25 48.0805 3.65 ;
      RECT MASK 1 48.2405 3.25 48.2805 3.65 ;
      RECT MASK 1 48.4405 3.25 48.4805 3.77 ;
      RECT MASK 1 48.6405 3.25 48.6805 3.65 ;
      RECT MASK 1 48.8405 3.25 48.8805 3.65 ;
      RECT MASK 1 49.0405 3.25 49.0805 3.65 ;
      RECT MASK 1 47.0405 3.258 47.0805 3.642 ;
      RECT MASK 1 47.6405 3.258 47.6805 3.642 ;
      RECT MASK 1 3.0905 3.294 3.1505 4.086 ;
      RECT MASK 1 5.3805 3.294 5.4405 4.086 ;
      RECT MASK 1 8.5865 3.294 8.6465 4.086 ;
      RECT MASK 1 9.9605 3.294 10.0205 4.086 ;
      RECT MASK 1 36.9165 3.294 36.9765 4.086 ;
      RECT MASK 1 38.2905 3.294 38.3505 4.086 ;
      RECT MASK 1 63.8 3.3 63.86 3.487 ;
      RECT MASK 1 58.536 3.361 58.596 4.799 ;
      RECT MASK 1 60.368 3.361 60.428 4.799 ;
      RECT MASK 1 65.635 3.445 65.695 3.842 ;
      RECT MASK 1 61.971 3.5225 62.031 4.6375 ;
      RECT MASK 1 72.7295 3.527 72.8295 8.8515 ;
      RECT MASK 1 113.8755 3.527 113.9755 8.8515 ;
      RECT MASK 1 73.9545 3.54 74.2745 8.822 ;
      RECT MASK 1 75.4865 3.54 75.8065 8.822 ;
      RECT MASK 1 78.6125 3.54 78.9325 10.538 ;
      RECT MASK 1 80.9105 3.54 81.2305 10.538 ;
      RECT MASK 1 82.2575 3.54 82.3575 10.5615 ;
      RECT MASK 1 104.3475 3.54 104.4475 10.5615 ;
      RECT MASK 1 105.4745 3.54 105.7945 10.538 ;
      RECT MASK 1 107.7725 3.54 108.0925 10.538 ;
      RECT MASK 1 110.8985 3.54 111.2185 8.822 ;
      RECT MASK 1 112.4305 3.54 112.7505 8.822 ;
      RECT MASK 1 50.1875 3.545 50.2275 10.375 ;
      RECT MASK 1 50.4095 3.545 50.4495 8.095 ;
      RECT MASK 1 50.8515 3.545 50.8915 10.375 ;
      RECT MASK 1 51.0735 3.545 51.1135 8.095 ;
      RECT MASK 1 51.5155 3.545 51.5555 10.375 ;
      RECT MASK 1 51.7375 3.545 51.7775 8.095 ;
      RECT MASK 1 52.1795 3.545 52.2195 10.375 ;
      RECT MASK 1 52.4015 3.545 52.4415 8.095 ;
      RECT MASK 1 66.5645 3.563 66.6245 8.221 ;
      RECT MASK 1 58.994 3.662 59.054 4.498 ;
      RECT MASK 1 59.452 3.662 59.512 4.498 ;
      RECT MASK 1 59.91 3.662 59.97 4.498 ;
      RECT MASK 1 63.803 3.662 63.863 3.875 ;
      RECT MASK 1 64.261 3.662 64.321 3.875 ;
      RECT MASK 1 64.719 3.662 64.779 3.875 ;
      RECT MASK 1 65.177 3.662 65.237 3.875 ;
      RECT MASK 1 47.0405 3.68 47.0805 3.94 ;
      RECT MASK 1 47.6405 3.68 47.6805 3.94 ;
      RECT MASK 1 90.9345 3.78 91.0345 5.289 ;
      RECT MASK 1 91.9305 3.78 92.0305 6.54 ;
      RECT MASK 1 92.5945 3.78 92.6945 6.54 ;
      RECT MASK 1 92.9535 3.78 93.0535 6.54 ;
      RECT MASK 1 93.6515 3.78 93.7515 6.54 ;
      RECT MASK 1 94.0105 3.78 94.1105 6.54 ;
      RECT MASK 1 94.6745 3.78 94.7745 6.54 ;
      RECT MASK 1 95.6705 3.78 95.7705 5.289 ;
      RECT MASK 1 22.3385 3.84 22.3985 4.525 ;
      RECT MASK 1 22.5385 3.84 22.5985 4.525 ;
      RECT MASK 1 22.7385 3.84 22.7985 4.525 ;
      RECT MASK 1 22.9385 3.84 22.9985 4.525 ;
      RECT MASK 1 23.1385 3.84 23.1985 4.525 ;
      RECT MASK 1 23.7385 3.84 23.7985 4.525 ;
      RECT MASK 1 23.9385 3.84 23.9985 4.525 ;
      RECT MASK 1 24.1385 3.84 24.1985 4.525 ;
      RECT MASK 1 24.3385 3.84 24.3985 4.525 ;
      RECT MASK 1 24.5385 3.84 24.5985 4.525 ;
      RECT MASK 1 48.6405 3.85 48.6805 4.225 ;
      RECT MASK 1 46.8405 3.97 46.8805 4.225 ;
      RECT MASK 1 47.2405 3.97 47.2805 4.225 ;
      RECT MASK 1 47.4405 3.97 47.4805 4.225 ;
      RECT MASK 1 47.8405 3.97 47.8805 4.225 ;
      RECT MASK 1 48.0405 3.97 48.0805 4.225 ;
      RECT MASK 1 48.2405 3.97 48.2805 4.225 ;
      RECT MASK 1 48.4405 3.97 48.4805 4.225 ;
      RECT MASK 1 48.8405 3.97 48.8805 4.225 ;
      RECT MASK 1 49.0405 3.97 49.0805 4.225 ;
      RECT MASK 1 47.0405 3.978 47.0805 4.225 ;
      RECT MASK 1 47.6405 3.978 47.6805 4.225 ;
      RECT MASK 1 9.2735 4.13 9.3335 4.348 ;
      RECT MASK 1 9.7315 4.13 9.7915 4.348 ;
      RECT MASK 1 37.1455 4.13 37.2055 4.348 ;
      RECT MASK 1 37.6035 4.13 37.6635 4.348 ;
      RECT MASK 1 8.8155 4.135 8.8755 4.348 ;
      RECT MASK 1 38.0615 4.135 38.1215 4.348 ;
      RECT MASK 1 80.1445 4.159 80.4645 5.015 ;
      RECT MASK 1 106.2405 4.159 106.5605 5.015 ;
      RECT MASK 1 74.7205 4.162 75.0405 5.36 ;
      RECT MASK 1 79.3785 4.162 79.6985 7.535 ;
      RECT MASK 1 107.0065 4.162 107.3265 7.535 ;
      RECT MASK 1 111.6645 4.162 111.9845 5.36 ;
      RECT MASK 1 2.4035 4.168 2.4635 5.252 ;
      RECT MASK 1 2.8615 4.168 2.9215 5.252 ;
      RECT MASK 1 3.5485 4.168 3.6085 5.252 ;
      RECT MASK 1 4.0065 4.168 4.0665 4.805 ;
      RECT MASK 1 4.4645 4.168 4.5245 5.252 ;
      RECT MASK 1 4.9225 4.168 4.9825 5.252 ;
      RECT MASK 1 6.0675 4.168 6.1275 5.252 ;
      RECT MASK 1 6.9835 4.168 7.0435 5.252 ;
      RECT MASK 1 7.8995 4.168 7.9595 5.252 ;
      RECT MASK 1 11.3455 4.168 11.4055 5.252 ;
      RECT MASK 1 11.8035 4.168 11.8635 5.252 ;
      RECT MASK 1 12.2615 4.168 12.3215 5.252 ;
      RECT MASK 1 12.7195 4.168 12.7795 5.252 ;
      RECT MASK 1 34.1575 4.168 34.2175 5.252 ;
      RECT MASK 1 34.6155 4.168 34.6755 5.252 ;
      RECT MASK 1 35.0735 4.168 35.1335 5.252 ;
      RECT MASK 1 35.5315 4.168 35.5915 5.252 ;
      RECT MASK 1 38.9775 4.168 39.0375 5.252 ;
      RECT MASK 1 39.8935 4.168 39.9535 5.252 ;
      RECT MASK 1 40.8095 4.168 40.8695 5.252 ;
      RECT MASK 1 41.9545 4.168 42.0145 5.252 ;
      RECT MASK 1 42.4125 4.168 42.4725 5.252 ;
      RECT MASK 1 42.8705 4.168 42.9305 4.805 ;
      RECT MASK 1 43.3285 4.168 43.3885 5.252 ;
      RECT MASK 1 44.0155 4.168 44.0755 5.252 ;
      RECT MASK 1 44.4735 4.168 44.5335 5.252 ;
      RECT MASK 1 63.803 4.285 63.863 4.498 ;
      RECT MASK 1 64.261 4.285 64.321 4.498 ;
      RECT MASK 1 64.719 4.285 64.779 4.498 ;
      RECT MASK 1 65.177 4.285 65.237 4.498 ;
      RECT MASK 1 62.887 4.318 62.947 5.402 ;
      RECT MASK 1 63.345 4.318 63.405 5.402 ;
      RECT MASK 1 65.635 4.318 65.695 4.715 ;
      RECT MASK 1 10.8455 4.37 10.9055 5.045 ;
      RECT MASK 1 36.0315 4.37 36.0915 5.045 ;
      RECT MASK 1 8.5865 4.375 8.6465 5.045 ;
      RECT MASK 1 38.2905 4.375 38.3505 5.045 ;
      RECT MASK 1 5.3805 4.468 5.4405 5.05 ;
      RECT MASK 1 6.2965 4.468 6.3565 5.285 ;
      RECT MASK 1 7.2125 4.468 7.2725 4.952 ;
      RECT MASK 1 39.6645 4.468 39.7245 4.952 ;
      RECT MASK 1 40.5805 4.468 40.6405 5.285 ;
      RECT MASK 1 41.4965 4.468 41.5565 5.05 ;
      RECT MASK 1 61.055 4.4825 61.115 5.725 ;
      RECT MASK 1 84.6265 4.488 84.7265 5.168 ;
      RECT MASK 1 85.6225 4.488 85.7225 5.168 ;
      RECT MASK 1 86.6185 4.488 86.7185 5.168 ;
      RECT MASK 1 87.6145 4.488 87.7145 5.168 ;
      RECT MASK 1 89.2745 4.488 89.3745 5.168 ;
      RECT MASK 1 90.2705 4.488 90.3705 5.168 ;
      RECT MASK 1 91.2665 4.488 91.3665 5.168 ;
      RECT MASK 1 95.3385 4.488 95.4385 5.168 ;
      RECT MASK 1 96.3345 4.488 96.4345 5.168 ;
      RECT MASK 1 97.3305 4.488 97.4305 5.168 ;
      RECT MASK 1 98.9905 4.488 99.0905 5.168 ;
      RECT MASK 1 99.9865 4.488 100.0865 5.168 ;
      RECT MASK 1 100.9825 4.488 101.0825 5.168 ;
      RECT MASK 1 101.9785 4.488 102.0785 5.168 ;
      RECT MASK 1 14.917 4.51 14.977 4.69 ;
      RECT MASK 1 15.375 4.51 15.435 4.69 ;
      RECT MASK 1 15.833 4.51 15.893 4.69 ;
      RECT MASK 1 16.291 4.51 16.351 4.69 ;
      RECT MASK 1 16.749 4.51 16.809 4.69 ;
      RECT MASK 1 17.665 4.51 17.725 4.69 ;
      RECT MASK 1 18.123 4.51 18.183 4.69 ;
      RECT MASK 1 19.039 4.51 19.099 4.69 ;
      RECT MASK 1 19.497 4.51 19.557 4.69 ;
      RECT MASK 1 19.955 4.51 20.015 4.69 ;
      RECT MASK 1 20.413 4.51 20.473 4.69 ;
      RECT MASK 1 20.871 4.51 20.931 4.69 ;
      RECT MASK 1 21.329 4.51 21.389 4.69 ;
      RECT MASK 1 25.548 4.51 25.608 4.69 ;
      RECT MASK 1 26.006 4.51 26.066 4.69 ;
      RECT MASK 1 26.464 4.51 26.524 4.69 ;
      RECT MASK 1 26.922 4.51 26.982 4.69 ;
      RECT MASK 1 27.38 4.51 27.44 4.69 ;
      RECT MASK 1 27.838 4.51 27.898 4.69 ;
      RECT MASK 1 28.754 4.51 28.814 4.69 ;
      RECT MASK 1 29.212 4.51 29.272 4.69 ;
      RECT MASK 1 30.128 4.51 30.188 4.69 ;
      RECT MASK 1 30.586 4.51 30.646 4.69 ;
      RECT MASK 1 31.044 4.51 31.104 4.69 ;
      RECT MASK 1 31.502 4.51 31.562 4.69 ;
      RECT MASK 1 31.96 4.51 32.02 4.69 ;
      RECT MASK 1 56.592 4.523 56.652 6.472 ;
      RECT MASK 1 66.882 4.523 66.942 5.6575 ;
      RECT MASK 1 87.2825 4.557 87.3825 5.9975 ;
      RECT MASK 1 99.3225 4.557 99.4225 5.9975 ;
      RECT MASK 1 9.0445 4.569 9.1045 4.749 ;
      RECT MASK 1 9.5025 4.569 9.5625 4.749 ;
      RECT MASK 1 37.3745 4.569 37.4345 4.749 ;
      RECT MASK 1 37.8325 4.569 37.8925 4.749 ;
      RECT MASK 1 85.2905 4.609 85.3905 6.625 ;
      RECT MASK 1 86.2865 4.609 86.3865 5.345 ;
      RECT MASK 1 88.9425 4.609 89.0425 5.289 ;
      RECT MASK 1 89.9385 4.609 90.0385 5.289 ;
      RECT MASK 1 96.6665 4.609 96.7665 5.289 ;
      RECT MASK 1 97.6625 4.609 97.7625 5.289 ;
      RECT MASK 1 100.3185 4.609 100.4185 5.345 ;
      RECT MASK 1 101.3145 4.609 101.4145 6.625 ;
      RECT MASK 1 11.0955 4.61 11.1555 4.851 ;
      RECT MASK 1 35.7815 4.61 35.8415 4.851 ;
      RECT MASK 1 9.9815 4.615 10.0415 4.851 ;
      RECT MASK 1 36.8955 4.615 36.9555 4.851 ;
      RECT MASK 1 63.574 4.618 63.634 4.955 ;
      RECT MASK 1 64.49 4.618 64.55 5.102 ;
      RECT MASK 1 65.177 4.645 65.237 5.402 ;
      RECT MASK 1 63.8 4.673 63.86 4.86 ;
      RECT MASK 1 23.7385 4.6795 23.7985 4.911 ;
      RECT MASK 1 22.9385 4.68 22.9985 4.82 ;
      RECT MASK 1 59.5665 4.719 59.6265 5.001 ;
      RECT MASK 1 88.3185 4.7235 88.3785 6.54 ;
      RECT MASK 1 98.3265 4.7235 98.3865 6.54 ;
      RECT MASK 1 8.8155 4.73 8.8755 5.252 ;
      RECT MASK 1 9.2735 4.73 9.3335 5.252 ;
      RECT MASK 1 12.9915 4.73 13.0515 4.91 ;
      RECT MASK 1 14.688 4.73 14.748 4.91 ;
      RECT MASK 1 15.146 4.73 15.206 4.91 ;
      RECT MASK 1 15.604 4.73 15.664 4.91 ;
      RECT MASK 1 16.062 4.73 16.122 4.91 ;
      RECT MASK 1 16.52 4.73 16.58 4.91 ;
      RECT MASK 1 16.978 4.73 17.038 4.91 ;
      RECT MASK 1 17.436 4.73 17.496 4.91 ;
      RECT MASK 1 18.352 4.73 18.412 4.91 ;
      RECT MASK 1 18.81 4.73 18.87 4.91 ;
      RECT MASK 1 19.726 4.73 19.786 4.91 ;
      RECT MASK 1 20.642 4.73 20.702 4.91 ;
      RECT MASK 1 21.1 4.73 21.16 4.91 ;
      RECT MASK 1 25.777 4.73 25.837 4.91 ;
      RECT MASK 1 26.235 4.73 26.295 4.91 ;
      RECT MASK 1 27.151 4.73 27.211 4.91 ;
      RECT MASK 1 28.067 4.73 28.127 4.91 ;
      RECT MASK 1 28.525 4.73 28.585 4.91 ;
      RECT MASK 1 29.441 4.73 29.501 4.91 ;
      RECT MASK 1 29.899 4.73 29.959 4.91 ;
      RECT MASK 1 30.357 4.73 30.417 4.91 ;
      RECT MASK 1 30.815 4.73 30.875 4.91 ;
      RECT MASK 1 31.273 4.73 31.333 4.91 ;
      RECT MASK 1 31.731 4.73 31.791 4.91 ;
      RECT MASK 1 32.189 4.73 32.249 4.91 ;
      RECT MASK 1 33.8855 4.73 33.9455 4.91 ;
      RECT MASK 1 37.6035 4.73 37.6635 5.252 ;
      RECT MASK 1 38.0615 4.73 38.1215 5.252 ;
      RECT MASK 1 84.9585 4.73 85.0585 5.41 ;
      RECT MASK 1 85.9545 4.73 86.0545 5.41 ;
      RECT MASK 1 86.9505 4.73 87.0505 5.41 ;
      RECT MASK 1 87.9465 4.73 88.0465 5.41 ;
      RECT MASK 1 89.6065 4.73 89.7065 5.41 ;
      RECT MASK 1 90.6025 4.73 90.7025 5.41 ;
      RECT MASK 1 91.5985 4.73 91.6985 5.4165 ;
      RECT MASK 1 95.0065 4.73 95.1065 5.4165 ;
      RECT MASK 1 96.0025 4.73 96.1025 5.41 ;
      RECT MASK 1 96.9985 4.73 97.0985 5.41 ;
      RECT MASK 1 98.6585 4.73 98.7585 5.41 ;
      RECT MASK 1 99.6545 4.73 99.7545 5.41 ;
      RECT MASK 1 100.6505 4.73 100.7505 5.41 ;
      RECT MASK 1 101.6465 4.73 101.7465 5.41 ;
      RECT MASK 1 9.7315 4.735 9.7915 5.252 ;
      RECT MASK 1 37.1455 4.735 37.2055 5.252 ;
      RECT MASK 1 57.053 4.762 57.113 5.371 ;
      RECT MASK 1 22.5385 4.94 22.5985 5.565 ;
      RECT MASK 1 22.7385 4.94 22.7985 5.565 ;
      RECT MASK 1 22.9385 4.94 22.9985 5.565 ;
      RECT MASK 1 23.9385 4.94 23.9985 5.565 ;
      RECT MASK 1 24.1385 4.94 24.1985 5.565 ;
      RECT MASK 1 24.3385 4.94 24.3985 5.565 ;
      RECT MASK 1 4.0065 4.975 4.0665 5.252 ;
      RECT MASK 1 9.0445 4.975 9.1045 5.252 ;
      RECT MASK 1 37.8325 4.975 37.8925 5.252 ;
      RECT MASK 1 42.8705 4.975 42.9305 5.252 ;
      RECT MASK 1 65.635 5.022 65.695 6.0775 ;
      RECT MASK 1 22.3385 5.031 22.3985 5.565 ;
      RECT MASK 1 23.1385 5.031 23.1985 5.565 ;
      RECT MASK 1 23.7385 5.031 23.7985 5.565 ;
      RECT MASK 1 24.5385 5.031 24.5985 5.565 ;
      RECT MASK 1 5.1515 5.071 5.2115 6.389 ;
      RECT MASK 1 41.7255 5.071 41.7855 6.389 ;
      RECT MASK 1 3.3195 5.072 3.3795 6.388 ;
      RECT MASK 1 3.7775 5.072 3.8375 6.388 ;
      RECT MASK 1 4.2355 5.072 4.2955 6.388 ;
      RECT MASK 1 4.6935 5.072 4.7535 6.388 ;
      RECT MASK 1 5.6095 5.072 5.6695 6.388 ;
      RECT MASK 1 6.5255 5.072 6.5855 6.388 ;
      RECT MASK 1 7.4415 5.072 7.5015 6.388 ;
      RECT MASK 1 9.5025 5.072 9.5625 5.29 ;
      RECT MASK 1 14.5735 5.072 14.6335 6.388 ;
      RECT MASK 1 15.0315 5.072 15.0915 6.388 ;
      RECT MASK 1 15.4895 5.072 15.5495 6.388 ;
      RECT MASK 1 15.9475 5.072 16.0075 6.388 ;
      RECT MASK 1 16.4055 5.072 16.4655 6.388 ;
      RECT MASK 1 16.8635 5.072 16.9235 6.388 ;
      RECT MASK 1 17.3215 5.072 17.3815 6.388 ;
      RECT MASK 1 17.7795 5.072 17.8395 6.388 ;
      RECT MASK 1 18.2375 5.072 18.2975 6.388 ;
      RECT MASK 1 18.6955 5.072 18.7555 6.388 ;
      RECT MASK 1 19.1535 5.072 19.2135 6.388 ;
      RECT MASK 1 19.6115 5.072 19.6715 6.388 ;
      RECT MASK 1 20.0695 5.072 20.1295 6.388 ;
      RECT MASK 1 20.5275 5.072 20.5875 6.388 ;
      RECT MASK 1 20.9855 5.072 21.0455 6.388 ;
      RECT MASK 1 21.4435 5.072 21.5035 6.388 ;
      RECT MASK 1 25.4335 5.072 25.4935 6.388 ;
      RECT MASK 1 25.8915 5.072 25.9515 6.388 ;
      RECT MASK 1 26.3495 5.072 26.4095 6.388 ;
      RECT MASK 1 26.8075 5.072 26.8675 6.388 ;
      RECT MASK 1 27.2655 5.072 27.3255 6.388 ;
      RECT MASK 1 27.7235 5.072 27.7835 6.388 ;
      RECT MASK 1 28.1815 5.072 28.2415 6.388 ;
      RECT MASK 1 28.6395 5.072 28.6995 6.388 ;
      RECT MASK 1 29.0975 5.072 29.1575 6.388 ;
      RECT MASK 1 29.5555 5.072 29.6155 6.388 ;
      RECT MASK 1 30.0135 5.072 30.0735 6.388 ;
      RECT MASK 1 30.4715 5.072 30.5315 6.388 ;
      RECT MASK 1 30.9295 5.072 30.9895 6.388 ;
      RECT MASK 1 31.3875 5.072 31.4475 6.388 ;
      RECT MASK 1 31.8455 5.072 31.9055 6.388 ;
      RECT MASK 1 32.3035 5.072 32.3635 6.388 ;
      RECT MASK 1 37.3745 5.072 37.4345 5.29 ;
      RECT MASK 1 39.4355 5.072 39.4955 6.388 ;
      RECT MASK 1 40.3515 5.072 40.4115 6.388 ;
      RECT MASK 1 41.2675 5.072 41.3275 6.388 ;
      RECT MASK 1 42.1835 5.072 42.2435 6.388 ;
      RECT MASK 1 42.6415 5.072 42.7015 6.388 ;
      RECT MASK 1 43.0995 5.072 43.1595 6.388 ;
      RECT MASK 1 43.5575 5.072 43.6175 6.388 ;
      RECT MASK 1 8.3575 5.0725 8.4175 6.3875 ;
      RECT MASK 1 38.5195 5.0725 38.5795 6.3875 ;
      RECT MASK 1 46.7995 5.135 46.8595 5.781 ;
      RECT MASK 1 47.1315 5.135 47.1915 5.786 ;
      RECT MASK 1 47.4635 5.135 47.5235 5.786 ;
      RECT MASK 1 47.7955 5.135 47.8555 5.781 ;
      RECT MASK 1 48.1275 5.135 48.1875 5.786 ;
      RECT MASK 1 48.4595 5.135 48.5195 5.781 ;
      RECT MASK 1 48.8745 5.135 48.9345 6.0475 ;
      RECT MASK 1 61.971 5.2025 62.031 5.73 ;
      RECT MASK 1 58.536 5.222 58.596 5.722 ;
      RECT MASK 1 58.994 5.222 59.054 5.722 ;
      RECT MASK 1 59.452 5.222 59.512 5.722 ;
      RECT MASK 1 59.91 5.222 59.97 5.722 ;
      RECT MASK 1 60.368 5.222 60.428 5.722 ;
      RECT MASK 1 63.803 5.222 63.863 5.435 ;
      RECT MASK 1 64.261 5.222 64.321 5.435 ;
      RECT MASK 1 64.719 5.222 64.779 5.435 ;
      RECT MASK 1 53.9295 5.255 53.9895 6.1675 ;
      RECT MASK 1 54.3445 5.255 54.4045 5.901 ;
      RECT MASK 1 54.6765 5.255 54.7365 5.906 ;
      RECT MASK 1 54.8425 5.255 54.9025 5.726 ;
      RECT MASK 1 55.1745 5.255 55.2345 5.901 ;
      RECT MASK 1 55.3405 5.255 55.4005 5.726 ;
      RECT MASK 1 55.5065 5.255 55.5665 5.906 ;
      RECT MASK 1 55.8385 5.255 55.8985 5.901 ;
      RECT MASK 1 56.0875 5.255 56.1475 6.1675 ;
      RECT MASK 1 49.3445 5.301 49.4045 7.3995 ;
      RECT MASK 1 3.0905 5.334 3.1505 6.126 ;
      RECT MASK 1 5.3805 5.334 5.4405 6.126 ;
      RECT MASK 1 8.5865 5.334 8.6465 6.126 ;
      RECT MASK 1 9.9605 5.334 10.0205 6.126 ;
      RECT MASK 1 36.9165 5.334 36.9765 6.126 ;
      RECT MASK 1 38.2905 5.334 38.3505 6.126 ;
      RECT MASK 1 41.4965 5.334 41.5565 6.126 ;
      RECT MASK 1 43.7865 5.334 43.8465 6.126 ;
      RECT MASK 1 58.765 5.558 58.825 6.058 ;
      RECT MASK 1 59.223 5.558 59.283 6.058 ;
      RECT MASK 1 59.681 5.558 59.741 6.058 ;
      RECT MASK 1 63.803 5.558 63.863 6.058 ;
      RECT MASK 1 64.261 5.558 64.321 6.058 ;
      RECT MASK 1 64.719 5.558 64.779 6.058 ;
      RECT MASK 1 87.6145 5.6585 87.7145 7.6 ;
      RECT MASK 1 98.9905 5.6585 99.0905 7.6 ;
      RECT MASK 1 89.0145 5.673 89.0745 6.54 ;
      RECT MASK 1 89.8305 5.673 89.8905 6.54 ;
      RECT MASK 1 90.0825 5.673 90.1425 6.54 ;
      RECT MASK 1 90.5745 5.673 90.6345 6.54 ;
      RECT MASK 1 96.0705 5.673 96.1305 6.54 ;
      RECT MASK 1 96.5625 5.673 96.6225 6.54 ;
      RECT MASK 1 96.8145 5.673 96.8745 6.54 ;
      RECT MASK 1 97.6305 5.673 97.6905 6.54 ;
      RECT MASK 1 86.9545 5.68 87.0545 6.54 ;
      RECT MASK 1 99.6505 5.68 99.7505 6.54 ;
      RECT MASK 1 89.5785 5.7275 89.6385 7.721 ;
      RECT MASK 1 97.0665 5.7275 97.1265 7.721 ;
      RECT MASK 1 88.5705 5.7995 88.6305 7.721 ;
      RECT MASK 1 98.0745 5.7995 98.1345 7.721 ;
      RECT MASK 1 90.3335 5.809 90.3935 7.721 ;
      RECT MASK 1 96.3115 5.809 96.3715 7.721 ;
      RECT MASK 1 60.826 5.845 60.886 7 ;
      RECT MASK 1 61.284 5.845 61.344 6.058 ;
      RECT MASK 1 61.742 5.845 61.802 6.058 ;
      RECT MASK 1 62.2 5.845 62.26 6.058 ;
      RECT MASK 1 62.658 5.845 62.718 6.058 ;
      RECT MASK 1 63.116 5.845 63.176 7 ;
      RECT MASK 1 86.6185 5.846 86.7185 7.6 ;
      RECT MASK 1 99.9865 5.846 100.0865 7.6 ;
      RECT MASK 1 90.834 5.8565 90.894 7.6 ;
      RECT MASK 1 95.811 5.8565 95.871 7.6 ;
      RECT MASK 1 22.3385 5.895 22.3985 6.429 ;
      RECT MASK 1 22.5385 5.895 22.5985 6.52 ;
      RECT MASK 1 22.7385 5.895 22.7985 6.52 ;
      RECT MASK 1 22.9385 5.895 22.9985 6.52 ;
      RECT MASK 1 23.1385 5.895 23.1985 6.429 ;
      RECT MASK 1 23.7385 5.895 23.7985 6.429 ;
      RECT MASK 1 23.9385 5.895 23.9985 6.52 ;
      RECT MASK 1 24.1385 5.895 24.1985 6.52 ;
      RECT MASK 1 24.3385 5.895 24.3985 6.52 ;
      RECT MASK 1 24.5385 5.895 24.5985 6.429 ;
      RECT MASK 1 47.1315 5.906 47.1915 6.514 ;
      RECT MASK 1 47.4635 5.906 47.5235 6.514 ;
      RECT MASK 1 88.7735 5.909 88.8335 7.6 ;
      RECT MASK 1 89.2555 5.909 89.3155 7.6 ;
      RECT MASK 1 97.3895 5.909 97.4495 7.6 ;
      RECT MASK 1 97.8715 5.909 97.9315 7.6 ;
      RECT MASK 1 54.8425 5.918 54.9025 6.742 ;
      RECT MASK 1 60.2275 5.9225 60.2875 8.4775 ;
      RECT MASK 1 84.6265 5.93 84.7265 7.6 ;
      RECT MASK 1 101.9785 5.93 102.0785 7.6 ;
      RECT MASK 1 55.1745 6.021 55.2345 6.639 ;
      RECT MASK 1 54.6765 6.026 54.7365 6.634 ;
      RECT MASK 1 55.5065 6.026 55.5665 6.634 ;
      RECT MASK 1 9.5025 6.17 9.5625 6.388 ;
      RECT MASK 1 37.3745 6.17 37.4345 6.388 ;
      RECT MASK 1 6.2965 6.175 6.3565 6.992 ;
      RECT MASK 1 40.5805 6.175 40.6405 6.992 ;
      RECT MASK 1 62.2 6.178 62.26 6.561 ;
      RECT MASK 1 62.658 6.178 62.718 6.561 ;
      RECT MASK 1 2.4035 6.208 2.4635 7.292 ;
      RECT MASK 1 2.8615 6.208 2.9215 7.292 ;
      RECT MASK 1 3.5485 6.208 3.6085 7.292 ;
      RECT MASK 1 4.0065 6.208 4.0665 6.485 ;
      RECT MASK 1 4.4645 6.208 4.5245 7.292 ;
      RECT MASK 1 4.9225 6.208 4.9825 7.292 ;
      RECT MASK 1 6.0675 6.208 6.1275 7.292 ;
      RECT MASK 1 6.9835 6.208 7.0435 7.292 ;
      RECT MASK 1 7.8995 6.208 7.9595 7.292 ;
      RECT MASK 1 8.8155 6.208 8.8755 6.73 ;
      RECT MASK 1 9.0445 6.208 9.1045 6.485 ;
      RECT MASK 1 9.2735 6.208 9.3335 6.73 ;
      RECT MASK 1 9.7315 6.208 9.7915 6.725 ;
      RECT MASK 1 11.3455 6.208 11.4055 7.292 ;
      RECT MASK 1 11.8035 6.208 11.8635 7.292 ;
      RECT MASK 1 12.2615 6.208 12.3215 7.292 ;
      RECT MASK 1 12.7195 6.208 12.7795 7.292 ;
      RECT MASK 1 34.1575 6.208 34.2175 7.292 ;
      RECT MASK 1 34.6155 6.208 34.6755 7.292 ;
      RECT MASK 1 35.0735 6.208 35.1335 7.292 ;
      RECT MASK 1 35.5315 6.208 35.5915 7.292 ;
      RECT MASK 1 37.1455 6.208 37.2055 6.725 ;
      RECT MASK 1 37.6035 6.208 37.6635 6.73 ;
      RECT MASK 1 37.8325 6.208 37.8925 6.485 ;
      RECT MASK 1 38.0615 6.208 38.1215 6.73 ;
      RECT MASK 1 38.9775 6.208 39.0375 7.292 ;
      RECT MASK 1 39.8935 6.208 39.9535 7.292 ;
      RECT MASK 1 40.8095 6.208 40.8695 7.292 ;
      RECT MASK 1 41.9545 6.208 42.0145 7.292 ;
      RECT MASK 1 42.4125 6.208 42.4725 7.292 ;
      RECT MASK 1 42.8705 6.208 42.9305 6.485 ;
      RECT MASK 1 43.3285 6.208 43.3885 7.292 ;
      RECT MASK 1 44.0155 6.208 44.0755 7.292 ;
      RECT MASK 1 44.4735 6.208 44.5335 7.292 ;
      RECT MASK 1 58.765 6.279 58.825 6.561 ;
      RECT MASK 1 59.223 6.279 59.283 6.561 ;
      RECT MASK 1 59.681 6.279 59.741 6.561 ;
      RECT MASK 1 61.284 6.279 61.344 6.662 ;
      RECT MASK 1 61.742 6.279 61.802 6.662 ;
      RECT MASK 1 63.803 6.279 63.863 6.561 ;
      RECT MASK 1 64.261 6.279 64.321 6.561 ;
      RECT MASK 1 64.719 6.279 64.779 6.561 ;
      RECT MASK 1 53.079 6.301 53.139 9.185 ;
      RECT MASK 1 5.3805 6.41 5.4405 6.992 ;
      RECT MASK 1 41.4965 6.41 41.5565 6.992 ;
      RECT MASK 1 8.5865 6.415 8.6465 7.085 ;
      RECT MASK 1 10.8455 6.415 10.9055 7.09 ;
      RECT MASK 1 36.0315 6.415 36.0915 7.09 ;
      RECT MASK 1 38.2905 6.415 38.3505 7.085 ;
      RECT MASK 1 7.2125 6.508 7.2725 6.992 ;
      RECT MASK 1 39.6645 6.508 39.7245 6.992 ;
      RECT MASK 1 23.3385 6.535 23.3985 6.9215 ;
      RECT MASK 1 12.9915 6.55 13.0515 6.73 ;
      RECT MASK 1 14.688 6.55 14.748 6.73 ;
      RECT MASK 1 15.146 6.55 15.206 6.73 ;
      RECT MASK 1 15.604 6.55 15.664 6.73 ;
      RECT MASK 1 16.062 6.55 16.122 6.73 ;
      RECT MASK 1 16.52 6.55 16.58 6.73 ;
      RECT MASK 1 16.978 6.55 17.038 6.73 ;
      RECT MASK 1 17.436 6.55 17.496 6.73 ;
      RECT MASK 1 18.352 6.55 18.412 6.73 ;
      RECT MASK 1 18.81 6.55 18.87 6.73 ;
      RECT MASK 1 19.726 6.55 19.786 6.73 ;
      RECT MASK 1 20.642 6.55 20.702 6.73 ;
      RECT MASK 1 21.1 6.55 21.16 6.73 ;
      RECT MASK 1 25.777 6.55 25.837 6.73 ;
      RECT MASK 1 26.235 6.55 26.295 6.73 ;
      RECT MASK 1 27.151 6.55 27.211 6.73 ;
      RECT MASK 1 28.067 6.55 28.127 6.73 ;
      RECT MASK 1 28.525 6.55 28.585 6.73 ;
      RECT MASK 1 29.441 6.55 29.501 6.73 ;
      RECT MASK 1 29.899 6.55 29.959 6.73 ;
      RECT MASK 1 30.357 6.55 30.417 6.73 ;
      RECT MASK 1 30.815 6.55 30.875 6.73 ;
      RECT MASK 1 31.273 6.55 31.333 6.73 ;
      RECT MASK 1 31.731 6.55 31.791 6.73 ;
      RECT MASK 1 32.189 6.55 32.249 6.73 ;
      RECT MASK 1 33.8855 6.55 33.9455 6.73 ;
      RECT MASK 1 23.7385 6.554 23.7985 6.78 ;
      RECT MASK 1 9.9815 6.609 10.0415 6.845 ;
      RECT MASK 1 11.0955 6.609 11.1555 6.85 ;
      RECT MASK 1 35.7815 6.609 35.8415 6.85 ;
      RECT MASK 1 36.8955 6.609 36.9555 6.845 ;
      RECT MASK 1 47.1315 6.634 47.1915 7.226 ;
      RECT MASK 1 47.4635 6.634 47.5235 7.226 ;
      RECT MASK 1 48.4595 6.634 48.5195 7.221 ;
      RECT MASK 1 46.7995 6.639 46.8595 7.221 ;
      RECT MASK 1 47.7955 6.639 47.8555 7.226 ;
      RECT MASK 1 48.2935 6.639 48.3535 7.221 ;
      RECT MASK 1 48.6255 6.639 48.6855 7.221 ;
      RECT MASK 1 65.635 6.6425 65.695 7.7575 ;
      RECT MASK 1 65.864 6.6425 65.924 7.7575 ;
      RECT MASK 1 4.0065 6.655 4.0665 7.292 ;
      RECT MASK 1 42.8705 6.655 42.9305 7.292 ;
      RECT MASK 1 9.0445 6.711 9.1045 6.891 ;
      RECT MASK 1 9.5025 6.711 9.5625 6.891 ;
      RECT MASK 1 37.3745 6.711 37.4345 6.891 ;
      RECT MASK 1 37.8325 6.711 37.8925 6.891 ;
      RECT MASK 1 49.9665 6.75 50.0065 9.122 ;
      RECT MASK 1 50.6305 6.75 50.6705 9.122 ;
      RECT MASK 1 51.2945 6.75 51.3345 9.122 ;
      RECT MASK 1 51.9585 6.75 51.9985 9.122 ;
      RECT MASK 1 52.6225 6.75 52.6625 9.122 ;
      RECT MASK 1 54.6765 6.754 54.7365 7.405 ;
      RECT MASK 1 55.5065 6.754 55.5665 7.405 ;
      RECT MASK 1 54.3445 6.759 54.4045 7.405 ;
      RECT MASK 1 55.1745 6.759 55.2345 7.405 ;
      RECT MASK 1 55.8385 6.759 55.8985 7.405 ;
      RECT MASK 1 14.917 6.77 14.977 6.95 ;
      RECT MASK 1 15.375 6.77 15.435 6.95 ;
      RECT MASK 1 15.833 6.77 15.893 6.95 ;
      RECT MASK 1 16.291 6.77 16.351 6.95 ;
      RECT MASK 1 16.749 6.77 16.809 6.95 ;
      RECT MASK 1 17.665 6.77 17.725 6.95 ;
      RECT MASK 1 18.123 6.77 18.183 6.95 ;
      RECT MASK 1 19.039 6.77 19.099 6.95 ;
      RECT MASK 1 19.497 6.77 19.557 6.95 ;
      RECT MASK 1 19.955 6.77 20.015 6.95 ;
      RECT MASK 1 20.413 6.77 20.473 6.95 ;
      RECT MASK 1 20.871 6.77 20.931 6.95 ;
      RECT MASK 1 21.329 6.77 21.389 6.95 ;
      RECT MASK 1 25.548 6.77 25.608 6.95 ;
      RECT MASK 1 26.006 6.77 26.066 6.95 ;
      RECT MASK 1 26.464 6.77 26.524 6.95 ;
      RECT MASK 1 26.922 6.77 26.982 6.95 ;
      RECT MASK 1 27.38 6.77 27.44 6.95 ;
      RECT MASK 1 27.838 6.77 27.898 6.95 ;
      RECT MASK 1 28.754 6.77 28.814 6.95 ;
      RECT MASK 1 29.212 6.77 29.272 6.95 ;
      RECT MASK 1 30.128 6.77 30.188 6.95 ;
      RECT MASK 1 30.586 6.77 30.646 6.95 ;
      RECT MASK 1 31.044 6.77 31.104 6.95 ;
      RECT MASK 1 31.502 6.77 31.562 6.95 ;
      RECT MASK 1 31.96 6.77 32.02 6.95 ;
      RECT MASK 1 58.765 6.782 58.825 7.618 ;
      RECT MASK 1 59.223 6.782 59.283 7.618 ;
      RECT MASK 1 59.681 6.782 59.741 7.618 ;
      RECT MASK 1 61.284 6.782 61.344 7 ;
      RECT MASK 1 61.742 6.782 61.802 7 ;
      RECT MASK 1 62.2 6.782 62.26 7 ;
      RECT MASK 1 62.658 6.782 62.718 7 ;
      RECT MASK 1 63.803 6.782 63.863 7.618 ;
      RECT MASK 1 64.261 6.782 64.321 7.618 ;
      RECT MASK 1 64.719 6.782 64.779 7.618 ;
      RECT MASK 1 47.9615 6.814 48.0215 7.046 ;
      RECT MASK 1 54.8425 6.934 54.9025 7.405 ;
      RECT MASK 1 55.3405 6.934 55.4005 7.405 ;
      RECT MASK 1 22.3385 6.935 22.3985 7.62 ;
      RECT MASK 1 22.5385 6.935 22.5985 7.62 ;
      RECT MASK 1 22.7385 6.935 22.7985 7.62 ;
      RECT MASK 1 22.9385 6.935 22.9985 7.62 ;
      RECT MASK 1 23.1385 6.935 23.1985 7.62 ;
      RECT MASK 1 23.7385 6.935 23.7985 7.62 ;
      RECT MASK 1 23.9385 6.935 23.9985 7.62 ;
      RECT MASK 1 24.1385 6.935 24.1985 7.62 ;
      RECT MASK 1 24.3385 6.935 24.3985 7.62 ;
      RECT MASK 1 24.5385 6.935 24.5985 7.62 ;
      RECT MASK 1 87.2825 6.96 87.3825 8.46 ;
      RECT MASK 1 99.3225 6.96 99.4225 8.46 ;
      RECT MASK 1 88.3185 6.965 88.3785 8.46 ;
      RECT MASK 1 89.0145 6.965 89.0745 8.46 ;
      RECT MASK 1 89.8305 6.965 89.8905 8.46 ;
      RECT MASK 1 90.0825 6.965 90.1425 8.46 ;
      RECT MASK 1 90.5865 6.965 90.6465 8.46 ;
      RECT MASK 1 91.0905 6.965 91.1505 8.46 ;
      RECT MASK 1 91.3425 6.965 91.4025 8.46 ;
      RECT MASK 1 95.3025 6.965 95.3625 8.46 ;
      RECT MASK 1 95.5545 6.965 95.6145 8.46 ;
      RECT MASK 1 96.0585 6.965 96.1185 8.46 ;
      RECT MASK 1 96.5625 6.965 96.6225 8.46 ;
      RECT MASK 1 96.8145 6.965 96.8745 8.46 ;
      RECT MASK 1 97.6305 6.965 97.6905 8.46 ;
      RECT MASK 1 98.3265 6.965 98.3865 8.46 ;
      RECT MASK 1 3.3195 7.112 3.3795 7.89 ;
      RECT MASK 1 3.7775 7.112 3.8375 7.89 ;
      RECT MASK 1 4.2355 7.112 4.2955 7.89 ;
      RECT MASK 1 4.6935 7.112 4.7535 7.89 ;
      RECT MASK 1 5.1515 7.112 5.2115 7.89 ;
      RECT MASK 1 5.6095 7.112 5.6695 7.89 ;
      RECT MASK 1 6.5255 7.112 6.5855 7.89 ;
      RECT MASK 1 7.4415 7.112 7.5015 7.89 ;
      RECT MASK 1 8.3575 7.112 8.4175 7.89 ;
      RECT MASK 1 8.8155 7.112 8.8755 7.325 ;
      RECT MASK 1 9.0445 7.112 9.1045 7.89 ;
      RECT MASK 1 9.2735 7.112 9.3335 7.33 ;
      RECT MASK 1 9.5025 7.112 9.5625 7.89 ;
      RECT MASK 1 9.7315 7.112 9.7915 7.33 ;
      RECT MASK 1 14.5735 7.112 14.6335 7.89 ;
      RECT MASK 1 15.0315 7.112 15.0915 7.89 ;
      RECT MASK 1 15.4895 7.112 15.5495 7.89 ;
      RECT MASK 1 15.9475 7.112 16.0075 7.89 ;
      RECT MASK 1 16.4055 7.112 16.4655 7.89 ;
      RECT MASK 1 16.8635 7.112 16.9235 7.89 ;
      RECT MASK 1 17.3215 7.112 17.3815 7.89 ;
      RECT MASK 1 17.7795 7.112 17.8395 7.89 ;
      RECT MASK 1 18.2375 7.112 18.2975 7.89 ;
      RECT MASK 1 18.6955 7.112 18.7555 7.89 ;
      RECT MASK 1 19.1535 7.112 19.2135 7.89 ;
      RECT MASK 1 19.6115 7.112 19.6715 7.89 ;
      RECT MASK 1 20.0695 7.112 20.1295 7.89 ;
      RECT MASK 1 20.5275 7.112 20.5875 7.89 ;
      RECT MASK 1 20.9855 7.112 21.0455 7.89 ;
      RECT MASK 1 21.4435 7.112 21.5035 7.89 ;
      RECT MASK 1 25.4335 7.112 25.4935 7.89 ;
      RECT MASK 1 25.8915 7.112 25.9515 7.89 ;
      RECT MASK 1 26.3495 7.112 26.4095 7.89 ;
      RECT MASK 1 26.8075 7.112 26.8675 7.89 ;
      RECT MASK 1 27.2655 7.112 27.3255 7.89 ;
      RECT MASK 1 27.7235 7.112 27.7835 7.89 ;
      RECT MASK 1 28.1815 7.112 28.2415 7.89 ;
      RECT MASK 1 28.6395 7.112 28.6995 7.89 ;
      RECT MASK 1 29.0975 7.112 29.1575 7.89 ;
      RECT MASK 1 29.5555 7.112 29.6155 7.89 ;
      RECT MASK 1 30.0135 7.112 30.0735 7.89 ;
      RECT MASK 1 30.4715 7.112 30.5315 7.89 ;
      RECT MASK 1 30.9295 7.112 30.9895 7.89 ;
      RECT MASK 1 31.3875 7.112 31.4475 7.89 ;
      RECT MASK 1 31.8455 7.112 31.9055 7.89 ;
      RECT MASK 1 32.3035 7.112 32.3635 7.89 ;
      RECT MASK 1 37.1455 7.112 37.2055 7.33 ;
      RECT MASK 1 37.3745 7.112 37.4345 7.89 ;
      RECT MASK 1 37.6035 7.112 37.6635 7.33 ;
      RECT MASK 1 37.8325 7.112 37.8925 7.89 ;
      RECT MASK 1 38.0615 7.112 38.1215 7.325 ;
      RECT MASK 1 38.5195 7.112 38.5795 7.89 ;
      RECT MASK 1 39.4355 7.112 39.4955 7.89 ;
      RECT MASK 1 40.3515 7.112 40.4115 7.89 ;
      RECT MASK 1 41.2675 7.112 41.3275 7.89 ;
      RECT MASK 1 41.7255 7.112 41.7855 7.89 ;
      RECT MASK 1 42.1835 7.112 42.2435 7.89 ;
      RECT MASK 1 42.6415 7.112 42.7015 7.89 ;
      RECT MASK 1 43.0995 7.112 43.1595 7.89 ;
      RECT MASK 1 43.5575 7.112 43.6175 7.89 ;
      RECT MASK 1 47.9615 7.238 48.0215 8.062 ;
      RECT MASK 1 74.7205 7.26 75.0405 8.176 ;
      RECT MASK 1 111.6645 7.26 111.9845 8.176 ;
      RECT MASK 1 84.9585 7.315 85.0585 7.721 ;
      RECT MASK 1 85.2905 7.315 85.3905 7.721 ;
      RECT MASK 1 85.6225 7.315 85.7225 7.721 ;
      RECT MASK 1 85.9545 7.315 86.0545 7.721 ;
      RECT MASK 1 86.2865 7.315 86.3865 7.721 ;
      RECT MASK 1 86.9505 7.315 87.0505 7.721 ;
      RECT MASK 1 87.9465 7.315 88.0465 7.721 ;
      RECT MASK 1 98.6585 7.315 98.7585 7.721 ;
      RECT MASK 1 99.6545 7.315 99.7545 7.721 ;
      RECT MASK 1 100.3185 7.315 100.4185 7.721 ;
      RECT MASK 1 100.6505 7.315 100.7505 7.721 ;
      RECT MASK 1 100.9825 7.315 101.0825 7.721 ;
      RECT MASK 1 101.3145 7.315 101.4145 7.721 ;
      RECT MASK 1 101.6465 7.315 101.7465 7.721 ;
      RECT MASK 1 48.2935 7.341 48.3535 7.959 ;
      RECT MASK 1 47.1315 7.346 47.1915 7.954 ;
      RECT MASK 1 47.4635 7.346 47.5235 7.954 ;
      RECT MASK 1 47.7955 7.346 47.8555 7.954 ;
      RECT MASK 1 3.0905 7.374 3.1505 7.89 ;
      RECT MASK 1 5.3805 7.374 5.4405 7.89 ;
      RECT MASK 1 8.5865 7.374 8.6465 7.89 ;
      RECT MASK 1 9.9605 7.374 10.0205 7.89 ;
      RECT MASK 1 36.9165 7.374 36.9765 7.89 ;
      RECT MASK 1 38.2905 7.374 38.3505 7.89 ;
      RECT MASK 1 41.4965 7.374 41.5565 7.89 ;
      RECT MASK 1 43.7865 7.374 43.8465 7.89 ;
      RECT MASK 1 60.826 7.4 60.886 8.555 ;
      RECT MASK 1 61.284 7.4 61.344 7.618 ;
      RECT MASK 1 61.742 7.4 61.802 7.618 ;
      RECT MASK 1 62.2 7.4 62.26 7.618 ;
      RECT MASK 1 62.658 7.4 62.718 7.618 ;
      RECT MASK 1 63.116 7.4 63.176 8.555 ;
      RECT MASK 1 49.6765 7.452 49.7365 8.745 ;
      RECT MASK 1 61.284 7.738 61.344 8.121 ;
      RECT MASK 1 61.742 7.738 61.802 8.121 ;
      RECT MASK 1 49.3445 7.751 49.4045 8.9845 ;
      RECT MASK 1 48.8745 7.8125 48.9345 8.9275 ;
      RECT MASK 1 58.765 7.839 58.825 8.121 ;
      RECT MASK 1 59.223 7.839 59.283 8.121 ;
      RECT MASK 1 59.681 7.839 59.741 8.121 ;
      RECT MASK 1 62.2 7.839 62.26 8.222 ;
      RECT MASK 1 62.658 7.839 62.718 8.222 ;
      RECT MASK 1 63.803 7.839 63.863 8.121 ;
      RECT MASK 1 64.261 7.839 64.321 8.121 ;
      RECT MASK 1 64.719 7.839 64.779 8.121 ;
      RECT MASK 1 79.3785 7.963 79.6985 9.929 ;
      RECT MASK 1 107.0065 7.963 107.3265 9.929 ;
      RECT MASK 1 71.1105 8.0455 71.1705 9.658 ;
      RECT MASK 1 3.0905 8.07 3.1505 8.586 ;
      RECT MASK 1 3.3195 8.07 3.3795 8.848 ;
      RECT MASK 1 3.7775 8.07 3.8375 8.848 ;
      RECT MASK 1 4.2355 8.07 4.2955 8.848 ;
      RECT MASK 1 4.6935 8.07 4.7535 8.848 ;
      RECT MASK 1 5.1515 8.07 5.2115 8.848 ;
      RECT MASK 1 5.3805 8.07 5.4405 8.586 ;
      RECT MASK 1 5.6095 8.07 5.6695 8.848 ;
      RECT MASK 1 6.5255 8.07 6.5855 8.848 ;
      RECT MASK 1 7.4415 8.07 7.5015 8.848 ;
      RECT MASK 1 8.3575 8.07 8.4175 8.848 ;
      RECT MASK 1 8.5865 8.07 8.6465 8.586 ;
      RECT MASK 1 9.0445 8.07 9.1045 8.848 ;
      RECT MASK 1 9.5025 8.07 9.5625 8.848 ;
      RECT MASK 1 9.9605 8.07 10.0205 8.586 ;
      RECT MASK 1 14.3445 8.07 14.4045 10.35 ;
      RECT MASK 1 14.5735 8.07 14.6335 8.848 ;
      RECT MASK 1 15.0315 8.07 15.0915 8.848 ;
      RECT MASK 1 15.4895 8.07 15.5495 8.848 ;
      RECT MASK 1 15.9475 8.07 16.0075 8.848 ;
      RECT MASK 1 16.4055 8.07 16.4655 8.848 ;
      RECT MASK 1 16.8635 8.07 16.9235 8.848 ;
      RECT MASK 1 17.3215 8.07 17.3815 8.848 ;
      RECT MASK 1 17.7795 8.07 17.8395 8.848 ;
      RECT MASK 1 18.2375 8.07 18.2975 8.848 ;
      RECT MASK 1 18.6955 8.07 18.7555 8.848 ;
      RECT MASK 1 19.1535 8.07 19.2135 8.848 ;
      RECT MASK 1 19.6115 8.07 19.6715 8.848 ;
      RECT MASK 1 20.0695 8.07 20.1295 8.848 ;
      RECT MASK 1 20.5275 8.07 20.5875 8.848 ;
      RECT MASK 1 20.9855 8.07 21.0455 8.848 ;
      RECT MASK 1 21.4435 8.07 21.5035 8.848 ;
      RECT MASK 1 21.6725 8.07 21.7325 10.35 ;
      RECT MASK 1 47.1315 8.074 47.1915 8.666 ;
      RECT MASK 1 47.4635 8.074 47.5235 8.666 ;
      RECT MASK 1 47.7955 8.074 47.8555 8.268 ;
      RECT MASK 1 46.7995 8.079 46.8595 8.661 ;
      RECT MASK 1 48.2935 8.079 48.3535 8.666 ;
      RECT MASK 1 48.6255 8.079 48.6855 8.661 ;
      RECT MASK 1 50.4095 8.225 50.4495 10.259 ;
      RECT MASK 1 51.0735 8.225 51.1135 10.259 ;
      RECT MASK 1 51.7375 8.225 51.7775 10.259 ;
      RECT MASK 1 52.4015 8.225 52.4415 10.259 ;
      RECT MASK 1 47.6295 8.254 47.6895 8.486 ;
      RECT MASK 1 47.9615 8.254 48.0215 8.661 ;
      RECT MASK 1 65.635 8.3225 65.695 9.378 ;
      RECT MASK 1 22.3385 8.34 22.3985 9.025 ;
      RECT MASK 1 22.5385 8.34 22.5985 9.025 ;
      RECT MASK 1 22.7385 8.34 22.7985 9.025 ;
      RECT MASK 1 22.9385 8.34 22.9985 9.025 ;
      RECT MASK 1 23.1385 8.34 23.1985 9.025 ;
      RECT MASK 1 58.765 8.342 58.825 8.842 ;
      RECT MASK 1 59.223 8.342 59.283 8.842 ;
      RECT MASK 1 59.681 8.342 59.741 8.842 ;
      RECT MASK 1 61.284 8.342 61.344 8.555 ;
      RECT MASK 1 61.742 8.342 61.802 8.555 ;
      RECT MASK 1 62.2 8.342 62.26 8.555 ;
      RECT MASK 1 62.658 8.342 62.718 8.555 ;
      RECT MASK 1 63.803 8.342 63.863 8.842 ;
      RECT MASK 1 64.261 8.342 64.321 8.842 ;
      RECT MASK 1 64.719 8.342 64.779 8.842 ;
      RECT MASK 1 67.659 8.495 67.719 9.4075 ;
      RECT MASK 1 67.888 8.495 67.948 8.966 ;
      RECT MASK 1 68.346 8.495 68.406 9.292 ;
      RECT MASK 1 68.575 8.495 68.635 8.725 ;
      RECT MASK 1 68.804 8.495 68.864 9.292 ;
      RECT MASK 1 69.033 8.495 69.093 8.725 ;
      RECT MASK 1 69.262 8.495 69.322 9.292 ;
      RECT MASK 1 69.491 8.495 69.551 8.725 ;
      RECT MASK 1 69.72 8.495 69.78 8.966 ;
      RECT MASK 1 69.949 8.495 70.009 9.292 ;
      RECT MASK 1 70.407 8.495 70.467 8.966 ;
      RECT MASK 1 70.636 8.495 70.696 9.4075 ;
      RECT MASK 1 53.7915 8.525 53.8515 9.4375 ;
      RECT MASK 1 54.0205 8.525 54.0805 8.996 ;
      RECT MASK 1 54.4785 8.525 54.5385 9.322 ;
      RECT MASK 1 54.7075 8.525 54.7675 8.755 ;
      RECT MASK 1 54.9365 8.525 54.9965 9.322 ;
      RECT MASK 1 55.1655 8.525 55.2255 8.755 ;
      RECT MASK 1 55.3945 8.525 55.4545 9.322 ;
      RECT MASK 1 55.6235 8.525 55.6835 8.996 ;
      RECT MASK 1 55.8525 8.525 55.9125 8.996 ;
      RECT MASK 1 56.0815 8.525 56.1415 9.4375 ;
      RECT MASK 1 9.2735 8.63 9.3335 8.848 ;
      RECT MASK 1 9.7315 8.63 9.7915 8.848 ;
      RECT MASK 1 8.8155 8.635 8.8755 8.848 ;
      RECT MASK 1 2.4035 8.668 2.4635 9.752 ;
      RECT MASK 1 2.8615 8.668 2.9215 9.752 ;
      RECT MASK 1 3.5485 8.668 3.6085 9.752 ;
      RECT MASK 1 4.0065 8.668 4.0665 9.305 ;
      RECT MASK 1 4.4645 8.668 4.5245 9.752 ;
      RECT MASK 1 4.9225 8.668 4.9825 9.752 ;
      RECT MASK 1 6.0675 8.668 6.1275 9.752 ;
      RECT MASK 1 6.9835 8.668 7.0435 9.752 ;
      RECT MASK 1 7.8995 8.668 7.9595 9.752 ;
      RECT MASK 1 11.3455 8.668 11.4055 9.752 ;
      RECT MASK 1 11.8035 8.668 11.8635 9.752 ;
      RECT MASK 1 12.2615 8.668 12.3215 9.752 ;
      RECT MASK 1 12.7195 8.668 12.7795 9.752 ;
      RECT MASK 1 61.971 8.67 62.031 9.1975 ;
      RECT MASK 1 61.055 8.675 61.115 9.9175 ;
      RECT MASK 1 47.6295 8.678 47.6895 9.502 ;
      RECT MASK 1 58.536 8.678 58.596 9.178 ;
      RECT MASK 1 58.994 8.678 59.054 9.178 ;
      RECT MASK 1 59.452 8.678 59.512 9.178 ;
      RECT MASK 1 59.91 8.678 59.97 9.178 ;
      RECT MASK 1 60.368 8.678 60.428 9.178 ;
      RECT MASK 1 47.9615 8.781 48.0215 9.399 ;
      RECT MASK 1 47.1315 8.786 47.1915 9.394 ;
      RECT MASK 1 47.4635 8.786 47.5235 9.394 ;
      RECT MASK 1 48.2935 8.786 48.3535 9.394 ;
      RECT MASK 1 10.8455 8.87 10.9055 9.545 ;
      RECT MASK 1 8.5865 8.875 8.6465 9.545 ;
      RECT MASK 1 63.803 8.965 63.863 9.178 ;
      RECT MASK 1 64.261 8.965 64.321 9.178 ;
      RECT MASK 1 64.719 8.965 64.779 9.178 ;
      RECT MASK 1 5.3805 8.968 5.4405 9.55 ;
      RECT MASK 1 6.2965 8.968 6.3565 9.785 ;
      RECT MASK 1 7.2125 8.968 7.2725 9.452 ;
      RECT MASK 1 31.5655 8.982 31.6255 9.4375 ;
      RECT MASK 1 39.1225 8.982 39.1825 9.4375 ;
      RECT MASK 1 62.887 8.998 62.947 10.082 ;
      RECT MASK 1 63.345 8.998 63.405 10.082 ;
      RECT MASK 1 65.177 8.998 65.237 9.755 ;
      RECT MASK 1 14.917 9.01 14.977 9.19 ;
      RECT MASK 1 15.375 9.01 15.435 9.19 ;
      RECT MASK 1 15.833 9.01 15.893 9.19 ;
      RECT MASK 1 16.291 9.01 16.351 9.19 ;
      RECT MASK 1 16.749 9.01 16.809 9.19 ;
      RECT MASK 1 17.665 9.01 17.725 9.19 ;
      RECT MASK 1 18.123 9.01 18.183 9.19 ;
      RECT MASK 1 19.039 9.01 19.099 9.19 ;
      RECT MASK 1 19.497 9.01 19.557 9.19 ;
      RECT MASK 1 19.955 9.01 20.015 9.19 ;
      RECT MASK 1 20.413 9.01 20.473 9.19 ;
      RECT MASK 1 20.871 9.01 20.931 9.19 ;
      RECT MASK 1 21.329 9.01 21.389 9.19 ;
      RECT MASK 1 32.367 9.0495 32.427 10.1015 ;
      RECT MASK 1 33.283 9.0495 33.343 10.1015 ;
      RECT MASK 1 34.199 9.0495 34.259 10.1015 ;
      RECT MASK 1 35.115 9.0495 35.175 10.1015 ;
      RECT MASK 1 36.031 9.0495 36.091 10.1015 ;
      RECT MASK 1 36.947 9.0495 37.007 10.1015 ;
      RECT MASK 1 37.863 9.0495 37.923 10.1015 ;
      RECT MASK 1 9.0445 9.069 9.1045 9.249 ;
      RECT MASK 1 9.5025 9.069 9.5625 9.249 ;
      RECT MASK 1 68.575 9.071 68.635 10.069 ;
      RECT MASK 1 69.033 9.071 69.093 10.069 ;
      RECT MASK 1 69.491 9.071 69.551 9.292 ;
      RECT MASK 1 54.7075 9.101 54.7675 10.099 ;
      RECT MASK 1 55.1655 9.101 55.2255 10.099 ;
      RECT MASK 1 11.0955 9.11 11.1555 9.351 ;
      RECT MASK 1 9.9815 9.115 10.0415 9.351 ;
      RECT MASK 1 69.72 9.193 69.78 10.069 ;
      RECT MASK 1 43.467 9.195 43.527 10.545 ;
      RECT MASK 1 8.8155 9.23 8.8755 9.752 ;
      RECT MASK 1 9.2735 9.23 9.3335 9.752 ;
      RECT MASK 1 12.9915 9.23 13.0515 9.41 ;
      RECT MASK 1 14.688 9.23 14.748 9.41 ;
      RECT MASK 1 15.146 9.23 15.206 9.41 ;
      RECT MASK 1 15.604 9.23 15.664 9.41 ;
      RECT MASK 1 16.062 9.23 16.122 9.41 ;
      RECT MASK 1 16.52 9.23 16.58 9.41 ;
      RECT MASK 1 16.978 9.23 17.038 9.41 ;
      RECT MASK 1 17.436 9.23 17.496 9.41 ;
      RECT MASK 1 18.352 9.23 18.412 9.41 ;
      RECT MASK 1 18.81 9.23 18.87 9.41 ;
      RECT MASK 1 19.726 9.23 19.786 9.41 ;
      RECT MASK 1 20.642 9.23 20.702 9.41 ;
      RECT MASK 1 21.1 9.23 21.16 9.41 ;
      RECT MASK 1 26.382 9.231 26.442 14.557 ;
      RECT MASK 1 9.7315 9.235 9.7915 9.752 ;
      RECT MASK 1 22.0365 9.235 22.0965 9.416 ;
      RECT MASK 1 32.825 9.291 32.885 9.909 ;
      RECT MASK 1 33.741 9.291 33.801 9.909 ;
      RECT MASK 1 34.657 9.291 34.717 9.909 ;
      RECT MASK 1 35.573 9.291 35.633 9.909 ;
      RECT MASK 1 36.489 9.291 36.549 9.909 ;
      RECT MASK 1 37.405 9.291 37.465 9.909 ;
      RECT MASK 1 38.321 9.291 38.381 9.909 ;
      RECT MASK 1 64.49 9.298 64.55 9.782 ;
      RECT MASK 1 49.9665 9.3 50.0065 10.77 ;
      RECT MASK 1 50.6305 9.3 50.6705 10.77 ;
      RECT MASK 1 51.2945 9.3 51.3345 10.77 ;
      RECT MASK 1 51.9585 9.3 51.9985 10.77 ;
      RECT MASK 1 52.6225 9.3 52.6625 10.77 ;
      RECT MASK 1 49.6765 9.3945 49.7365 10.353 ;
      RECT MASK 1 59.5665 9.399 59.6265 9.681 ;
      RECT MASK 1 22.5385 9.44 22.5985 10.065 ;
      RECT MASK 1 22.7385 9.44 22.7985 10.065 ;
      RECT MASK 1 22.9385 9.44 22.9985 10.065 ;
      RECT MASK 1 63.574 9.445 63.634 9.782 ;
      RECT MASK 1 4.0065 9.475 4.0665 9.752 ;
      RECT MASK 1 9.0445 9.475 9.1045 9.752 ;
      RECT MASK 1 47.1315 9.514 47.1915 10.165 ;
      RECT MASK 1 47.4635 9.514 47.5235 10.165 ;
      RECT MASK 1 48.2935 9.514 48.3535 10.165 ;
      RECT MASK 1 56.939 9.517 56.999 9.8755 ;
      RECT MASK 1 46.7995 9.519 46.8595 10.165 ;
      RECT MASK 1 47.9615 9.519 48.0215 10.165 ;
      RECT MASK 1 48.6255 9.519 48.6855 10.165 ;
      RECT MASK 1 43.1215 9.529 43.1815 10.941 ;
      RECT MASK 1 22.3385 9.531 22.3985 10.065 ;
      RECT MASK 1 23.1385 9.531 23.1985 10.065 ;
      RECT MASK 1 63.8 9.54 63.86 9.727 ;
      RECT MASK 1 5.1515 9.571 5.2115 10.35 ;
      RECT MASK 1 3.3195 9.572 3.3795 10.35 ;
      RECT MASK 1 3.7775 9.572 3.8375 10.35 ;
      RECT MASK 1 4.2355 9.572 4.2955 10.35 ;
      RECT MASK 1 4.6935 9.572 4.7535 10.35 ;
      RECT MASK 1 5.6095 9.572 5.6695 10.35 ;
      RECT MASK 1 6.5255 9.572 6.5855 10.35 ;
      RECT MASK 1 7.4415 9.572 7.5015 10.35 ;
      RECT MASK 1 9.5025 9.572 9.5625 9.79 ;
      RECT MASK 1 14.5735 9.572 14.6335 10.35 ;
      RECT MASK 1 15.0315 9.572 15.0915 10.35 ;
      RECT MASK 1 15.4895 9.572 15.5495 10.35 ;
      RECT MASK 1 15.9475 9.572 16.0075 10.35 ;
      RECT MASK 1 16.4055 9.572 16.4655 10.35 ;
      RECT MASK 1 16.8635 9.572 16.9235 10.35 ;
      RECT MASK 1 17.3215 9.572 17.3815 10.35 ;
      RECT MASK 1 17.7795 9.572 17.8395 10.35 ;
      RECT MASK 1 18.2375 9.572 18.2975 10.35 ;
      RECT MASK 1 18.6955 9.572 18.7555 10.35 ;
      RECT MASK 1 19.1535 9.572 19.2135 10.35 ;
      RECT MASK 1 19.6115 9.572 19.6715 10.35 ;
      RECT MASK 1 20.0695 9.572 20.1295 10.35 ;
      RECT MASK 1 20.5275 9.572 20.5875 10.35 ;
      RECT MASK 1 20.9855 9.572 21.0455 10.35 ;
      RECT MASK 1 21.4435 9.572 21.5035 10.35 ;
      RECT MASK 1 8.3575 9.5725 8.4175 10.35 ;
      RECT MASK 1 58.536 9.601 58.596 10.68 ;
      RECT MASK 1 60.368 9.601 60.428 10.68 ;
      RECT MASK 1 65.635 9.685 65.695 10.082 ;
      RECT MASK 1 66.101 9.685 66.161 9.9385 ;
      RECT MASK 1 47.6295 9.694 47.6895 10.165 ;
      RECT MASK 1 48.1275 9.694 48.1875 10.165 ;
      RECT MASK 1 42.7895 9.702 42.8495 11.133 ;
      RECT MASK 1 61.971 9.7625 62.031 10.68 ;
      RECT MASK 1 41.156 9.803 41.216 12.923 ;
      RECT MASK 1 3.0905 9.834 3.1505 10.35 ;
      RECT MASK 1 5.3805 9.834 5.4405 10.35 ;
      RECT MASK 1 8.5865 9.834 8.6465 10.35 ;
      RECT MASK 1 9.9605 9.834 10.0205 10.35 ;
      RECT MASK 1 68.346 9.848 68.406 10.645 ;
      RECT MASK 1 68.804 9.848 68.864 10.645 ;
      RECT MASK 1 69.262 9.848 69.322 10.645 ;
      RECT MASK 1 69.491 9.848 69.551 10.188 ;
      RECT MASK 1 69.949 9.848 70.009 10.645 ;
      RECT MASK 1 54.4785 9.878 54.5385 10.675 ;
      RECT MASK 1 54.9365 9.878 54.9965 10.675 ;
      RECT MASK 1 55.3945 9.878 55.4545 10.675 ;
      RECT MASK 1 58.994 9.902 59.054 10.68 ;
      RECT MASK 1 59.452 9.902 59.512 10.68 ;
      RECT MASK 1 59.91 9.902 59.97 10.68 ;
      RECT MASK 1 63.803 9.902 63.863 10.115 ;
      RECT MASK 1 64.261 9.902 64.321 10.115 ;
      RECT MASK 1 64.719 9.902 64.779 10.115 ;
      RECT MASK 1 65.177 9.902 65.237 10.115 ;
      RECT MASK 1 27.212 9.903 27.272 13.113 ;
      RECT MASK 1 38.832 9.903 38.892 13.156 ;
      RECT MASK 1 67.888 10.174 67.948 10.645 ;
      RECT MASK 1 70.178 10.174 70.238 10.645 ;
      RECT MASK 1 70.407 10.174 70.467 10.645 ;
      RECT MASK 1 54.0205 10.204 54.0805 10.675 ;
      RECT MASK 1 55.6235 10.204 55.6835 10.675 ;
      RECT MASK 1 55.8525 10.204 55.9125 10.675 ;
      RECT MASK 1 68.575 10.415 68.635 10.645 ;
      RECT MASK 1 69.033 10.415 69.093 10.645 ;
      RECT MASK 1 69.491 10.415 69.551 10.645 ;
      RECT MASK 1 69.72 10.415 69.78 10.645 ;
      RECT MASK 1 54.7075 10.445 54.7675 10.675 ;
      RECT MASK 1 55.1655 10.445 55.2255 10.675 ;
      RECT MASK 1 59.223 10.445 59.283 10.675 ;
      RECT MASK 1 59.681 10.445 59.741 10.675 ;
      RECT MASK 1 62.429 10.445 62.489 10.675 ;
      RECT MASK 1 62.887 10.445 62.947 10.675 ;
      RECT MASK 1 63.345 10.445 63.405 10.675 ;
      RECT MASK 1 63.803 10.445 63.863 10.675 ;
      RECT MASK 1 64.032 10.445 64.092 10.675 ;
      RECT MASK 1 64.261 10.445 64.321 10.675 ;
      RECT MASK 1 64.719 10.445 64.779 10.675 ;
      RECT MASK 1 64.948 10.445 65.008 10.675 ;
      RECT MASK 1 65.177 10.445 65.237 10.675 ;
      RECT MASK 1 65.635 10.445 65.695 10.675 ;
      RECT MASK 1 62.238 10.871 62.298 12.923 ;
      RECT MASK 1 59.914 10.967 59.974 13.019 ;
      RECT MASK 1 55.432 11.063 55.492 12.9695 ;
      RECT MASK 1 79.668 11.246 79.728 13.019 ;
      RECT MASK 1 35.512 11.253 35.572 13.113 ;
      RECT MASK 1 23.062 11.255 23.122 12.731 ;
      RECT MASK 1 42.982 11.255 43.042 12.731 ;
      RECT MASK 1 89.628 11.255 89.688 13.019 ;
      RECT MASK 1 33.022 11.33 33.082 13.27 ;
      RECT MASK 1 47.132 11.349 47.192 13.113 ;
      RECT MASK 1 10.612 11.351 10.672 12.938 ;
      RECT MASK 1 68.878 11.351 68.938 13.019 ;
      RECT MASK 1 102.078 11.351 102.138 12.977 ;
      RECT MASK 1 83.818 11.433 83.878 13.019 ;
      RECT MASK 1 28.872 11.447 28.932 12.637 ;
      RECT MASK 1 36.342 11.537 36.402 13.113 ;
      RECT MASK 1 24.722 11.543 24.782 12.635 ;
      RECT MASK 1 38.002 11.543 38.062 12.731 ;
      RECT MASK 1 78.008 11.543 78.068 13.019 ;
      RECT MASK 1 91.288 11.543 91.348 12.637 ;
      RECT MASK 1 50.452 11.637 50.512 13.113 ;
      RECT MASK 1 8.952 11.639 9.012 12.923 ;
      RECT MASK 1 67.218 11.639 67.278 13.019 ;
      RECT MASK 1 103.738 11.639 103.798 13.019 ;
      RECT MASK 1 4.626 11.76 4.706 12.416 ;
      RECT MASK 1 4.792 11.76 4.872 12.416 ;
      RECT MASK 1 4.958 11.76 5.038 12.416 ;
      RECT MASK 1 5.124 11.76 5.204 12.416 ;
      RECT MASK 1 5.29 11.76 5.37 12.416 ;
      RECT MASK 1 5.456 11.76 5.536 12.416 ;
      RECT MASK 1 5.622 11.76 5.702 12.416 ;
      RECT MASK 1 5.788 11.76 5.868 12.416 ;
      RECT MASK 1 5.954 11.76 6.034 12.416 ;
      RECT MASK 1 6.12 11.76 6.2 12.416 ;
      RECT MASK 1 6.286 11.76 6.366 12.416 ;
      RECT MASK 1 6.452 11.76 6.532 12.416 ;
      RECT MASK 1 6.618 11.76 6.698 12.416 ;
      RECT MASK 1 6.784 11.76 6.864 12.416 ;
      RECT MASK 1 6.95 11.76 7.03 12.416 ;
      RECT MASK 1 7.116 11.76 7.196 12.416 ;
      RECT MASK 1 7.282 11.76 7.362 12.416 ;
      RECT MASK 1 7.448 11.76 7.528 12.416 ;
      RECT MASK 1 7.614 11.76 7.694 12.416 ;
      RECT MASK 1 7.78 11.76 7.86 12.416 ;
      RECT MASK 1 7.946 11.76 8.026 12.416 ;
      RECT MASK 1 8.112 11.76 8.192 12.416 ;
      RECT MASK 1 8.278 11.76 8.358 12.416 ;
      RECT MASK 1 9.606 11.76 9.686 12.416 ;
      RECT MASK 1 9.772 11.76 9.852 12.416 ;
      RECT MASK 1 9.938 11.76 10.018 12.416 ;
      RECT MASK 1 11.266 11.76 11.346 12.416 ;
      RECT MASK 1 11.432 11.76 11.512 12.416 ;
      RECT MASK 1 11.598 11.76 11.678 12.416 ;
      RECT MASK 1 11.764 11.76 11.844 12.416 ;
      RECT MASK 1 11.93 11.76 12.01 12.416 ;
      RECT MASK 1 12.096 11.76 12.176 12.416 ;
      RECT MASK 1 12.262 11.76 12.342 12.416 ;
      RECT MASK 1 12.428 11.76 12.508 12.416 ;
      RECT MASK 1 12.594 11.76 12.674 12.416 ;
      RECT MASK 1 12.76 11.76 12.84 12.416 ;
      RECT MASK 1 12.926 11.76 13.006 12.416 ;
      RECT MASK 1 13.092 11.76 13.172 12.416 ;
      RECT MASK 1 13.258 11.76 13.338 12.416 ;
      RECT MASK 1 13.424 11.76 13.504 12.416 ;
      RECT MASK 1 13.59 11.76 13.67 12.416 ;
      RECT MASK 1 13.756 11.76 13.836 12.416 ;
      RECT MASK 1 13.922 11.76 14.002 12.416 ;
      RECT MASK 1 14.088 11.76 14.168 12.416 ;
      RECT MASK 1 14.254 11.76 14.334 12.416 ;
      RECT MASK 1 14.42 11.76 14.5 12.416 ;
      RECT MASK 1 14.586 11.76 14.666 12.416 ;
      RECT MASK 1 14.752 11.76 14.832 12.416 ;
      RECT MASK 1 14.918 11.76 14.998 12.416 ;
      RECT MASK 1 15.084 11.76 15.164 12.416 ;
      RECT MASK 1 15.25 11.76 15.33 12.416 ;
      RECT MASK 1 15.416 11.76 15.496 12.416 ;
      RECT MASK 1 15.582 11.76 15.662 12.416 ;
      RECT MASK 1 15.748 11.76 15.828 12.416 ;
      RECT MASK 1 15.914 11.76 15.994 12.416 ;
      RECT MASK 1 16.08 11.76 16.16 12.416 ;
      RECT MASK 1 16.246 11.76 16.326 12.416 ;
      RECT MASK 1 16.412 11.76 16.492 12.416 ;
      RECT MASK 1 16.578 11.76 16.658 12.416 ;
      RECT MASK 1 16.744 11.76 16.824 12.416 ;
      RECT MASK 1 16.91 11.76 16.99 12.416 ;
      RECT MASK 1 17.076 11.76 17.156 12.416 ;
      RECT MASK 1 17.242 11.76 17.322 12.416 ;
      RECT MASK 1 17.408 11.76 17.488 12.416 ;
      RECT MASK 1 17.574 11.76 17.654 12.416 ;
      RECT MASK 1 17.74 11.76 17.82 12.416 ;
      RECT MASK 1 17.906 11.76 17.986 12.416 ;
      RECT MASK 1 18.072 11.76 18.152 12.416 ;
      RECT MASK 1 18.238 11.76 18.318 12.416 ;
      RECT MASK 1 18.404 11.76 18.484 12.416 ;
      RECT MASK 1 18.57 11.76 18.65 12.416 ;
      RECT MASK 1 18.736 11.76 18.816 12.416 ;
      RECT MASK 1 18.902 11.76 18.982 12.416 ;
      RECT MASK 1 19.068 11.76 19.148 12.416 ;
      RECT MASK 1 19.234 11.76 19.314 12.416 ;
      RECT MASK 1 19.4 11.76 19.48 12.416 ;
      RECT MASK 1 19.566 11.76 19.646 12.416 ;
      RECT MASK 1 19.732 11.76 19.812 12.416 ;
      RECT MASK 1 19.898 11.76 19.978 12.416 ;
      RECT MASK 1 20.064 11.76 20.144 12.416 ;
      RECT MASK 1 20.23 11.76 20.31 12.416 ;
      RECT MASK 1 20.396 11.76 20.476 12.416 ;
      RECT MASK 1 20.562 11.76 20.642 12.416 ;
      RECT MASK 1 20.728 11.76 20.808 12.416 ;
      RECT MASK 1 20.894 11.76 20.974 12.416 ;
      RECT MASK 1 21.06 11.76 21.14 12.416 ;
      RECT MASK 1 21.226 11.76 21.306 12.416 ;
      RECT MASK 1 21.392 11.76 21.472 12.416 ;
      RECT MASK 1 21.558 11.76 21.638 12.416 ;
      RECT MASK 1 21.724 11.76 21.804 12.416 ;
      RECT MASK 1 21.89 11.76 21.97 12.416 ;
      RECT MASK 1 22.056 11.76 22.136 12.416 ;
      RECT MASK 1 22.222 11.76 22.302 12.5115 ;
      RECT MASK 1 22.388 11.76 22.468 12.241 ;
      RECT MASK 1 22.886 11.76 22.966 12.416 ;
      RECT MASK 1 23.218 11.76 23.298 12.416 ;
      RECT MASK 1 23.716 11.76 23.796 12.2605 ;
      RECT MASK 1 23.882 11.76 23.962 12.464 ;
      RECT MASK 1 24.048 11.76 24.128 12.2605 ;
      RECT MASK 1 24.546 11.76 24.626 12.416 ;
      RECT MASK 1 24.878 11.76 24.958 12.416 ;
      RECT MASK 1 25.376 11.76 25.456 12.241 ;
      RECT MASK 1 25.542 11.76 25.622 12.5025 ;
      RECT MASK 1 25.708 11.76 25.788 12.241 ;
      RECT MASK 1 26.206 11.76 26.286 12.416 ;
      RECT MASK 1 26.538 11.76 26.618 12.416 ;
      RECT MASK 1 27.036 11.76 27.116 12.241 ;
      RECT MASK 1 27.368 11.76 27.448 12.481 ;
      RECT MASK 1 27.534 11.76 27.614 12.241 ;
      RECT MASK 1 27.7 11.76 27.78 12.4895 ;
      RECT MASK 1 27.866 11.76 27.946 12.4245 ;
      RECT MASK 1 28.032 11.76 28.112 12.4245 ;
      RECT MASK 1 28.198 11.76 28.278 12.416 ;
      RECT MASK 1 28.696 11.76 28.776 12.241 ;
      RECT MASK 1 29.028 11.76 29.108 12.241 ;
      RECT MASK 1 29.526 11.76 29.606 12.416 ;
      RECT MASK 1 29.692 11.76 29.772 12.421 ;
      RECT MASK 1 29.858 11.76 29.938 12.4765 ;
      RECT MASK 1 30.024 11.76 30.104 12.241 ;
      RECT MASK 1 30.19 11.76 30.27 12.4715 ;
      RECT MASK 1 30.356 11.76 30.436 12.421 ;
      RECT MASK 1 30.522 11.76 30.602 12.4765 ;
      RECT MASK 1 30.688 11.76 30.768 12.241 ;
      RECT MASK 1 31.186 11.76 31.266 12.416 ;
      RECT MASK 1 31.352 11.76 31.432 12.413 ;
      RECT MASK 1 31.518 11.76 31.598 12.416 ;
      RECT MASK 1 32.016 11.76 32.096 12.241 ;
      RECT MASK 1 32.182 11.76 32.262 12.515 ;
      RECT MASK 1 32.348 11.76 32.428 12.241 ;
      RECT MASK 1 32.846 11.76 32.926 12.416 ;
      RECT MASK 1 33.178 11.76 33.258 12.416 ;
      RECT MASK 1 33.676 11.76 33.756 12.241 ;
      RECT MASK 1 33.842 11.76 33.922 12.543 ;
      RECT MASK 1 34.008 11.76 34.088 12.416 ;
      RECT MASK 1 34.506 11.76 34.586 12.241 ;
      RECT MASK 1 34.672 11.76 34.752 12.5215 ;
      RECT MASK 1 34.838 11.76 34.918 12.241 ;
      RECT MASK 1 35.336 11.76 35.416 12.416 ;
      RECT MASK 1 35.668 11.76 35.748 12.241 ;
      RECT MASK 1 36.166 11.76 36.246 12.416 ;
      RECT MASK 1 36.498 11.76 36.578 12.416 ;
      RECT MASK 1 36.996 11.76 37.076 12.241 ;
      RECT MASK 1 37.162 11.76 37.242 12.4735 ;
      RECT MASK 1 37.328 11.76 37.408 12.241 ;
      RECT MASK 1 37.826 11.76 37.906 12.416 ;
      RECT MASK 1 38.158 11.76 38.238 12.416 ;
      RECT MASK 1 38.656 11.76 38.736 12.241 ;
      RECT MASK 1 38.988 11.76 39.068 12.241 ;
      RECT MASK 1 39.486 11.76 39.566 12.416 ;
      RECT MASK 1 39.818 11.76 39.898 12.416 ;
      RECT MASK 1 40.316 11.76 40.396 12.241 ;
      RECT MASK 1 40.482 11.76 40.562 12.4855 ;
      RECT MASK 1 40.648 11.76 40.728 12.4855 ;
      RECT MASK 1 40.814 11.76 40.894 12.241 ;
      RECT MASK 1 40.98 11.76 41.06 12.4775 ;
      RECT MASK 1 41.312 11.76 41.392 12.416 ;
      RECT MASK 1 41.478 11.76 41.558 12.4765 ;
      RECT MASK 1 41.644 11.76 41.724 12.2495 ;
      RECT MASK 1 41.81 11.76 41.89 12.4755 ;
      RECT MASK 1 41.976 11.76 42.056 12.4305 ;
      RECT MASK 1 42.142 11.76 42.222 12.4755 ;
      RECT MASK 1 42.308 11.76 42.388 12.241 ;
      RECT MASK 1 42.806 11.76 42.886 12.416 ;
      RECT MASK 1 43.138 11.76 43.218 12.416 ;
      RECT MASK 1 43.636 11.76 43.716 12.241 ;
      RECT MASK 1 43.802 11.76 43.882 12.468 ;
      RECT MASK 1 43.968 11.76 44.048 12.241 ;
      RECT MASK 1 44.466 11.76 44.546 12.416 ;
      RECT MASK 1 44.632 11.76 44.712 12.4345 ;
      RECT MASK 1 44.798 11.76 44.878 12.416 ;
      RECT MASK 1 45.296 11.76 45.376 12.241 ;
      RECT MASK 1 45.628 11.76 45.708 12.416 ;
      RECT MASK 1 46.126 11.76 46.206 12.241 ;
      RECT MASK 1 46.458 11.76 46.538 12.416 ;
      RECT MASK 1 46.956 11.76 47.036 12.241 ;
      RECT MASK 1 47.288 11.76 47.368 12.241 ;
      RECT MASK 1 47.786 11.76 47.866 12.416 ;
      RECT MASK 1 47.952 11.76 48.032 12.416 ;
      RECT MASK 1 48.118 11.76 48.198 12.416 ;
      RECT MASK 1 48.616 11.76 48.696 12.241 ;
      RECT MASK 1 48.782 11.76 48.862 12.4565 ;
      RECT MASK 1 48.948 11.76 49.028 12.241 ;
      RECT MASK 1 49.446 11.76 49.526 12.416 ;
      RECT MASK 1 49.612 11.76 49.692 12.416 ;
      RECT MASK 1 49.778 11.76 49.858 12.416 ;
      RECT MASK 1 50.276 11.76 50.356 12.241 ;
      RECT MASK 1 50.608 11.76 50.688 12.241 ;
      RECT MASK 1 51.106 11.76 51.186 12.416 ;
      RECT MASK 1 51.272 11.76 51.352 12.4195 ;
      RECT MASK 1 51.438 11.76 51.518 12.416 ;
      RECT MASK 1 51.936 11.76 52.016 12.241 ;
      RECT MASK 1 52.102 11.76 52.182 12.4605 ;
      RECT MASK 1 52.268 11.76 52.348 12.241 ;
      RECT MASK 1 52.766 11.76 52.846 12.416 ;
      RECT MASK 1 52.932 11.76 53.012 12.4265 ;
      RECT MASK 1 53.098 11.76 53.178 12.416 ;
      RECT MASK 1 53.596 11.76 53.676 12.241 ;
      RECT MASK 1 53.762 11.76 53.842 12.461 ;
      RECT MASK 1 53.928 11.76 54.008 12.241 ;
      RECT MASK 1 54.426 11.76 54.506 12.416 ;
      RECT MASK 1 54.592 11.76 54.672 12.416 ;
      RECT MASK 1 54.758 11.76 54.838 12.416 ;
      RECT MASK 1 55.256 11.76 55.336 12.241 ;
      RECT MASK 1 55.588 11.76 55.668 12.241 ;
      RECT MASK 1 55.754 11.76 55.834 12.4615 ;
      RECT MASK 1 55.92 11.76 56 12.4235 ;
      RECT MASK 1 56.086 11.76 56.166 12.4235 ;
      RECT MASK 1 56.252 11.76 56.332 12.4235 ;
      RECT MASK 1 56.418 11.76 56.498 12.4235 ;
      RECT MASK 1 56.584 11.76 56.664 12.416 ;
      RECT MASK 1 57.082 11.76 57.162 12.241 ;
      RECT MASK 1 57.248 11.76 57.328 12.4605 ;
      RECT MASK 1 57.414 11.76 57.494 12.241 ;
      RECT MASK 1 57.912 11.76 57.992 12.416 ;
      RECT MASK 1 58.078 11.76 58.158 12.419 ;
      RECT MASK 1 58.244 11.76 58.324 12.416 ;
      RECT MASK 1 58.742 11.76 58.822 12.241 ;
      RECT MASK 1 58.908 11.76 58.988 12.541 ;
      RECT MASK 1 59.074 11.76 59.154 12.241 ;
      RECT MASK 1 59.572 11.76 59.652 12.416 ;
      RECT MASK 1 59.738 11.76 59.818 12.541 ;
      RECT MASK 1 60.07 11.76 60.15 12.241 ;
      RECT MASK 1 60.236 11.76 60.316 12.4615 ;
      RECT MASK 1 60.402 11.76 60.482 12.448 ;
      RECT MASK 1 60.568 11.76 60.648 12.448 ;
      RECT MASK 1 60.734 11.76 60.814 12.241 ;
      RECT MASK 1 61.232 11.76 61.312 12.416 ;
      RECT MASK 1 61.398 11.76 61.478 12.417 ;
      RECT MASK 1 61.564 11.76 61.644 12.416 ;
      RECT MASK 1 62.062 11.76 62.142 12.241 ;
      RECT MASK 1 62.394 11.76 62.474 12.4615 ;
      RECT MASK 1 62.56 11.76 62.64 12.241 ;
      RECT MASK 1 62.726 11.76 62.806 12.4685 ;
      RECT MASK 1 62.892 11.76 62.972 12.423 ;
      RECT MASK 1 63.058 11.76 63.138 12.423 ;
      RECT MASK 1 63.224 11.76 63.304 12.416 ;
      RECT MASK 1 63.722 11.76 63.802 12.241 ;
      RECT MASK 1 63.888 11.76 63.968 12.444 ;
      RECT MASK 1 64.054 11.76 64.134 12.241 ;
      RECT MASK 1 64.552 11.76 64.632 12.416 ;
      RECT MASK 1 64.718 11.76 64.798 12.416 ;
      RECT MASK 1 64.884 11.76 64.964 12.416 ;
      RECT MASK 1 65.382 11.76 65.462 12.241 ;
      RECT MASK 1 65.548 11.76 65.628 12.4535 ;
      RECT MASK 1 65.714 11.76 65.794 12.241 ;
      RECT MASK 1 66.212 11.76 66.292 12.416 ;
      RECT MASK 1 66.378 11.76 66.458 12.415 ;
      RECT MASK 1 66.544 11.76 66.624 12.416 ;
      RECT MASK 1 67.042 11.76 67.122 12.241 ;
      RECT MASK 1 67.374 11.76 67.454 12.241 ;
      RECT MASK 1 67.872 11.76 67.952 12.416 ;
      RECT MASK 1 68.038 11.76 68.118 12.241 ;
      RECT MASK 1 68.204 11.76 68.284 12.416 ;
      RECT MASK 1 68.702 11.76 68.782 12.241 ;
      RECT MASK 1 69.034 11.76 69.114 12.241 ;
      RECT MASK 1 69.532 11.76 69.612 12.416 ;
      RECT MASK 1 69.698 11.76 69.778 12.241 ;
      RECT MASK 1 69.864 11.76 69.944 12.416 ;
      RECT MASK 1 70.362 11.76 70.442 12.241 ;
      RECT MASK 1 70.528 11.76 70.608 12.456 ;
      RECT MASK 1 70.694 11.76 70.774 12.241 ;
      RECT MASK 1 71.192 11.76 71.272 12.416 ;
      RECT MASK 1 71.358 11.76 71.438 12.417 ;
      RECT MASK 1 71.524 11.76 71.604 12.416 ;
      RECT MASK 1 72.022 11.76 72.102 12.241 ;
      RECT MASK 1 72.188 11.76 72.268 12.4575 ;
      RECT MASK 1 72.354 11.76 72.434 12.241 ;
      RECT MASK 1 72.852 11.76 72.932 12.416 ;
      RECT MASK 1 73.018 11.76 73.098 12.417 ;
      RECT MASK 1 73.184 11.76 73.264 12.417 ;
      RECT MASK 1 73.35 11.76 73.43 12.25 ;
      RECT MASK 1 73.516 11.76 73.596 12.416 ;
      RECT MASK 1 73.682 11.76 73.762 12.416 ;
      RECT MASK 1 73.848 11.76 73.928 12.416 ;
      RECT MASK 1 74.014 11.76 74.094 12.416 ;
      RECT MASK 1 74.18 11.76 74.26 12.416 ;
      RECT MASK 1 74.346 11.76 74.426 12.416 ;
      RECT MASK 1 74.512 11.76 74.592 12.416 ;
      RECT MASK 1 74.678 11.76 74.758 12.416 ;
      RECT MASK 1 74.844 11.76 74.924 12.416 ;
      RECT MASK 1 75.01 11.76 75.09 12.416 ;
      RECT MASK 1 75.176 11.76 75.256 12.416 ;
      RECT MASK 1 75.342 11.76 75.422 12.416 ;
      RECT MASK 1 75.508 11.76 75.588 12.416 ;
      RECT MASK 1 75.674 11.76 75.754 12.416 ;
      RECT MASK 1 75.84 11.76 75.92 12.416 ;
      RECT MASK 1 76.006 11.76 76.086 12.416 ;
      RECT MASK 1 76.172 11.76 76.252 12.416 ;
      RECT MASK 1 76.338 11.76 76.418 12.416 ;
      RECT MASK 1 76.504 11.76 76.584 12.416 ;
      RECT MASK 1 76.67 11.76 76.75 12.416 ;
      RECT MASK 1 76.836 11.76 76.916 12.416 ;
      RECT MASK 1 77.002 11.76 77.082 12.416 ;
      RECT MASK 1 77.168 11.76 77.248 12.464 ;
      RECT MASK 1 77.334 11.76 77.414 12.241 ;
      RECT MASK 1 77.832 11.76 77.912 12.416 ;
      RECT MASK 1 78.164 11.76 78.244 12.416 ;
      RECT MASK 1 78.662 11.76 78.742 12.241 ;
      RECT MASK 1 78.828 11.76 78.908 12.4785 ;
      RECT MASK 1 78.994 11.76 79.074 12.241 ;
      RECT MASK 1 79.492 11.76 79.572 12.416 ;
      RECT MASK 1 79.824 11.76 79.904 12.416 ;
      RECT MASK 1 80.322 11.76 80.402 12.241 ;
      RECT MASK 1 80.488 11.76 80.568 12.4575 ;
      RECT MASK 1 80.654 11.76 80.734 12.421 ;
      RECT MASK 1 80.82 11.76 80.9 12.424 ;
      RECT MASK 1 80.986 11.76 81.066 12.421 ;
      RECT MASK 1 81.152 11.76 81.232 12.421 ;
      RECT MASK 1 81.318 11.76 81.398 12.421 ;
      RECT MASK 1 81.484 11.76 81.564 12.421 ;
      RECT MASK 1 81.65 11.76 81.73 12.421 ;
      RECT MASK 1 81.816 11.76 81.896 12.421 ;
      RECT MASK 1 81.982 11.76 82.062 12.421 ;
      RECT MASK 1 82.148 11.76 82.228 12.421 ;
      RECT MASK 1 82.314 11.76 82.394 12.421 ;
      RECT MASK 1 82.48 11.76 82.56 12.421 ;
      RECT MASK 1 82.646 11.76 82.726 12.421 ;
      RECT MASK 1 82.812 11.76 82.892 12.421 ;
      RECT MASK 1 82.978 11.76 83.058 12.421 ;
      RECT MASK 1 83.144 11.76 83.224 12.416 ;
      RECT MASK 1 83.642 11.76 83.722 12.241 ;
      RECT MASK 1 83.974 11.76 84.054 12.241 ;
      RECT MASK 1 84.472 11.76 84.552 12.416 ;
      RECT MASK 1 84.638 11.76 84.718 12.416 ;
      RECT MASK 1 84.804 11.76 84.884 12.416 ;
      RECT MASK 1 84.97 11.76 85.05 12.416 ;
      RECT MASK 1 85.136 11.76 85.216 12.416 ;
      RECT MASK 1 85.302 11.76 85.382 12.416 ;
      RECT MASK 1 85.468 11.76 85.548 12.416 ;
      RECT MASK 1 85.634 11.76 85.714 12.416 ;
      RECT MASK 1 85.8 11.76 85.88 12.416 ;
      RECT MASK 1 85.966 11.76 86.046 12.416 ;
      RECT MASK 1 86.132 11.76 86.212 12.416 ;
      RECT MASK 1 86.298 11.76 86.378 12.416 ;
      RECT MASK 1 86.464 11.76 86.544 12.416 ;
      RECT MASK 1 86.63 11.76 86.71 12.416 ;
      RECT MASK 1 86.796 11.76 86.876 12.416 ;
      RECT MASK 1 86.962 11.76 87.042 12.416 ;
      RECT MASK 1 87.128 11.76 87.208 12.416 ;
      RECT MASK 1 87.294 11.76 87.374 12.416 ;
      RECT MASK 1 87.46 11.76 87.54 12.416 ;
      RECT MASK 1 87.626 11.76 87.706 12.416 ;
      RECT MASK 1 87.792 11.76 87.872 12.416 ;
      RECT MASK 1 87.958 11.76 88.038 12.416 ;
      RECT MASK 1 88.124 11.76 88.204 12.416 ;
      RECT MASK 1 88.29 11.76 88.37 12.416 ;
      RECT MASK 1 88.456 11.76 88.536 12.416 ;
      RECT MASK 1 88.622 11.76 88.702 12.416 ;
      RECT MASK 1 88.788 11.76 88.868 12.4645 ;
      RECT MASK 1 88.954 11.76 89.034 12.241 ;
      RECT MASK 1 89.452 11.76 89.532 12.416 ;
      RECT MASK 1 89.784 11.76 89.864 12.416 ;
      RECT MASK 1 90.282 11.76 90.362 12.241 ;
      RECT MASK 1 90.448 11.76 90.528 12.4355 ;
      RECT MASK 1 90.614 11.76 90.694 12.241 ;
      RECT MASK 1 91.112 11.76 91.192 12.416 ;
      RECT MASK 1 91.444 11.76 91.524 12.416 ;
      RECT MASK 1 91.942 11.76 92.022 12.241 ;
      RECT MASK 1 92.108 11.76 92.188 12.471 ;
      RECT MASK 1 92.274 11.76 92.354 12.416 ;
      RECT MASK 1 92.44 11.76 92.52 12.416 ;
      RECT MASK 1 92.606 11.76 92.686 12.416 ;
      RECT MASK 1 92.772 11.76 92.852 12.416 ;
      RECT MASK 1 92.938 11.76 93.018 12.416 ;
      RECT MASK 1 93.104 11.76 93.184 12.416 ;
      RECT MASK 1 93.27 11.76 93.35 12.416 ;
      RECT MASK 1 93.436 11.76 93.516 12.416 ;
      RECT MASK 1 93.602 11.76 93.682 12.416 ;
      RECT MASK 1 93.768 11.76 93.848 12.416 ;
      RECT MASK 1 93.934 11.76 94.014 12.416 ;
      RECT MASK 1 94.1 11.76 94.18 12.416 ;
      RECT MASK 1 94.266 11.76 94.346 12.416 ;
      RECT MASK 1 94.432 11.76 94.512 12.416 ;
      RECT MASK 1 94.598 11.76 94.678 12.416 ;
      RECT MASK 1 94.764 11.76 94.844 12.416 ;
      RECT MASK 1 94.93 11.76 95.01 12.416 ;
      RECT MASK 1 95.096 11.76 95.176 12.416 ;
      RECT MASK 1 95.262 11.76 95.342 12.416 ;
      RECT MASK 1 95.428 11.76 95.508 12.416 ;
      RECT MASK 1 95.594 11.76 95.674 12.416 ;
      RECT MASK 1 95.76 11.76 95.84 12.416 ;
      RECT MASK 1 95.926 11.76 96.006 12.416 ;
      RECT MASK 1 96.092 11.76 96.172 12.416 ;
      RECT MASK 1 96.258 11.76 96.338 12.416 ;
      RECT MASK 1 96.424 11.76 96.504 12.416 ;
      RECT MASK 1 96.59 11.76 96.67 12.416 ;
      RECT MASK 1 96.756 11.76 96.836 12.416 ;
      RECT MASK 1 96.922 11.76 97.002 12.416 ;
      RECT MASK 1 97.088 11.76 97.168 12.416 ;
      RECT MASK 1 97.254 11.76 97.334 12.416 ;
      RECT MASK 1 97.42 11.76 97.5 12.416 ;
      RECT MASK 1 97.586 11.76 97.666 12.416 ;
      RECT MASK 1 97.752 11.76 97.832 12.416 ;
      RECT MASK 1 97.918 11.76 97.998 12.416 ;
      RECT MASK 1 98.084 11.76 98.164 12.416 ;
      RECT MASK 1 98.25 11.76 98.33 12.416 ;
      RECT MASK 1 98.416 11.76 98.496 12.416 ;
      RECT MASK 1 98.582 11.76 98.662 12.416 ;
      RECT MASK 1 98.748 11.76 98.828 12.416 ;
      RECT MASK 1 98.914 11.76 98.994 12.416 ;
      RECT MASK 1 99.08 11.76 99.16 12.416 ;
      RECT MASK 1 99.246 11.76 99.326 12.416 ;
      RECT MASK 1 99.412 11.76 99.492 12.416 ;
      RECT MASK 1 99.578 11.76 99.658 12.416 ;
      RECT MASK 1 99.744 11.76 99.824 12.416 ;
      RECT MASK 1 99.91 11.76 99.99 12.416 ;
      RECT MASK 1 100.076 11.76 100.156 12.416 ;
      RECT MASK 1 100.242 11.76 100.322 12.416 ;
      RECT MASK 1 100.408 11.76 100.488 12.416 ;
      RECT MASK 1 100.574 11.76 100.654 12.416 ;
      RECT MASK 1 100.74 11.76 100.82 12.416 ;
      RECT MASK 1 100.906 11.76 100.986 12.416 ;
      RECT MASK 1 101.072 11.76 101.152 12.416 ;
      RECT MASK 1 101.238 11.76 101.318 12.416 ;
      RECT MASK 1 101.404 11.76 101.484 12.416 ;
      RECT MASK 1 101.902 11.76 101.982 12.241 ;
      RECT MASK 1 102.234 11.76 102.314 12.241 ;
      RECT MASK 1 102.732 11.76 102.812 12.416 ;
      RECT MASK 1 102.898 11.76 102.978 12.416 ;
      RECT MASK 1 103.064 11.76 103.144 12.416 ;
      RECT MASK 1 103.562 11.76 103.642 12.241 ;
      RECT MASK 1 103.894 11.76 103.974 12.241 ;
      RECT MASK 1 104.392 11.76 104.472 12.416 ;
      RECT MASK 1 104.558 11.76 104.638 12.416 ;
      RECT MASK 1 104.724 11.76 104.804 12.416 ;
      RECT MASK 1 104.89 11.76 104.97 12.416 ;
      RECT MASK 1 105.056 11.76 105.136 12.416 ;
      RECT MASK 1 105.222 11.76 105.302 12.416 ;
      RECT MASK 1 105.388 11.76 105.468 12.416 ;
      RECT MASK 1 105.554 11.76 105.634 12.416 ;
      RECT MASK 1 105.72 11.76 105.8 12.416 ;
      RECT MASK 1 105.886 11.76 105.966 12.416 ;
      RECT MASK 1 106.052 11.76 106.132 12.416 ;
      RECT MASK 1 106.218 11.76 106.298 12.416 ;
      RECT MASK 1 106.384 11.76 106.464 12.416 ;
      RECT MASK 1 106.55 11.76 106.63 12.416 ;
      RECT MASK 1 106.716 11.76 106.796 12.416 ;
      RECT MASK 1 106.882 11.76 106.962 12.416 ;
      RECT MASK 1 107.048 11.76 107.128 12.416 ;
      RECT MASK 1 107.214 11.76 107.294 12.416 ;
      RECT MASK 1 107.38 11.76 107.46 12.416 ;
      RECT MASK 1 107.546 11.76 107.626 12.416 ;
      RECT MASK 1 107.712 11.76 107.792 12.416 ;
      RECT MASK 1 107.878 11.76 107.958 12.416 ;
      RECT MASK 1 108.044 11.76 108.124 12.416 ;
      RECT MASK 1 108.21 11.76 108.29 12.416 ;
      RECT MASK 1 108.376 11.76 108.456 12.416 ;
      RECT MASK 1 108.542 11.76 108.622 12.416 ;
      RECT MASK 1 108.708 11.76 108.788 12.416 ;
      RECT MASK 1 108.874 11.76 108.954 12.416 ;
      RECT MASK 1 109.04 11.76 109.12 12.416 ;
      RECT MASK 1 109.206 11.76 109.286 12.416 ;
      RECT MASK 1 109.372 11.76 109.452 12.416 ;
      RECT MASK 1 109.538 11.76 109.618 12.416 ;
      RECT MASK 1 109.704 11.76 109.784 12.416 ;
      RECT MASK 1 109.87 11.76 109.95 12.416 ;
      RECT MASK 1 110.036 11.76 110.116 12.416 ;
      RECT MASK 1 110.202 11.76 110.282 12.416 ;
      RECT MASK 1 110.368 11.76 110.448 12.416 ;
      RECT MASK 1 110.534 11.76 110.614 12.416 ;
      RECT MASK 1 110.7 11.76 110.78 12.416 ;
      RECT MASK 1 110.866 11.76 110.946 12.416 ;
      RECT MASK 1 111.032 11.76 111.112 12.416 ;
      RECT MASK 1 111.198 11.76 111.278 12.416 ;
      RECT MASK 1 111.364 11.76 111.444 12.416 ;
      RECT MASK 1 8.288 12.536 8.348 13.144 ;
      RECT MASK 1 8.62 12.536 8.68 13.144 ;
      RECT MASK 1 9.284 12.536 9.344 13.144 ;
      RECT MASK 1 9.616 12.536 9.676 13.144 ;
      RECT MASK 1 9.948 12.536 10.008 13.144 ;
      RECT MASK 1 10.28 12.536 10.34 13.144 ;
      RECT MASK 1 10.944 12.536 11.004 13.144 ;
      RECT MASK 1 11.276 12.536 11.336 13.144 ;
      RECT MASK 1 22.564 12.536 22.624 13.144 ;
      RECT MASK 1 22.896 12.536 22.956 13.144 ;
      RECT MASK 1 23.228 12.536 23.288 13.144 ;
      RECT MASK 1 23.56 12.536 23.62 13.144 ;
      RECT MASK 1 24.224 12.536 24.284 13.144 ;
      RECT MASK 1 24.556 12.536 24.616 13.144 ;
      RECT MASK 1 24.888 12.536 24.948 13.144 ;
      RECT MASK 1 25.22 12.536 25.28 13.144 ;
      RECT MASK 1 25.884 12.536 25.944 13.144 ;
      RECT MASK 1 26.216 12.536 26.276 13.144 ;
      RECT MASK 1 26.548 12.536 26.608 13.144 ;
      RECT MASK 1 26.88 12.536 26.94 13.144 ;
      RECT MASK 1 28.208 12.536 28.268 13.144 ;
      RECT MASK 1 28.54 12.536 28.6 13.144 ;
      RECT MASK 1 29.204 12.536 29.264 13.144 ;
      RECT MASK 1 29.536 12.536 29.596 13.144 ;
      RECT MASK 1 30.864 12.536 30.924 13.144 ;
      RECT MASK 1 31.196 12.536 31.256 13.144 ;
      RECT MASK 1 31.528 12.536 31.588 13.144 ;
      RECT MASK 1 31.86 12.536 31.92 13.144 ;
      RECT MASK 1 32.524 12.536 32.584 13.144 ;
      RECT MASK 1 32.856 12.536 32.916 13.144 ;
      RECT MASK 1 33.188 12.536 33.248 13.144 ;
      RECT MASK 1 33.52 12.536 33.58 13.144 ;
      RECT MASK 1 34.018 12.536 34.078 13.144 ;
      RECT MASK 1 34.35 12.536 34.41 13.144 ;
      RECT MASK 1 35.014 12.536 35.074 13.144 ;
      RECT MASK 1 35.346 12.536 35.406 13.144 ;
      RECT MASK 1 35.844 12.536 35.904 13.144 ;
      RECT MASK 1 36.176 12.536 36.236 13.144 ;
      RECT MASK 1 36.508 12.536 36.568 13.144 ;
      RECT MASK 1 36.84 12.536 36.9 13.144 ;
      RECT MASK 1 37.504 12.536 37.564 13.144 ;
      RECT MASK 1 37.836 12.536 37.896 13.144 ;
      RECT MASK 1 38.168 12.536 38.228 13.144 ;
      RECT MASK 1 38.5 12.536 38.56 13.144 ;
      RECT MASK 1 39.164 12.536 39.224 13.144 ;
      RECT MASK 1 39.496 12.536 39.556 13.144 ;
      RECT MASK 1 39.828 12.536 39.888 13.144 ;
      RECT MASK 1 40.16 12.536 40.22 13.144 ;
      RECT MASK 1 42.484 12.536 42.544 13.144 ;
      RECT MASK 1 42.816 12.536 42.876 13.144 ;
      RECT MASK 1 43.148 12.536 43.208 13.144 ;
      RECT MASK 1 43.48 12.536 43.54 13.144 ;
      RECT MASK 1 44.144 12.536 44.204 13.144 ;
      RECT MASK 1 44.476 12.536 44.536 13.144 ;
      RECT MASK 1 44.808 12.536 44.868 13.144 ;
      RECT MASK 1 45.14 12.536 45.2 13.144 ;
      RECT MASK 1 45.638 12.536 45.698 13.144 ;
      RECT MASK 1 45.97 12.536 46.03 13.144 ;
      RECT MASK 1 46.468 12.536 46.528 13.144 ;
      RECT MASK 1 46.8 12.536 46.86 13.144 ;
      RECT MASK 1 47.464 12.536 47.524 13.144 ;
      RECT MASK 1 47.796 12.536 47.856 13.144 ;
      RECT MASK 1 48.128 12.536 48.188 13.144 ;
      RECT MASK 1 48.46 12.536 48.52 13.144 ;
      RECT MASK 1 49.124 12.536 49.184 13.144 ;
      RECT MASK 1 49.456 12.536 49.516 13.144 ;
      RECT MASK 1 49.788 12.536 49.848 13.144 ;
      RECT MASK 1 50.12 12.536 50.18 13.144 ;
      RECT MASK 1 50.784 12.536 50.844 13.144 ;
      RECT MASK 1 51.116 12.536 51.176 13.144 ;
      RECT MASK 1 51.448 12.536 51.508 13.144 ;
      RECT MASK 1 51.78 12.536 51.84 13.144 ;
      RECT MASK 1 52.444 12.536 52.504 13.144 ;
      RECT MASK 1 52.776 12.536 52.836 13.144 ;
      RECT MASK 1 53.108 12.536 53.168 13.144 ;
      RECT MASK 1 53.44 12.536 53.5 13.144 ;
      RECT MASK 1 54.104 12.536 54.164 13.144 ;
      RECT MASK 1 54.436 12.536 54.496 13.144 ;
      RECT MASK 1 54.768 12.536 54.828 13.144 ;
      RECT MASK 1 55.1 12.536 55.16 13.144 ;
      RECT MASK 1 56.594 12.536 56.654 13.144 ;
      RECT MASK 1 56.926 12.536 56.986 13.144 ;
      RECT MASK 1 57.59 12.536 57.65 13.144 ;
      RECT MASK 1 57.922 12.536 57.982 13.144 ;
      RECT MASK 1 58.254 12.536 58.314 13.144 ;
      RECT MASK 1 58.586 12.536 58.646 13.144 ;
      RECT MASK 1 59.25 12.536 59.31 13.144 ;
      RECT MASK 1 59.582 12.536 59.642 13.144 ;
      RECT MASK 1 60.91 12.536 60.97 13.144 ;
      RECT MASK 1 61.242 12.536 61.302 13.144 ;
      RECT MASK 1 61.574 12.536 61.634 13.144 ;
      RECT MASK 1 61.906 12.536 61.966 13.144 ;
      RECT MASK 1 63.234 12.536 63.294 13.144 ;
      RECT MASK 1 63.566 12.536 63.626 13.144 ;
      RECT MASK 1 64.23 12.536 64.29 13.144 ;
      RECT MASK 1 64.562 12.536 64.622 13.144 ;
      RECT MASK 1 64.894 12.536 64.954 13.144 ;
      RECT MASK 1 65.226 12.536 65.286 13.144 ;
      RECT MASK 1 65.89 12.536 65.95 13.144 ;
      RECT MASK 1 66.222 12.536 66.282 13.144 ;
      RECT MASK 1 66.554 12.536 66.614 13.144 ;
      RECT MASK 1 66.886 12.536 66.946 13.144 ;
      RECT MASK 1 67.55 12.536 67.61 13.144 ;
      RECT MASK 1 67.882 12.536 67.942 13.144 ;
      RECT MASK 1 68.214 12.536 68.274 13.144 ;
      RECT MASK 1 68.546 12.536 68.606 13.144 ;
      RECT MASK 1 69.21 12.536 69.27 13.144 ;
      RECT MASK 1 69.542 12.536 69.602 13.144 ;
      RECT MASK 1 69.874 12.536 69.934 13.144 ;
      RECT MASK 1 70.206 12.536 70.266 13.144 ;
      RECT MASK 1 70.87 12.536 70.93 13.144 ;
      RECT MASK 1 71.202 12.536 71.262 13.144 ;
      RECT MASK 1 71.534 12.536 71.594 13.144 ;
      RECT MASK 1 71.866 12.536 71.926 13.144 ;
      RECT MASK 1 72.53 12.536 72.59 13.144 ;
      RECT MASK 1 72.862 12.536 72.922 13.144 ;
      RECT MASK 1 77.51 12.536 77.57 13.144 ;
      RECT MASK 1 77.842 12.536 77.902 13.144 ;
      RECT MASK 1 78.174 12.536 78.234 13.144 ;
      RECT MASK 1 78.506 12.536 78.566 13.144 ;
      RECT MASK 1 79.17 12.536 79.23 13.144 ;
      RECT MASK 1 79.502 12.536 79.562 13.144 ;
      RECT MASK 1 79.834 12.536 79.894 13.144 ;
      RECT MASK 1 80.166 12.536 80.226 13.144 ;
      RECT MASK 1 83.154 12.536 83.214 13.144 ;
      RECT MASK 1 83.486 12.536 83.546 13.144 ;
      RECT MASK 1 84.15 12.536 84.21 13.144 ;
      RECT MASK 1 84.482 12.536 84.542 13.144 ;
      RECT MASK 1 89.13 12.536 89.19 13.144 ;
      RECT MASK 1 89.462 12.536 89.522 13.144 ;
      RECT MASK 1 89.794 12.536 89.854 13.144 ;
      RECT MASK 1 90.126 12.536 90.186 13.144 ;
      RECT MASK 1 90.79 12.536 90.85 13.144 ;
      RECT MASK 1 91.122 12.536 91.182 13.144 ;
      RECT MASK 1 91.454 12.536 91.514 13.144 ;
      RECT MASK 1 91.786 12.536 91.846 13.144 ;
      RECT MASK 1 101.414 12.536 101.474 13.144 ;
      RECT MASK 1 101.746 12.536 101.806 13.144 ;
      RECT MASK 1 102.41 12.536 102.47 13.144 ;
      RECT MASK 1 102.742 12.536 102.802 13.144 ;
      RECT MASK 1 103.074 12.536 103.134 13.144 ;
      RECT MASK 1 103.406 12.536 103.466 13.144 ;
      RECT MASK 1 104.07 12.536 104.13 13.144 ;
      RECT MASK 1 104.402 12.536 104.462 13.144 ;
      RECT MASK 1 40.99 12.659 41.05 13.113 ;
      RECT MASK 1 48.792 12.659 48.852 13.113 ;
      RECT MASK 1 60.578 12.661 60.638 14.935 ;
      RECT MASK 1 30.2 12.685 30.26 13.113 ;
      RECT MASK 1 40.658 12.685 40.718 13.113 ;
      RECT MASK 1 27.378 12.687 27.438 12.993 ;
      RECT MASK 1 41.488 12.687 41.548 12.993 ;
      RECT MASK 1 55.764 12.687 55.824 13.019 ;
      RECT MASK 1 60.246 12.687 60.306 12.993 ;
      RECT MASK 1 62.404 12.687 62.464 13.142 ;
      RECT MASK 1 59.748 12.853 59.808 13.113 ;
      RECT MASK 1 54.6015 12.949 54.6615 13.211 ;
      RECT MASK 1 70.538 12.949 70.598 14.453 ;
      RECT MASK 1 4.387 13.0025 4.447 14.5975 ;
      RECT MASK 1 111.623 13.0025 111.683 14.5975 ;
      RECT MASK 1 63.068 13.014 63.128 14.935 ;
      RECT MASK 1 73.028 13.041 73.088 15.033 ;
      RECT MASK 1 24.722 13.043 24.782 14.939 ;
      RECT MASK 1 31.362 13.043 31.422 14.557 ;
      RECT MASK 1 33.852 13.043 33.912 14.557 ;
      RECT MASK 1 42.152 13.043 42.212 14.557 ;
      RECT MASK 1 51.282 13.043 51.342 14.459 ;
      RECT MASK 1 64.728 13.043 64.788 16.477 ;
      RECT MASK 1 8.952 13.141 9.012 14.939 ;
      RECT MASK 1 10.612 13.141 10.672 16.763 ;
      RECT MASK 1 14.762 13.141 14.822 16.763 ;
      RECT MASK 1 16.422 13.141 16.482 16.763 ;
      RECT MASK 1 18.082 13.141 18.142 16.763 ;
      RECT MASK 1 18.912 13.141 18.972 16.763 ;
      RECT MASK 1 23.062 13.141 23.122 16.763 ;
      RECT MASK 1 28.042 13.141 28.102 16.763 ;
      RECT MASK 1 29.702 13.141 29.762 16.763 ;
      RECT MASK 1 34.682 13.141 34.742 14.939 ;
      RECT MASK 1 38.002 13.141 38.062 16.763 ;
      RECT MASK 1 41.322 13.141 41.382 16.763 ;
      RECT MASK 1 42.982 13.141 43.042 16.763 ;
      RECT MASK 1 44.642 13.141 44.702 16.859 ;
      RECT MASK 1 46.302 13.141 46.362 14.557 ;
      RECT MASK 1 47.962 13.141 48.022 14.459 ;
      RECT MASK 1 49.622 13.141 49.682 16.763 ;
      RECT MASK 1 57.258 13.141 57.318 14.453 ;
      RECT MASK 1 58.088 13.141 58.148 14.747 ;
      RECT MASK 1 61.408 13.141 61.468 16.571 ;
      RECT MASK 1 65.558 13.141 65.618 14.651 ;
      RECT MASK 1 67.218 13.141 67.278 14.557 ;
      RECT MASK 1 68.048 13.141 68.108 16.763 ;
      RECT MASK 1 69.708 13.141 69.768 16.763 ;
      RECT MASK 1 72.198 13.141 72.258 16.763 ;
      RECT MASK 1 76.348 13.141 76.408 14.939 ;
      RECT MASK 1 79.668 13.141 79.728 16.763 ;
      RECT MASK 1 84.648 13.141 84.708 16.763 ;
      RECT MASK 1 89.628 13.141 89.688 14.939 ;
      RECT MASK 1 91.288 13.141 91.348 16.763 ;
      RECT MASK 1 94.608 13.141 94.668 16.763 ;
      RECT MASK 1 96.268 13.141 96.328 16.763 ;
      RECT MASK 1 97.928 13.141 97.988 16.763 ;
      RECT MASK 1 104.568 13.145 104.628 16.763 ;
      RECT MASK 1 107.888 13.145 107.948 16.661 ;
      RECT MASK 1 110.378 13.145 110.438 14.843 ;
      RECT MASK 1 102.078 13.1525 102.138 14.939 ;
      RECT MASK 1 4.636 13.264 4.696 14.336 ;
      RECT MASK 1 4.802 13.264 4.862 14.336 ;
      RECT MASK 1 4.968 13.264 5.028 14.336 ;
      RECT MASK 1 5.466 13.264 5.526 14.161 ;
      RECT MASK 1 5.632 13.264 5.692 14.161 ;
      RECT MASK 1 5.798 13.264 5.858 14.161 ;
      RECT MASK 1 6.296 13.264 6.356 14.336 ;
      RECT MASK 1 6.462 13.264 6.522 14.161 ;
      RECT MASK 1 6.628 13.264 6.688 14.336 ;
      RECT MASK 1 7.126 13.264 7.186 14.161 ;
      RECT MASK 1 7.292 13.264 7.352 14.161 ;
      RECT MASK 1 7.458 13.264 7.518 14.161 ;
      RECT MASK 1 7.956 13.264 8.016 14.336 ;
      RECT MASK 1 8.122 13.264 8.182 14.161 ;
      RECT MASK 1 8.288 13.264 8.348 14.336 ;
      RECT MASK 1 9.616 13.264 9.676 14.336 ;
      RECT MASK 1 9.948 13.264 10.008 14.336 ;
      RECT MASK 1 11.276 13.264 11.336 14.336 ;
      RECT MASK 1 11.608 13.264 11.668 14.336 ;
      RECT MASK 1 12.106 13.264 12.166 14.161 ;
      RECT MASK 1 12.272 13.264 12.332 14.161 ;
      RECT MASK 1 12.438 13.264 12.498 14.161 ;
      RECT MASK 1 12.936 13.264 12.996 14.336 ;
      RECT MASK 1 13.102 13.264 13.162 14.161 ;
      RECT MASK 1 13.268 13.264 13.328 14.336 ;
      RECT MASK 1 13.766 13.264 13.826 14.161 ;
      RECT MASK 1 13.932 13.264 13.992 14.161 ;
      RECT MASK 1 14.098 13.264 14.158 14.161 ;
      RECT MASK 1 14.596 13.264 14.656 14.336 ;
      RECT MASK 1 14.928 13.264 14.988 14.336 ;
      RECT MASK 1 15.426 13.264 15.486 14.161 ;
      RECT MASK 1 15.592 13.264 15.652 14.161 ;
      RECT MASK 1 15.758 13.264 15.818 14.161 ;
      RECT MASK 1 16.256 13.264 16.316 14.336 ;
      RECT MASK 1 16.588 13.264 16.648 14.336 ;
      RECT MASK 1 17.086 13.264 17.146 14.161 ;
      RECT MASK 1 17.252 13.264 17.312 14.161 ;
      RECT MASK 1 17.418 13.264 17.478 14.161 ;
      RECT MASK 1 17.916 13.264 17.976 14.336 ;
      RECT MASK 1 18.248 13.264 18.308 14.336 ;
      RECT MASK 1 18.746 13.264 18.806 14.161 ;
      RECT MASK 1 19.078 13.264 19.138 14.161 ;
      RECT MASK 1 19.576 13.264 19.636 14.336 ;
      RECT MASK 1 19.742 13.264 19.802 14.161 ;
      RECT MASK 1 19.908 13.264 19.968 14.336 ;
      RECT MASK 1 20.406 13.264 20.466 14.161 ;
      RECT MASK 1 20.572 13.264 20.632 14.161 ;
      RECT MASK 1 20.738 13.264 20.798 14.161 ;
      RECT MASK 1 21.236 13.264 21.296 14.336 ;
      RECT MASK 1 21.402 13.264 21.462 14.161 ;
      RECT MASK 1 21.568 13.264 21.628 14.336 ;
      RECT MASK 1 22.066 13.264 22.126 14.161 ;
      RECT MASK 1 22.896 13.264 22.956 14.336 ;
      RECT MASK 1 23.228 13.264 23.288 14.336 ;
      RECT MASK 1 24.556 13.264 24.616 14.336 ;
      RECT MASK 1 24.888 13.264 24.948 14.336 ;
      RECT MASK 1 26.216 13.264 26.276 14.336 ;
      RECT MASK 1 26.548 13.264 26.608 14.336 ;
      RECT MASK 1 27.378 13.264 27.438 13.458 ;
      RECT MASK 1 28.208 13.264 28.268 14.336 ;
      RECT MASK 1 29.536 13.264 29.596 14.336 ;
      RECT MASK 1 30.2 13.264 30.26 14.161 ;
      RECT MASK 1 31.196 13.264 31.256 14.336 ;
      RECT MASK 1 31.528 13.264 31.588 14.336 ;
      RECT MASK 1 32.856 13.264 32.916 14.336 ;
      RECT MASK 1 33.188 13.264 33.248 14.336 ;
      RECT MASK 1 34.018 13.264 34.078 13.458 ;
      RECT MASK 1 35.346 13.264 35.406 13.458 ;
      RECT MASK 1 36.176 13.264 36.236 14.336 ;
      RECT MASK 1 36.508 13.264 36.568 14.336 ;
      RECT MASK 1 37.836 13.264 37.896 14.336 ;
      RECT MASK 1 38.168 13.264 38.228 14.336 ;
      RECT MASK 1 39.496 13.264 39.556 14.336 ;
      RECT MASK 1 39.828 13.264 39.888 14.336 ;
      RECT MASK 1 40.658 13.264 40.718 13.458 ;
      RECT MASK 1 41.488 13.264 41.548 14.336 ;
      RECT MASK 1 42.816 13.264 42.876 14.336 ;
      RECT MASK 1 43.148 13.264 43.208 14.336 ;
      RECT MASK 1 44.476 13.264 44.536 14.336 ;
      RECT MASK 1 44.808 13.264 44.868 14.336 ;
      RECT MASK 1 45.638 13.264 45.698 13.458 ;
      RECT MASK 1 46.468 13.264 46.528 14.336 ;
      RECT MASK 1 47.796 13.264 47.856 14.336 ;
      RECT MASK 1 48.128 13.264 48.188 14.336 ;
      RECT MASK 1 49.456 13.264 49.516 14.336 ;
      RECT MASK 1 49.788 13.264 49.848 14.336 ;
      RECT MASK 1 51.116 13.264 51.176 14.336 ;
      RECT MASK 1 51.448 13.264 51.508 14.336 ;
      RECT MASK 1 52.776 13.264 52.836 14.336 ;
      RECT MASK 1 53.108 13.264 53.168 14.336 ;
      RECT MASK 1 54.436 13.264 54.496 14.336 ;
      RECT MASK 1 54.768 13.264 54.828 14.336 ;
      RECT MASK 1 55.764 13.264 55.824 13.458 ;
      RECT MASK 1 56.096 13.264 56.156 14.336 ;
      RECT MASK 1 56.262 13.264 56.322 14.161 ;
      RECT MASK 1 56.428 13.264 56.488 14.161 ;
      RECT MASK 1 56.594 13.264 56.654 14.336 ;
      RECT MASK 1 57.922 13.264 57.982 14.336 ;
      RECT MASK 1 58.254 13.264 58.314 14.336 ;
      RECT MASK 1 59.582 13.264 59.642 14.336 ;
      RECT MASK 1 60.246 13.264 60.306 13.458 ;
      RECT MASK 1 61.242 13.264 61.302 14.336 ;
      RECT MASK 1 61.574 13.264 61.634 14.336 ;
      RECT MASK 1 62.404 13.264 62.464 13.458 ;
      RECT MASK 1 63.234 13.264 63.294 14.336 ;
      RECT MASK 1 64.562 13.264 64.622 14.336 ;
      RECT MASK 1 64.894 13.264 64.954 14.336 ;
      RECT MASK 1 66.222 13.264 66.282 14.336 ;
      RECT MASK 1 66.554 13.264 66.614 14.336 ;
      RECT MASK 1 67.882 13.264 67.942 14.336 ;
      RECT MASK 1 68.214 13.264 68.274 14.336 ;
      RECT MASK 1 69.542 13.264 69.602 14.336 ;
      RECT MASK 1 69.874 13.264 69.934 14.336 ;
      RECT MASK 1 71.202 13.264 71.262 14.336 ;
      RECT MASK 1 71.534 13.264 71.594 14.336 ;
      RECT MASK 1 72.862 13.264 72.922 14.336 ;
      RECT MASK 1 73.692 13.264 73.752 14.161 ;
      RECT MASK 1 73.858 13.264 73.918 14.161 ;
      RECT MASK 1 74.024 13.264 74.084 14.161 ;
      RECT MASK 1 74.522 13.264 74.582 14.336 ;
      RECT MASK 1 74.688 13.264 74.748 14.161 ;
      RECT MASK 1 74.854 13.264 74.914 14.336 ;
      RECT MASK 1 75.352 13.264 75.412 14.161 ;
      RECT MASK 1 75.518 13.264 75.578 14.161 ;
      RECT MASK 1 75.684 13.264 75.744 14.161 ;
      RECT MASK 1 76.182 13.264 76.242 14.336 ;
      RECT MASK 1 76.514 13.264 76.574 14.336 ;
      RECT MASK 1 77.012 13.264 77.072 14.161 ;
      RECT MASK 1 77.178 13.264 77.238 14.161 ;
      RECT MASK 1 77.842 13.264 77.902 14.336 ;
      RECT MASK 1 78.174 13.264 78.234 14.336 ;
      RECT MASK 1 79.502 13.264 79.562 14.336 ;
      RECT MASK 1 79.834 13.264 79.894 14.336 ;
      RECT MASK 1 80.664 13.264 80.724 14.161 ;
      RECT MASK 1 81.162 13.264 81.222 14.336 ;
      RECT MASK 1 81.328 13.264 81.388 14.161 ;
      RECT MASK 1 81.494 13.264 81.554 14.336 ;
      RECT MASK 1 81.992 13.264 82.052 14.161 ;
      RECT MASK 1 82.158 13.264 82.218 14.161 ;
      RECT MASK 1 82.324 13.264 82.384 14.161 ;
      RECT MASK 1 82.822 13.264 82.882 14.336 ;
      RECT MASK 1 82.988 13.264 83.048 14.161 ;
      RECT MASK 1 83.154 13.264 83.214 14.336 ;
      RECT MASK 1 84.482 13.264 84.542 14.336 ;
      RECT MASK 1 84.814 13.264 84.874 14.336 ;
      RECT MASK 1 85.312 13.264 85.372 14.161 ;
      RECT MASK 1 85.478 13.264 85.538 14.161 ;
      RECT MASK 1 85.644 13.264 85.704 14.161 ;
      RECT MASK 1 86.142 13.264 86.202 14.336 ;
      RECT MASK 1 86.308 13.264 86.368 14.161 ;
      RECT MASK 1 86.474 13.264 86.534 14.336 ;
      RECT MASK 1 86.972 13.264 87.032 14.161 ;
      RECT MASK 1 87.138 13.264 87.198 14.161 ;
      RECT MASK 1 87.304 13.264 87.364 14.161 ;
      RECT MASK 1 87.802 13.264 87.862 14.336 ;
      RECT MASK 1 87.968 13.264 88.028 14.161 ;
      RECT MASK 1 88.134 13.264 88.194 14.336 ;
      RECT MASK 1 88.632 13.264 88.692 14.161 ;
      RECT MASK 1 88.798 13.264 88.858 14.161 ;
      RECT MASK 1 89.462 13.264 89.522 14.336 ;
      RECT MASK 1 89.794 13.264 89.854 14.336 ;
      RECT MASK 1 91.122 13.264 91.182 14.336 ;
      RECT MASK 1 91.454 13.264 91.514 14.336 ;
      RECT MASK 1 92.118 13.264 92.178 14.161 ;
      RECT MASK 1 92.284 13.264 92.344 14.161 ;
      RECT MASK 1 92.782 13.264 92.842 14.336 ;
      RECT MASK 1 92.948 13.264 93.008 14.161 ;
      RECT MASK 1 93.114 13.264 93.174 14.336 ;
      RECT MASK 1 93.612 13.264 93.672 14.161 ;
      RECT MASK 1 93.778 13.264 93.838 14.161 ;
      RECT MASK 1 93.944 13.264 94.004 14.161 ;
      RECT MASK 1 94.442 13.264 94.502 14.336 ;
      RECT MASK 1 94.774 13.264 94.834 14.336 ;
      RECT MASK 1 95.272 13.264 95.332 14.161 ;
      RECT MASK 1 95.438 13.264 95.498 14.161 ;
      RECT MASK 1 95.604 13.264 95.664 14.161 ;
      RECT MASK 1 96.102 13.264 96.162 14.336 ;
      RECT MASK 1 96.434 13.264 96.494 14.336 ;
      RECT MASK 1 96.932 13.264 96.992 14.161 ;
      RECT MASK 1 97.098 13.264 97.158 14.161 ;
      RECT MASK 1 97.264 13.264 97.324 14.161 ;
      RECT MASK 1 97.762 13.264 97.822 14.336 ;
      RECT MASK 1 98.094 13.264 98.154 14.336 ;
      RECT MASK 1 98.592 13.264 98.652 14.161 ;
      RECT MASK 1 98.758 13.264 98.818 14.161 ;
      RECT MASK 1 98.924 13.264 98.984 14.161 ;
      RECT MASK 1 99.422 13.264 99.482 14.336 ;
      RECT MASK 1 99.588 13.264 99.648 14.161 ;
      RECT MASK 1 99.754 13.264 99.814 14.336 ;
      RECT MASK 1 100.252 13.264 100.312 14.161 ;
      RECT MASK 1 100.418 13.264 100.478 14.161 ;
      RECT MASK 1 100.584 13.264 100.644 14.161 ;
      RECT MASK 1 101.082 13.264 101.142 14.336 ;
      RECT MASK 1 101.248 13.264 101.308 14.161 ;
      RECT MASK 1 101.414 13.264 101.474 14.336 ;
      RECT MASK 1 102.742 13.264 102.802 14.336 ;
      RECT MASK 1 103.074 13.264 103.134 14.336 ;
      RECT MASK 1 104.402 13.264 104.462 14.336 ;
      RECT MASK 1 104.734 13.264 104.794 14.336 ;
      RECT MASK 1 105.232 13.264 105.292 14.161 ;
      RECT MASK 1 105.398 13.264 105.458 14.161 ;
      RECT MASK 1 105.564 13.264 105.624 14.161 ;
      RECT MASK 1 106.062 13.264 106.122 14.336 ;
      RECT MASK 1 106.228 13.264 106.288 14.161 ;
      RECT MASK 1 106.394 13.264 106.454 14.336 ;
      RECT MASK 1 106.892 13.264 106.952 14.161 ;
      RECT MASK 1 107.058 13.264 107.118 14.161 ;
      RECT MASK 1 107.224 13.264 107.284 14.161 ;
      RECT MASK 1 107.722 13.264 107.782 14.336 ;
      RECT MASK 1 108.054 13.264 108.114 14.336 ;
      RECT MASK 1 108.552 13.264 108.612 14.161 ;
      RECT MASK 1 108.718 13.264 108.778 14.161 ;
      RECT MASK 1 108.884 13.264 108.944 14.161 ;
      RECT MASK 1 109.382 13.264 109.442 14.336 ;
      RECT MASK 1 109.548 13.264 109.608 14.161 ;
      RECT MASK 1 109.714 13.264 109.774 14.336 ;
      RECT MASK 1 110.212 13.264 110.272 14.161 ;
      RECT MASK 1 110.544 13.264 110.604 14.161 ;
      RECT MASK 1 111.042 13.264 111.102 14.336 ;
      RECT MASK 1 111.208 13.264 111.268 14.161 ;
      RECT MASK 1 111.374 13.264 111.434 14.161 ;
      RECT MASK 1 8.786 13.439 8.846 14.161 ;
      RECT MASK 1 9.118 13.439 9.178 14.161 ;
      RECT MASK 1 9.782 13.439 9.842 14.161 ;
      RECT MASK 1 10.446 13.439 10.506 14.161 ;
      RECT MASK 1 10.778 13.439 10.838 14.161 ;
      RECT MASK 1 11.442 13.439 11.502 14.161 ;
      RECT MASK 1 22.232 13.439 22.292 14.161 ;
      RECT MASK 1 22.398 13.439 22.458 14.161 ;
      RECT MASK 1 23.726 13.439 23.786 14.161 ;
      RECT MASK 1 23.892 13.439 23.952 14.161 ;
      RECT MASK 1 24.058 13.439 24.118 14.161 ;
      RECT MASK 1 25.386 13.439 25.446 14.161 ;
      RECT MASK 1 25.552 13.439 25.612 14.161 ;
      RECT MASK 1 25.718 13.439 25.778 14.161 ;
      RECT MASK 1 27.046 13.439 27.106 14.161 ;
      RECT MASK 1 27.212 13.439 27.272 14.161 ;
      RECT MASK 1 27.876 13.439 27.936 14.336 ;
      RECT MASK 1 28.706 13.439 28.766 14.161 ;
      RECT MASK 1 28.872 13.439 28.932 14.161 ;
      RECT MASK 1 29.038 13.439 29.098 14.161 ;
      RECT MASK 1 29.868 13.439 29.928 14.336 ;
      RECT MASK 1 30.366 13.439 30.426 14.161 ;
      RECT MASK 1 30.532 13.439 30.592 14.161 ;
      RECT MASK 1 30.698 13.439 30.758 14.161 ;
      RECT MASK 1 32.026 13.439 32.086 14.161 ;
      RECT MASK 1 32.192 13.439 32.252 14.161 ;
      RECT MASK 1 32.358 13.439 32.418 14.161 ;
      RECT MASK 1 33.022 13.439 33.082 14.161 ;
      RECT MASK 1 33.686 13.439 33.746 14.161 ;
      RECT MASK 1 34.516 13.439 34.576 14.336 ;
      RECT MASK 1 34.848 13.439 34.908 14.336 ;
      RECT MASK 1 35.512 13.439 35.572 14.161 ;
      RECT MASK 1 35.678 13.439 35.738 14.161 ;
      RECT MASK 1 36.342 13.439 36.402 14.161 ;
      RECT MASK 1 37.006 13.439 37.066 14.161 ;
      RECT MASK 1 37.172 13.439 37.232 14.161 ;
      RECT MASK 1 37.338 13.439 37.398 14.161 ;
      RECT MASK 1 38.666 13.439 38.726 14.161 ;
      RECT MASK 1 38.832 13.439 38.892 14.161 ;
      RECT MASK 1 38.998 13.439 39.058 14.161 ;
      RECT MASK 1 39.662 13.439 39.722 14.161 ;
      RECT MASK 1 40.326 13.439 40.386 14.161 ;
      RECT MASK 1 40.492 13.439 40.552 14.161 ;
      RECT MASK 1 41.156 13.439 41.216 14.336 ;
      RECT MASK 1 41.986 13.439 42.046 14.161 ;
      RECT MASK 1 42.318 13.439 42.378 14.161 ;
      RECT MASK 1 43.646 13.439 43.706 14.161 ;
      RECT MASK 1 43.812 13.439 43.872 14.161 ;
      RECT MASK 1 43.978 13.439 44.038 14.161 ;
      RECT MASK 1 45.306 13.439 45.366 14.161 ;
      RECT MASK 1 46.136 13.439 46.196 14.336 ;
      RECT MASK 1 46.966 13.439 47.026 14.161 ;
      RECT MASK 1 47.132 13.439 47.192 14.161 ;
      RECT MASK 1 47.298 13.439 47.358 14.161 ;
      RECT MASK 1 48.626 13.439 48.686 14.161 ;
      RECT MASK 1 48.792 13.439 48.852 14.161 ;
      RECT MASK 1 48.958 13.439 49.018 14.161 ;
      RECT MASK 1 50.286 13.439 50.346 14.161 ;
      RECT MASK 1 50.452 13.439 50.512 14.161 ;
      RECT MASK 1 50.618 13.439 50.678 14.161 ;
      RECT MASK 1 51.946 13.439 52.006 14.161 ;
      RECT MASK 1 52.112 13.439 52.172 14.161 ;
      RECT MASK 1 52.278 13.439 52.338 14.161 ;
      RECT MASK 1 52.942 13.439 53.002 14.161 ;
      RECT MASK 1 53.606 13.439 53.666 14.161 ;
      RECT MASK 1 53.772 13.439 53.832 14.161 ;
      RECT MASK 1 53.938 13.439 53.998 14.161 ;
      RECT MASK 1 54.602 13.439 54.662 14.161 ;
      RECT MASK 1 55.266 13.439 55.326 14.161 ;
      RECT MASK 1 55.432 13.439 55.492 14.161 ;
      RECT MASK 1 55.598 13.439 55.658 14.161 ;
      RECT MASK 1 57.092 13.439 57.152 14.161 ;
      RECT MASK 1 57.424 13.439 57.484 14.161 ;
      RECT MASK 1 58.752 13.439 58.812 14.161 ;
      RECT MASK 1 58.918 13.439 58.978 14.161 ;
      RECT MASK 1 59.084 13.439 59.144 14.161 ;
      RECT MASK 1 59.748 13.439 59.808 14.161 ;
      RECT MASK 1 59.914 13.439 59.974 14.336 ;
      RECT MASK 1 60.412 13.439 60.472 14.161 ;
      RECT MASK 1 60.744 13.439 60.804 14.161 ;
      RECT MASK 1 62.072 13.439 62.132 14.161 ;
      RECT MASK 1 62.238 13.439 62.298 14.161 ;
      RECT MASK 1 62.902 13.439 62.962 14.336 ;
      RECT MASK 1 63.732 13.439 63.792 14.161 ;
      RECT MASK 1 63.898 13.439 63.958 14.161 ;
      RECT MASK 1 64.064 13.439 64.124 14.161 ;
      RECT MASK 1 65.392 13.439 65.452 14.161 ;
      RECT MASK 1 65.724 13.439 65.784 14.161 ;
      RECT MASK 1 66.388 13.439 66.448 14.161 ;
      RECT MASK 1 67.052 13.439 67.112 14.161 ;
      RECT MASK 1 67.384 13.439 67.444 14.161 ;
      RECT MASK 1 68.712 13.439 68.772 14.161 ;
      RECT MASK 1 68.878 13.439 68.938 14.161 ;
      RECT MASK 1 69.044 13.439 69.104 14.161 ;
      RECT MASK 1 70.372 13.439 70.432 14.161 ;
      RECT MASK 1 70.704 13.439 70.764 14.161 ;
      RECT MASK 1 71.368 13.439 71.428 14.161 ;
      RECT MASK 1 72.032 13.439 72.092 14.161 ;
      RECT MASK 1 72.364 13.439 72.424 14.161 ;
      RECT MASK 1 73.194 13.439 73.254 14.336 ;
      RECT MASK 1 77.344 13.439 77.404 14.161 ;
      RECT MASK 1 78.008 13.439 78.068 14.161 ;
      RECT MASK 1 78.672 13.439 78.732 14.161 ;
      RECT MASK 1 78.838 13.439 78.898 14.161 ;
      RECT MASK 1 79.004 13.439 79.064 14.161 ;
      RECT MASK 1 80.332 13.439 80.392 14.161 ;
      RECT MASK 1 80.498 13.439 80.558 14.161 ;
      RECT MASK 1 83.652 13.439 83.712 14.161 ;
      RECT MASK 1 83.818 13.439 83.878 14.161 ;
      RECT MASK 1 83.984 13.439 84.044 14.161 ;
      RECT MASK 1 88.964 13.439 89.024 14.161 ;
      RECT MASK 1 90.292 13.439 90.352 14.161 ;
      RECT MASK 1 90.458 13.439 90.518 14.161 ;
      RECT MASK 1 90.624 13.439 90.684 14.161 ;
      RECT MASK 1 91.952 13.439 92.012 14.161 ;
      RECT MASK 1 101.912 13.439 101.972 14.161 ;
      RECT MASK 1 102.244 13.439 102.304 14.161 ;
      RECT MASK 1 102.908 13.439 102.968 14.161 ;
      RECT MASK 1 103.572 13.439 103.632 14.161 ;
      RECT MASK 1 103.738 13.439 103.798 14.161 ;
      RECT MASK 1 103.904 13.439 103.964 14.161 ;
      RECT MASK 1 4.968 14.456 5.028 15.064 ;
      RECT MASK 1 5.3 14.456 5.36 15.064 ;
      RECT MASK 1 5.964 14.456 6.024 15.064 ;
      RECT MASK 1 6.296 14.456 6.356 15.064 ;
      RECT MASK 1 6.628 14.456 6.688 15.064 ;
      RECT MASK 1 6.96 14.456 7.02 15.064 ;
      RECT MASK 1 7.624 14.456 7.684 15.064 ;
      RECT MASK 1 7.956 14.456 8.016 15.064 ;
      RECT MASK 1 8.288 14.456 8.348 15.064 ;
      RECT MASK 1 8.62 14.456 8.68 15.064 ;
      RECT MASK 1 9.284 14.456 9.344 15.064 ;
      RECT MASK 1 9.616 14.456 9.676 15.064 ;
      RECT MASK 1 9.948 14.456 10.008 15.064 ;
      RECT MASK 1 10.28 14.456 10.34 15.064 ;
      RECT MASK 1 10.944 14.456 11.004 15.064 ;
      RECT MASK 1 11.276 14.456 11.336 15.064 ;
      RECT MASK 1 11.608 14.456 11.668 15.064 ;
      RECT MASK 1 11.94 14.456 12 15.064 ;
      RECT MASK 1 12.604 14.456 12.664 15.064 ;
      RECT MASK 1 12.936 14.456 12.996 15.064 ;
      RECT MASK 1 13.268 14.456 13.328 15.064 ;
      RECT MASK 1 13.6 14.456 13.66 15.064 ;
      RECT MASK 1 14.264 14.456 14.324 15.064 ;
      RECT MASK 1 14.596 14.456 14.656 15.064 ;
      RECT MASK 1 14.928 14.456 14.988 15.064 ;
      RECT MASK 1 15.26 14.456 15.32 15.064 ;
      RECT MASK 1 15.924 14.456 15.984 15.064 ;
      RECT MASK 1 16.256 14.456 16.316 15.064 ;
      RECT MASK 1 16.588 14.456 16.648 15.064 ;
      RECT MASK 1 16.92 14.456 16.98 15.064 ;
      RECT MASK 1 17.584 14.456 17.644 15.064 ;
      RECT MASK 1 17.916 14.456 17.976 15.064 ;
      RECT MASK 1 18.248 14.456 18.308 15.064 ;
      RECT MASK 1 18.58 14.456 18.64 15.064 ;
      RECT MASK 1 19.244 14.456 19.304 15.064 ;
      RECT MASK 1 19.576 14.456 19.636 15.064 ;
      RECT MASK 1 19.908 14.456 19.968 15.064 ;
      RECT MASK 1 20.24 14.456 20.3 15.064 ;
      RECT MASK 1 20.904 14.456 20.964 15.064 ;
      RECT MASK 1 21.236 14.456 21.296 15.064 ;
      RECT MASK 1 21.568 14.456 21.628 15.064 ;
      RECT MASK 1 21.9 14.456 21.96 15.064 ;
      RECT MASK 1 22.564 14.456 22.624 15.064 ;
      RECT MASK 1 22.896 14.456 22.956 15.064 ;
      RECT MASK 1 23.228 14.456 23.288 15.064 ;
      RECT MASK 1 23.56 14.456 23.62 15.064 ;
      RECT MASK 1 24.224 14.456 24.284 15.064 ;
      RECT MASK 1 24.556 14.456 24.616 15.064 ;
      RECT MASK 1 24.888 14.456 24.948 15.064 ;
      RECT MASK 1 25.22 14.456 25.28 15.064 ;
      RECT MASK 1 25.884 14.456 25.944 15.064 ;
      RECT MASK 1 26.216 14.456 26.276 15.064 ;
      RECT MASK 1 26.548 14.456 26.608 15.064 ;
      RECT MASK 1 26.88 14.456 26.94 15.064 ;
      RECT MASK 1 27.544 14.456 27.604 15.064 ;
      RECT MASK 1 27.876 14.456 27.936 15.064 ;
      RECT MASK 1 28.208 14.456 28.268 15.064 ;
      RECT MASK 1 28.54 14.456 28.6 15.064 ;
      RECT MASK 1 29.204 14.456 29.264 15.064 ;
      RECT MASK 1 29.536 14.456 29.596 15.064 ;
      RECT MASK 1 29.868 14.456 29.928 15.064 ;
      RECT MASK 1 30.2 14.456 30.26 15.064 ;
      RECT MASK 1 30.864 14.456 30.924 15.064 ;
      RECT MASK 1 31.196 14.456 31.256 15.064 ;
      RECT MASK 1 31.528 14.456 31.588 15.064 ;
      RECT MASK 1 31.86 14.456 31.92 15.064 ;
      RECT MASK 1 32.524 14.456 32.584 15.064 ;
      RECT MASK 1 32.856 14.456 32.916 15.064 ;
      RECT MASK 1 33.188 14.456 33.248 15.064 ;
      RECT MASK 1 33.52 14.456 33.58 15.064 ;
      RECT MASK 1 34.184 14.456 34.244 15.064 ;
      RECT MASK 1 34.516 14.456 34.576 15.064 ;
      RECT MASK 1 34.848 14.456 34.908 15.064 ;
      RECT MASK 1 35.18 14.456 35.24 15.064 ;
      RECT MASK 1 35.844 14.456 35.904 15.064 ;
      RECT MASK 1 36.176 14.456 36.236 15.064 ;
      RECT MASK 1 36.508 14.456 36.568 15.064 ;
      RECT MASK 1 36.84 14.456 36.9 15.064 ;
      RECT MASK 1 37.504 14.456 37.564 15.064 ;
      RECT MASK 1 37.836 14.456 37.896 15.064 ;
      RECT MASK 1 38.168 14.456 38.228 15.064 ;
      RECT MASK 1 38.5 14.456 38.56 15.064 ;
      RECT MASK 1 39.164 14.456 39.224 15.064 ;
      RECT MASK 1 39.496 14.456 39.556 15.064 ;
      RECT MASK 1 39.828 14.456 39.888 15.064 ;
      RECT MASK 1 40.16 14.456 40.22 15.064 ;
      RECT MASK 1 40.824 14.456 40.884 15.064 ;
      RECT MASK 1 41.156 14.456 41.216 15.064 ;
      RECT MASK 1 41.488 14.456 41.548 15.064 ;
      RECT MASK 1 41.82 14.456 41.88 15.064 ;
      RECT MASK 1 42.484 14.456 42.544 15.064 ;
      RECT MASK 1 42.816 14.456 42.876 15.064 ;
      RECT MASK 1 43.148 14.456 43.208 15.064 ;
      RECT MASK 1 43.48 14.456 43.54 15.064 ;
      RECT MASK 1 44.144 14.456 44.204 15.064 ;
      RECT MASK 1 44.476 14.456 44.536 15.064 ;
      RECT MASK 1 44.808 14.456 44.868 15.064 ;
      RECT MASK 1 45.14 14.456 45.2 15.064 ;
      RECT MASK 1 45.804 14.456 45.864 15.064 ;
      RECT MASK 1 46.136 14.456 46.196 15.064 ;
      RECT MASK 1 46.468 14.456 46.528 15.064 ;
      RECT MASK 1 46.8 14.456 46.86 15.064 ;
      RECT MASK 1 47.464 14.456 47.524 15.064 ;
      RECT MASK 1 47.796 14.456 47.856 15.064 ;
      RECT MASK 1 48.128 14.456 48.188 15.064 ;
      RECT MASK 1 48.46 14.456 48.52 15.064 ;
      RECT MASK 1 49.124 14.456 49.184 15.064 ;
      RECT MASK 1 49.456 14.456 49.516 15.064 ;
      RECT MASK 1 49.788 14.456 49.848 15.064 ;
      RECT MASK 1 50.12 14.456 50.18 15.064 ;
      RECT MASK 1 50.784 14.456 50.844 15.064 ;
      RECT MASK 1 51.116 14.456 51.176 15.064 ;
      RECT MASK 1 51.448 14.456 51.508 15.064 ;
      RECT MASK 1 51.78 14.456 51.84 15.064 ;
      RECT MASK 1 52.444 14.456 52.504 15.064 ;
      RECT MASK 1 52.776 14.456 52.836 15.064 ;
      RECT MASK 1 53.108 14.456 53.168 15.064 ;
      RECT MASK 1 53.44 14.456 53.5 15.064 ;
      RECT MASK 1 54.104 14.456 54.164 15.064 ;
      RECT MASK 1 54.436 14.456 54.496 15.064 ;
      RECT MASK 1 54.768 14.456 54.828 15.064 ;
      RECT MASK 1 55.1 14.456 55.16 15.064 ;
      RECT MASK 1 55.764 14.456 55.824 15.064 ;
      RECT MASK 1 56.096 14.456 56.156 15.064 ;
      RECT MASK 1 56.594 14.456 56.654 15.064 ;
      RECT MASK 1 56.926 14.456 56.986 15.064 ;
      RECT MASK 1 57.59 14.456 57.65 15.064 ;
      RECT MASK 1 57.922 14.456 57.982 15.064 ;
      RECT MASK 1 58.254 14.456 58.314 15.064 ;
      RECT MASK 1 58.586 14.456 58.646 15.064 ;
      RECT MASK 1 59.25 14.456 59.31 15.064 ;
      RECT MASK 1 59.582 14.456 59.642 15.064 ;
      RECT MASK 1 59.914 14.456 59.974 15.064 ;
      RECT MASK 1 60.246 14.456 60.306 15.064 ;
      RECT MASK 1 60.91 14.456 60.97 15.064 ;
      RECT MASK 1 61.242 14.456 61.302 15.064 ;
      RECT MASK 1 61.574 14.456 61.634 15.064 ;
      RECT MASK 1 61.906 14.456 61.966 15.064 ;
      RECT MASK 1 62.57 14.456 62.63 15.064 ;
      RECT MASK 1 62.902 14.456 62.962 15.064 ;
      RECT MASK 1 63.234 14.456 63.294 15.064 ;
      RECT MASK 1 63.566 14.456 63.626 15.064 ;
      RECT MASK 1 64.23 14.456 64.29 15.064 ;
      RECT MASK 1 64.562 14.456 64.622 15.064 ;
      RECT MASK 1 64.894 14.456 64.954 15.064 ;
      RECT MASK 1 65.226 14.456 65.286 15.064 ;
      RECT MASK 1 65.89 14.456 65.95 15.064 ;
      RECT MASK 1 66.222 14.456 66.282 15.064 ;
      RECT MASK 1 66.554 14.456 66.614 15.064 ;
      RECT MASK 1 66.886 14.456 66.946 15.064 ;
      RECT MASK 1 67.55 14.456 67.61 15.064 ;
      RECT MASK 1 67.882 14.456 67.942 15.064 ;
      RECT MASK 1 68.214 14.456 68.274 15.064 ;
      RECT MASK 1 68.546 14.456 68.606 15.064 ;
      RECT MASK 1 69.21 14.456 69.27 15.064 ;
      RECT MASK 1 69.542 14.456 69.602 15.064 ;
      RECT MASK 1 69.874 14.456 69.934 15.064 ;
      RECT MASK 1 70.206 14.456 70.266 15.064 ;
      RECT MASK 1 70.87 14.456 70.93 15.064 ;
      RECT MASK 1 71.202 14.456 71.262 15.064 ;
      RECT MASK 1 71.534 14.456 71.594 15.064 ;
      RECT MASK 1 71.866 14.456 71.926 15.064 ;
      RECT MASK 1 72.53 14.456 72.59 15.064 ;
      RECT MASK 1 72.862 14.456 72.922 15.064 ;
      RECT MASK 1 73.194 14.456 73.254 15.064 ;
      RECT MASK 1 73.526 14.456 73.586 15.064 ;
      RECT MASK 1 74.19 14.456 74.25 15.064 ;
      RECT MASK 1 74.522 14.456 74.582 15.064 ;
      RECT MASK 1 74.854 14.456 74.914 15.064 ;
      RECT MASK 1 75.186 14.456 75.246 15.064 ;
      RECT MASK 1 75.85 14.456 75.91 15.064 ;
      RECT MASK 1 76.182 14.456 76.242 15.064 ;
      RECT MASK 1 76.514 14.456 76.574 15.064 ;
      RECT MASK 1 76.846 14.456 76.906 15.064 ;
      RECT MASK 1 77.51 14.456 77.57 15.064 ;
      RECT MASK 1 77.842 14.456 77.902 15.064 ;
      RECT MASK 1 78.174 14.456 78.234 15.064 ;
      RECT MASK 1 78.506 14.456 78.566 15.064 ;
      RECT MASK 1 79.17 14.456 79.23 15.064 ;
      RECT MASK 1 79.502 14.456 79.562 15.064 ;
      RECT MASK 1 79.834 14.456 79.894 15.064 ;
      RECT MASK 1 80.166 14.456 80.226 15.064 ;
      RECT MASK 1 80.83 14.456 80.89 15.064 ;
      RECT MASK 1 81.162 14.456 81.222 15.064 ;
      RECT MASK 1 81.494 14.456 81.554 15.064 ;
      RECT MASK 1 81.826 14.456 81.886 15.064 ;
      RECT MASK 1 82.49 14.456 82.55 15.064 ;
      RECT MASK 1 82.822 14.456 82.882 15.064 ;
      RECT MASK 1 83.154 14.456 83.214 15.064 ;
      RECT MASK 1 83.486 14.456 83.546 15.064 ;
      RECT MASK 1 84.15 14.456 84.21 15.064 ;
      RECT MASK 1 84.482 14.456 84.542 15.064 ;
      RECT MASK 1 84.814 14.456 84.874 15.064 ;
      RECT MASK 1 85.146 14.456 85.206 15.064 ;
      RECT MASK 1 85.81 14.456 85.87 15.064 ;
      RECT MASK 1 86.142 14.456 86.202 15.064 ;
      RECT MASK 1 86.474 14.456 86.534 15.064 ;
      RECT MASK 1 86.806 14.456 86.866 15.064 ;
      RECT MASK 1 87.47 14.456 87.53 15.064 ;
      RECT MASK 1 87.802 14.456 87.862 15.064 ;
      RECT MASK 1 88.134 14.456 88.194 15.064 ;
      RECT MASK 1 88.466 14.456 88.526 15.064 ;
      RECT MASK 1 89.13 14.456 89.19 15.064 ;
      RECT MASK 1 89.462 14.456 89.522 15.064 ;
      RECT MASK 1 89.794 14.456 89.854 15.064 ;
      RECT MASK 1 90.126 14.456 90.186 15.064 ;
      RECT MASK 1 90.79 14.456 90.85 15.064 ;
      RECT MASK 1 91.122 14.456 91.182 15.064 ;
      RECT MASK 1 91.454 14.456 91.514 15.064 ;
      RECT MASK 1 91.786 14.456 91.846 15.064 ;
      RECT MASK 1 92.45 14.456 92.51 15.064 ;
      RECT MASK 1 92.782 14.456 92.842 15.064 ;
      RECT MASK 1 93.114 14.456 93.174 15.064 ;
      RECT MASK 1 93.446 14.456 93.506 15.064 ;
      RECT MASK 1 94.11 14.456 94.17 15.064 ;
      RECT MASK 1 94.442 14.456 94.502 15.064 ;
      RECT MASK 1 94.774 14.456 94.834 15.064 ;
      RECT MASK 1 95.106 14.456 95.166 15.064 ;
      RECT MASK 1 95.77 14.456 95.83 15.064 ;
      RECT MASK 1 96.102 14.456 96.162 15.064 ;
      RECT MASK 1 96.434 14.456 96.494 15.064 ;
      RECT MASK 1 96.766 14.456 96.826 15.064 ;
      RECT MASK 1 97.43 14.456 97.49 15.064 ;
      RECT MASK 1 97.762 14.456 97.822 15.064 ;
      RECT MASK 1 98.094 14.456 98.154 15.064 ;
      RECT MASK 1 98.426 14.456 98.486 15.064 ;
      RECT MASK 1 99.09 14.456 99.15 15.064 ;
      RECT MASK 1 99.422 14.456 99.482 15.064 ;
      RECT MASK 1 99.754 14.456 99.814 15.064 ;
      RECT MASK 1 100.086 14.456 100.146 15.064 ;
      RECT MASK 1 100.75 14.456 100.81 15.064 ;
      RECT MASK 1 101.082 14.456 101.142 15.064 ;
      RECT MASK 1 101.414 14.456 101.474 15.064 ;
      RECT MASK 1 101.746 14.456 101.806 15.064 ;
      RECT MASK 1 102.41 14.456 102.47 15.064 ;
      RECT MASK 1 102.742 14.456 102.802 15.064 ;
      RECT MASK 1 103.074 14.456 103.134 15.064 ;
      RECT MASK 1 103.406 14.456 103.466 15.064 ;
      RECT MASK 1 104.07 14.456 104.13 15.064 ;
      RECT MASK 1 104.402 14.456 104.462 15.064 ;
      RECT MASK 1 104.734 14.456 104.794 15.064 ;
      RECT MASK 1 105.066 14.456 105.126 15.064 ;
      RECT MASK 1 105.73 14.456 105.79 15.064 ;
      RECT MASK 1 106.062 14.456 106.122 15.064 ;
      RECT MASK 1 106.394 14.456 106.454 15.064 ;
      RECT MASK 1 106.726 14.456 106.786 15.064 ;
      RECT MASK 1 107.39 14.456 107.45 15.064 ;
      RECT MASK 1 107.722 14.456 107.782 15.064 ;
      RECT MASK 1 108.054 14.456 108.114 15.064 ;
      RECT MASK 1 108.386 14.456 108.446 15.064 ;
      RECT MASK 1 109.05 14.456 109.11 15.064 ;
      RECT MASK 1 109.382 14.456 109.442 15.064 ;
      RECT MASK 1 109.714 14.456 109.774 15.064 ;
      RECT MASK 1 110.046 14.456 110.106 15.064 ;
      RECT MASK 1 110.71 14.456 110.77 15.064 ;
      RECT MASK 1 111.042 14.456 111.102 15.064 ;
      RECT MASK 1 52.112 14.487 52.172 16.765 ;
      RECT MASK 1 109.548 14.581 109.608 16.763 ;
      RECT MASK 1 13.932 14.773 13.992 16.763 ;
      RECT MASK 1 5.632 14.869 5.692 16.859 ;
      RECT MASK 1 54.602 14.869 54.662 16.763 ;
      RECT MASK 1 56.428 14.869 56.488 16.763 ;
      RECT MASK 1 58.918 14.869 58.978 16.763 ;
      RECT MASK 1 66.388 14.869 66.448 16.763 ;
      RECT MASK 1 17.252 14.961 17.312 16.953 ;
      RECT MASK 1 30.532 14.961 30.592 16.953 ;
      RECT MASK 1 43.812 14.961 43.872 16.953 ;
      RECT MASK 1 57.258 14.961 57.318 16.953 ;
      RECT MASK 1 70.538 14.961 70.598 16.953 ;
      RECT MASK 1 82.158 14.961 82.218 16.859 ;
      RECT MASK 1 83.818 14.961 83.878 16.953 ;
      RECT MASK 1 97.098 14.961 97.158 16.953 ;
      RECT MASK 1 108.718 14.961 108.778 16.859 ;
      RECT MASK 1 11.442 14.963 11.502 16.477 ;
      RECT MASK 1 12.272 14.963 12.332 16.571 ;
      RECT MASK 1 13.102 14.963 13.162 16.667 ;
      RECT MASK 1 15.592 14.963 15.652 16.859 ;
      RECT MASK 1 23.892 14.963 23.952 16.477 ;
      RECT MASK 1 25.552 14.963 25.612 16.571 ;
      RECT MASK 1 27.212 14.963 27.272 16.667 ;
      RECT MASK 1 28.872 14.963 28.932 16.859 ;
      RECT MASK 1 37.172 14.963 37.232 16.477 ;
      RECT MASK 1 38.832 14.963 38.892 16.571 ;
      RECT MASK 1 40.492 14.963 40.552 16.667 ;
      RECT MASK 1 42.152 14.963 42.212 16.859 ;
      RECT MASK 1 50.452 14.963 50.512 16.477 ;
      RECT MASK 1 51.282 14.963 51.342 16.477 ;
      RECT MASK 1 53.772 14.963 53.832 16.667 ;
      RECT MASK 1 55.432 14.963 55.492 16.859 ;
      RECT MASK 1 63.898 14.963 63.958 16.477 ;
      RECT MASK 1 65.558 14.963 65.618 16.571 ;
      RECT MASK 1 67.218 14.963 67.278 16.667 ;
      RECT MASK 1 68.878 14.963 68.938 16.859 ;
      RECT MASK 1 77.178 14.963 77.238 16.477 ;
      RECT MASK 1 78.838 14.963 78.898 16.571 ;
      RECT MASK 1 90.458 14.963 90.518 16.477 ;
      RECT MASK 1 92.118 14.963 92.178 16.571 ;
      RECT MASK 1 93.778 14.963 93.838 16.667 ;
      RECT MASK 1 95.438 14.963 95.498 16.859 ;
      RECT MASK 1 103.738 14.963 103.798 16.477 ;
      RECT MASK 1 105.398 14.963 105.458 16.571 ;
      RECT MASK 1 107.058 14.963 107.118 16.667 ;
      RECT MASK 1 110.378 14.963 110.438 16.953 ;
      RECT MASK 1 31.362 15.055 31.422 17.429 ;
      RECT MASK 1 71.368 15.055 71.428 17.429 ;
      RECT MASK 1 78.008 15.055 78.068 17.429 ;
      RECT MASK 1 4.636 15.184 4.696 16.256 ;
      RECT MASK 1 4.802 15.184 4.862 16.256 ;
      RECT MASK 1 4.968 15.184 5.028 16.256 ;
      RECT MASK 1 6.296 15.184 6.356 16.256 ;
      RECT MASK 1 6.628 15.184 6.688 16.256 ;
      RECT MASK 1 7.956 15.184 8.016 16.256 ;
      RECT MASK 1 8.288 15.184 8.348 16.256 ;
      RECT MASK 1 9.616 15.184 9.676 16.256 ;
      RECT MASK 1 9.948 15.184 10.008 16.256 ;
      RECT MASK 1 11.276 15.184 11.336 16.256 ;
      RECT MASK 1 11.608 15.184 11.668 16.256 ;
      RECT MASK 1 12.936 15.184 12.996 16.256 ;
      RECT MASK 1 13.268 15.184 13.328 16.256 ;
      RECT MASK 1 14.596 15.184 14.656 16.256 ;
      RECT MASK 1 14.928 15.184 14.988 16.256 ;
      RECT MASK 1 16.256 15.184 16.316 16.256 ;
      RECT MASK 1 16.588 15.184 16.648 16.256 ;
      RECT MASK 1 17.916 15.184 17.976 16.256 ;
      RECT MASK 1 18.248 15.184 18.308 16.256 ;
      RECT MASK 1 19.576 15.184 19.636 16.256 ;
      RECT MASK 1 19.908 15.184 19.968 16.256 ;
      RECT MASK 1 21.236 15.184 21.296 16.256 ;
      RECT MASK 1 21.568 15.184 21.628 16.256 ;
      RECT MASK 1 22.896 15.184 22.956 16.256 ;
      RECT MASK 1 23.228 15.184 23.288 16.256 ;
      RECT MASK 1 24.556 15.184 24.616 16.256 ;
      RECT MASK 1 24.888 15.184 24.948 16.256 ;
      RECT MASK 1 26.216 15.184 26.276 16.256 ;
      RECT MASK 1 26.548 15.184 26.608 16.256 ;
      RECT MASK 1 27.876 15.184 27.936 16.256 ;
      RECT MASK 1 28.208 15.184 28.268 16.256 ;
      RECT MASK 1 29.536 15.184 29.596 16.256 ;
      RECT MASK 1 29.868 15.184 29.928 16.256 ;
      RECT MASK 1 31.196 15.184 31.256 16.256 ;
      RECT MASK 1 31.528 15.184 31.588 16.256 ;
      RECT MASK 1 32.856 15.184 32.916 16.256 ;
      RECT MASK 1 33.188 15.184 33.248 16.256 ;
      RECT MASK 1 34.516 15.184 34.576 16.256 ;
      RECT MASK 1 34.848 15.184 34.908 16.256 ;
      RECT MASK 1 36.176 15.184 36.236 16.256 ;
      RECT MASK 1 36.508 15.184 36.568 16.256 ;
      RECT MASK 1 37.836 15.184 37.896 16.256 ;
      RECT MASK 1 38.168 15.184 38.228 16.256 ;
      RECT MASK 1 39.496 15.184 39.556 16.256 ;
      RECT MASK 1 39.828 15.184 39.888 16.256 ;
      RECT MASK 1 41.156 15.184 41.216 16.256 ;
      RECT MASK 1 41.488 15.184 41.548 16.256 ;
      RECT MASK 1 42.816 15.184 42.876 16.256 ;
      RECT MASK 1 43.148 15.184 43.208 16.256 ;
      RECT MASK 1 44.476 15.184 44.536 16.256 ;
      RECT MASK 1 44.808 15.184 44.868 16.256 ;
      RECT MASK 1 46.136 15.184 46.196 16.256 ;
      RECT MASK 1 46.468 15.184 46.528 16.256 ;
      RECT MASK 1 47.796 15.184 47.856 16.256 ;
      RECT MASK 1 48.128 15.184 48.188 16.256 ;
      RECT MASK 1 49.456 15.184 49.516 16.256 ;
      RECT MASK 1 49.788 15.184 49.848 16.256 ;
      RECT MASK 1 51.116 15.184 51.176 16.256 ;
      RECT MASK 1 51.448 15.184 51.508 16.256 ;
      RECT MASK 1 52.776 15.184 52.836 16.256 ;
      RECT MASK 1 53.108 15.184 53.168 16.256 ;
      RECT MASK 1 54.436 15.184 54.496 16.256 ;
      RECT MASK 1 54.768 15.184 54.828 16.256 ;
      RECT MASK 1 56.096 15.184 56.156 16.256 ;
      RECT MASK 1 56.594 15.184 56.654 16.256 ;
      RECT MASK 1 57.902 15.184 58.002 16.256 ;
      RECT MASK 1 58.234 15.184 58.334 16.256 ;
      RECT MASK 1 59.582 15.184 59.642 16.256 ;
      RECT MASK 1 59.748 15.184 59.808 16.256 ;
      RECT MASK 1 59.914 15.184 59.974 16.256 ;
      RECT MASK 1 60.578 15.184 60.638 16.256 ;
      RECT MASK 1 61.242 15.184 61.302 16.256 ;
      RECT MASK 1 61.574 15.184 61.634 16.256 ;
      RECT MASK 1 62.902 15.184 62.962 16.256 ;
      RECT MASK 1 63.234 15.184 63.294 16.256 ;
      RECT MASK 1 64.562 15.184 64.622 16.256 ;
      RECT MASK 1 64.894 15.184 64.954 16.256 ;
      RECT MASK 1 66.222 15.184 66.282 16.256 ;
      RECT MASK 1 66.554 15.184 66.614 16.256 ;
      RECT MASK 1 67.882 15.184 67.942 16.256 ;
      RECT MASK 1 68.214 15.184 68.274 16.256 ;
      RECT MASK 1 69.542 15.184 69.602 16.256 ;
      RECT MASK 1 69.874 15.184 69.934 16.256 ;
      RECT MASK 1 71.202 15.184 71.262 16.256 ;
      RECT MASK 1 71.534 15.184 71.594 16.256 ;
      RECT MASK 1 72.862 15.184 72.922 16.256 ;
      RECT MASK 1 73.194 15.184 73.254 16.256 ;
      RECT MASK 1 74.522 15.184 74.582 16.256 ;
      RECT MASK 1 74.854 15.184 74.914 16.256 ;
      RECT MASK 1 76.182 15.184 76.242 16.256 ;
      RECT MASK 1 76.514 15.184 76.574 16.256 ;
      RECT MASK 1 77.842 15.184 77.902 16.256 ;
      RECT MASK 1 78.174 15.184 78.234 16.256 ;
      RECT MASK 1 79.502 15.184 79.562 16.256 ;
      RECT MASK 1 79.834 15.184 79.894 16.256 ;
      RECT MASK 1 81.162 15.184 81.222 16.256 ;
      RECT MASK 1 81.494 15.184 81.554 16.256 ;
      RECT MASK 1 82.822 15.184 82.882 16.256 ;
      RECT MASK 1 83.154 15.184 83.214 16.256 ;
      RECT MASK 1 84.482 15.184 84.542 16.256 ;
      RECT MASK 1 84.814 15.184 84.874 16.256 ;
      RECT MASK 1 86.142 15.184 86.202 16.256 ;
      RECT MASK 1 86.474 15.184 86.534 16.256 ;
      RECT MASK 1 87.802 15.184 87.862 16.256 ;
      RECT MASK 1 88.134 15.184 88.194 16.256 ;
      RECT MASK 1 89.462 15.184 89.522 16.256 ;
      RECT MASK 1 89.794 15.184 89.854 16.256 ;
      RECT MASK 1 91.122 15.184 91.182 16.256 ;
      RECT MASK 1 91.454 15.184 91.514 16.256 ;
      RECT MASK 1 92.782 15.184 92.842 16.256 ;
      RECT MASK 1 93.114 15.184 93.174 16.256 ;
      RECT MASK 1 94.442 15.184 94.502 16.256 ;
      RECT MASK 1 94.774 15.184 94.834 16.256 ;
      RECT MASK 1 96.102 15.184 96.162 16.256 ;
      RECT MASK 1 96.434 15.184 96.494 16.256 ;
      RECT MASK 1 97.762 15.184 97.822 16.256 ;
      RECT MASK 1 98.094 15.184 98.154 16.256 ;
      RECT MASK 1 99.422 15.184 99.482 16.256 ;
      RECT MASK 1 99.754 15.184 99.814 16.256 ;
      RECT MASK 1 101.082 15.184 101.142 16.256 ;
      RECT MASK 1 101.414 15.184 101.474 16.256 ;
      RECT MASK 1 102.742 15.184 102.802 16.256 ;
      RECT MASK 1 103.074 15.184 103.134 16.256 ;
      RECT MASK 1 104.402 15.184 104.462 16.256 ;
      RECT MASK 1 104.734 15.184 104.794 16.256 ;
      RECT MASK 1 106.062 15.184 106.122 16.256 ;
      RECT MASK 1 106.394 15.184 106.454 16.256 ;
      RECT MASK 1 107.722 15.184 107.782 16.256 ;
      RECT MASK 1 108.054 15.184 108.114 16.256 ;
      RECT MASK 1 109.382 15.184 109.442 16.256 ;
      RECT MASK 1 109.714 15.184 109.774 16.256 ;
      RECT MASK 1 111.042 15.184 111.102 16.256 ;
      RECT MASK 1 111.208 15.184 111.268 16.256 ;
      RECT MASK 1 111.374 15.184 111.434 16.256 ;
      RECT MASK 1 5.466 15.359 5.526 16.081 ;
      RECT MASK 1 5.798 15.359 5.858 16.081 ;
      RECT MASK 1 6.462 15.359 6.522 16.081 ;
      RECT MASK 1 7.126 15.359 7.186 16.081 ;
      RECT MASK 1 7.292 15.359 7.352 16.081 ;
      RECT MASK 1 7.458 15.359 7.518 16.081 ;
      RECT MASK 1 8.122 15.359 8.182 16.081 ;
      RECT MASK 1 8.786 15.359 8.846 16.081 ;
      RECT MASK 1 8.952 15.359 9.012 16.081 ;
      RECT MASK 1 9.118 15.359 9.178 16.081 ;
      RECT MASK 1 9.782 15.359 9.842 16.081 ;
      RECT MASK 1 10.446 15.359 10.506 16.081 ;
      RECT MASK 1 10.778 15.359 10.838 16.081 ;
      RECT MASK 1 12.106 15.359 12.166 16.081 ;
      RECT MASK 1 12.438 15.359 12.498 16.081 ;
      RECT MASK 1 13.766 15.359 13.826 16.081 ;
      RECT MASK 1 14.098 15.359 14.158 16.081 ;
      RECT MASK 1 15.426 15.359 15.486 16.081 ;
      RECT MASK 1 15.758 15.359 15.818 16.081 ;
      RECT MASK 1 17.086 15.359 17.146 16.081 ;
      RECT MASK 1 17.418 15.359 17.478 16.081 ;
      RECT MASK 1 18.746 15.359 18.806 16.081 ;
      RECT MASK 1 19.078 15.359 19.138 16.081 ;
      RECT MASK 1 19.742 15.359 19.802 16.081 ;
      RECT MASK 1 20.406 15.359 20.466 16.081 ;
      RECT MASK 1 20.572 15.359 20.632 16.081 ;
      RECT MASK 1 20.738 15.359 20.798 16.081 ;
      RECT MASK 1 21.402 15.359 21.462 16.081 ;
      RECT MASK 1 22.066 15.359 22.126 16.081 ;
      RECT MASK 1 22.232 15.359 22.292 16.081 ;
      RECT MASK 1 22.398 15.359 22.458 16.081 ;
      RECT MASK 1 23.726 15.359 23.786 16.081 ;
      RECT MASK 1 24.058 15.359 24.118 16.081 ;
      RECT MASK 1 24.722 15.359 24.782 16.081 ;
      RECT MASK 1 25.386 15.359 25.446 16.081 ;
      RECT MASK 1 25.718 15.359 25.778 16.081 ;
      RECT MASK 1 26.382 15.359 26.442 16.081 ;
      RECT MASK 1 27.046 15.359 27.106 16.081 ;
      RECT MASK 1 27.378 15.359 27.438 16.081 ;
      RECT MASK 1 28.706 15.359 28.766 16.081 ;
      RECT MASK 1 29.038 15.359 29.098 16.081 ;
      RECT MASK 1 30.366 15.359 30.426 16.081 ;
      RECT MASK 1 30.698 15.359 30.758 16.081 ;
      RECT MASK 1 32.026 15.359 32.086 16.081 ;
      RECT MASK 1 32.192 15.359 32.252 16.081 ;
      RECT MASK 1 32.358 15.359 32.418 16.081 ;
      RECT MASK 1 33.022 15.359 33.082 16.081 ;
      RECT MASK 1 33.686 15.359 33.746 16.081 ;
      RECT MASK 1 33.852 15.359 33.912 16.081 ;
      RECT MASK 1 34.018 15.359 34.078 16.081 ;
      RECT MASK 1 34.682 15.359 34.742 16.081 ;
      RECT MASK 1 35.346 15.359 35.406 16.081 ;
      RECT MASK 1 35.512 15.359 35.572 16.081 ;
      RECT MASK 1 35.678 15.359 35.738 16.081 ;
      RECT MASK 1 36.342 15.359 36.402 16.081 ;
      RECT MASK 1 37.006 15.359 37.066 16.081 ;
      RECT MASK 1 37.338 15.359 37.398 16.081 ;
      RECT MASK 1 38.666 15.359 38.726 16.081 ;
      RECT MASK 1 38.998 15.359 39.058 16.081 ;
      RECT MASK 1 39.662 15.359 39.722 16.081 ;
      RECT MASK 1 40.326 15.359 40.386 16.081 ;
      RECT MASK 1 40.658 15.359 40.718 16.081 ;
      RECT MASK 1 41.986 15.359 42.046 16.081 ;
      RECT MASK 1 42.318 15.359 42.378 16.081 ;
      RECT MASK 1 43.646 15.359 43.706 16.081 ;
      RECT MASK 1 43.978 15.359 44.038 16.081 ;
      RECT MASK 1 45.306 15.359 45.366 16.081 ;
      RECT MASK 1 45.472 15.359 45.532 16.081 ;
      RECT MASK 1 45.638 15.359 45.698 16.081 ;
      RECT MASK 1 46.302 15.359 46.362 16.081 ;
      RECT MASK 1 46.966 15.359 47.026 16.081 ;
      RECT MASK 1 47.132 15.359 47.192 16.081 ;
      RECT MASK 1 47.298 15.359 47.358 16.081 ;
      RECT MASK 1 47.962 15.359 48.022 16.081 ;
      RECT MASK 1 48.626 15.359 48.686 16.081 ;
      RECT MASK 1 48.792 15.359 48.852 16.081 ;
      RECT MASK 1 48.958 15.359 49.018 16.081 ;
      RECT MASK 1 50.286 15.359 50.346 16.081 ;
      RECT MASK 1 50.618 15.359 50.678 16.081 ;
      RECT MASK 1 51.946 15.359 52.006 16.081 ;
      RECT MASK 1 52.278 15.359 52.338 16.081 ;
      RECT MASK 1 52.942 15.359 53.002 16.081 ;
      RECT MASK 1 53.606 15.359 53.666 16.081 ;
      RECT MASK 1 53.938 15.359 53.998 16.081 ;
      RECT MASK 1 55.266 15.359 55.326 16.081 ;
      RECT MASK 1 55.598 15.359 55.658 16.081 ;
      RECT MASK 1 56.262 15.359 56.322 16.081 ;
      RECT MASK 1 57.092 15.359 57.152 16.081 ;
      RECT MASK 1 57.424 15.359 57.484 16.081 ;
      RECT MASK 1 58.752 15.359 58.812 16.081 ;
      RECT MASK 1 59.084 15.359 59.144 16.081 ;
      RECT MASK 1 60.412 15.359 60.472 16.081 ;
      RECT MASK 1 60.744 15.359 60.804 16.081 ;
      RECT MASK 1 62.072 15.359 62.132 16.081 ;
      RECT MASK 1 62.238 15.359 62.298 16.081 ;
      RECT MASK 1 62.404 15.359 62.464 16.081 ;
      RECT MASK 1 63.068 15.359 63.128 16.081 ;
      RECT MASK 1 63.732 15.359 63.792 16.081 ;
      RECT MASK 1 64.064 15.359 64.124 16.081 ;
      RECT MASK 1 65.392 15.359 65.452 16.081 ;
      RECT MASK 1 65.724 15.359 65.784 16.081 ;
      RECT MASK 1 67.052 15.359 67.112 16.081 ;
      RECT MASK 1 67.384 15.359 67.444 16.081 ;
      RECT MASK 1 68.712 15.359 68.772 16.081 ;
      RECT MASK 1 69.044 15.359 69.104 16.081 ;
      RECT MASK 1 70.372 15.359 70.432 16.081 ;
      RECT MASK 1 70.704 15.359 70.764 16.081 ;
      RECT MASK 1 72.032 15.359 72.092 16.081 ;
      RECT MASK 1 72.364 15.359 72.424 16.081 ;
      RECT MASK 1 73.028 15.359 73.088 16.081 ;
      RECT MASK 1 73.692 15.359 73.752 16.081 ;
      RECT MASK 1 73.858 15.359 73.918 16.081 ;
      RECT MASK 1 74.024 15.359 74.084 16.081 ;
      RECT MASK 1 74.688 15.359 74.748 16.081 ;
      RECT MASK 1 75.352 15.359 75.412 16.081 ;
      RECT MASK 1 75.518 15.359 75.578 16.081 ;
      RECT MASK 1 75.684 15.359 75.744 16.081 ;
      RECT MASK 1 76.348 15.359 76.408 16.081 ;
      RECT MASK 1 77.012 15.359 77.072 16.081 ;
      RECT MASK 1 77.344 15.359 77.404 16.081 ;
      RECT MASK 1 78.672 15.359 78.732 16.081 ;
      RECT MASK 1 79.004 15.359 79.064 16.081 ;
      RECT MASK 1 80.332 15.359 80.392 16.081 ;
      RECT MASK 1 80.498 15.359 80.558 16.081 ;
      RECT MASK 1 80.664 15.359 80.724 16.081 ;
      RECT MASK 1 81.328 15.359 81.388 16.081 ;
      RECT MASK 1 81.992 15.359 82.052 16.081 ;
      RECT MASK 1 82.324 15.359 82.384 16.081 ;
      RECT MASK 1 82.988 15.359 83.048 16.081 ;
      RECT MASK 1 83.652 15.359 83.712 16.081 ;
      RECT MASK 1 83.984 15.359 84.044 16.081 ;
      RECT MASK 1 85.312 15.359 85.372 16.081 ;
      RECT MASK 1 85.478 15.359 85.538 16.081 ;
      RECT MASK 1 85.644 15.359 85.704 16.081 ;
      RECT MASK 1 86.308 15.359 86.368 16.081 ;
      RECT MASK 1 86.972 15.359 87.032 16.081 ;
      RECT MASK 1 87.138 15.359 87.198 16.081 ;
      RECT MASK 1 87.304 15.359 87.364 16.081 ;
      RECT MASK 1 87.968 15.359 88.028 16.081 ;
      RECT MASK 1 88.632 15.359 88.692 16.081 ;
      RECT MASK 1 88.798 15.359 88.858 16.081 ;
      RECT MASK 1 88.964 15.359 89.024 16.081 ;
      RECT MASK 1 89.628 15.359 89.688 16.081 ;
      RECT MASK 1 90.292 15.359 90.352 16.081 ;
      RECT MASK 1 90.624 15.359 90.684 16.081 ;
      RECT MASK 1 91.952 15.359 92.012 16.081 ;
      RECT MASK 1 92.284 15.359 92.344 16.081 ;
      RECT MASK 1 92.948 15.359 93.008 16.081 ;
      RECT MASK 1 93.612 15.359 93.672 16.081 ;
      RECT MASK 1 93.944 15.359 94.004 16.081 ;
      RECT MASK 1 95.272 15.359 95.332 16.081 ;
      RECT MASK 1 95.604 15.359 95.664 16.081 ;
      RECT MASK 1 96.932 15.359 96.992 16.081 ;
      RECT MASK 1 97.264 15.359 97.324 16.081 ;
      RECT MASK 1 98.592 15.359 98.652 16.081 ;
      RECT MASK 1 98.758 15.359 98.818 16.081 ;
      RECT MASK 1 98.924 15.359 98.984 16.081 ;
      RECT MASK 1 99.588 15.359 99.648 16.081 ;
      RECT MASK 1 100.252 15.359 100.312 16.081 ;
      RECT MASK 1 100.418 15.359 100.478 16.081 ;
      RECT MASK 1 100.584 15.359 100.644 16.081 ;
      RECT MASK 1 101.248 15.359 101.308 16.081 ;
      RECT MASK 1 101.912 15.359 101.972 16.081 ;
      RECT MASK 1 102.078 15.359 102.138 16.081 ;
      RECT MASK 1 102.244 15.359 102.304 16.081 ;
      RECT MASK 1 102.908 15.359 102.968 16.081 ;
      RECT MASK 1 103.572 15.359 103.632 16.081 ;
      RECT MASK 1 103.904 15.359 103.964 16.081 ;
      RECT MASK 1 105.232 15.359 105.292 16.081 ;
      RECT MASK 1 105.564 15.359 105.624 16.081 ;
      RECT MASK 1 106.228 15.359 106.288 16.081 ;
      RECT MASK 1 106.892 15.359 106.952 16.081 ;
      RECT MASK 1 107.224 15.359 107.284 16.081 ;
      RECT MASK 1 108.552 15.359 108.612 16.081 ;
      RECT MASK 1 108.884 15.359 108.944 16.081 ;
      RECT MASK 1 110.212 15.359 110.272 16.081 ;
      RECT MASK 1 110.544 15.359 110.604 16.081 ;
      RECT MASK 1 32.192 16.303 32.252 16.763 ;
      RECT MASK 1 45.472 16.309 45.532 16.763 ;
      RECT MASK 1 4.968 16.376 5.028 16.984 ;
      RECT MASK 1 5.3 16.376 5.36 16.984 ;
      RECT MASK 1 5.964 16.376 6.024 16.984 ;
      RECT MASK 1 6.296 16.376 6.356 16.984 ;
      RECT MASK 1 6.628 16.376 6.688 16.984 ;
      RECT MASK 1 6.96 16.376 7.02 16.984 ;
      RECT MASK 1 7.624 16.376 7.684 16.984 ;
      RECT MASK 1 7.956 16.376 8.016 16.984 ;
      RECT MASK 1 8.288 16.376 8.348 16.984 ;
      RECT MASK 1 8.62 16.376 8.68 16.984 ;
      RECT MASK 1 9.284 16.376 9.344 16.984 ;
      RECT MASK 1 9.616 16.376 9.676 16.984 ;
      RECT MASK 1 9.948 16.376 10.008 16.984 ;
      RECT MASK 1 10.28 16.376 10.34 16.984 ;
      RECT MASK 1 10.944 16.376 11.004 16.984 ;
      RECT MASK 1 11.276 16.376 11.336 16.984 ;
      RECT MASK 1 11.608 16.376 11.668 16.984 ;
      RECT MASK 1 11.94 16.376 12 16.984 ;
      RECT MASK 1 12.604 16.376 12.664 16.984 ;
      RECT MASK 1 12.936 16.376 12.996 16.984 ;
      RECT MASK 1 13.268 16.376 13.328 16.984 ;
      RECT MASK 1 13.6 16.376 13.66 16.984 ;
      RECT MASK 1 14.264 16.376 14.324 16.984 ;
      RECT MASK 1 14.596 16.376 14.656 16.984 ;
      RECT MASK 1 14.928 16.376 14.988 16.984 ;
      RECT MASK 1 15.26 16.376 15.32 16.984 ;
      RECT MASK 1 15.924 16.376 15.984 16.984 ;
      RECT MASK 1 16.256 16.376 16.316 16.984 ;
      RECT MASK 1 16.588 16.376 16.648 16.984 ;
      RECT MASK 1 16.92 16.376 16.98 16.984 ;
      RECT MASK 1 17.584 16.376 17.644 16.984 ;
      RECT MASK 1 17.916 16.376 17.976 16.984 ;
      RECT MASK 1 18.248 16.376 18.308 16.984 ;
      RECT MASK 1 18.58 16.376 18.64 16.984 ;
      RECT MASK 1 19.244 16.376 19.304 16.984 ;
      RECT MASK 1 19.576 16.376 19.636 16.984 ;
      RECT MASK 1 19.908 16.376 19.968 16.984 ;
      RECT MASK 1 20.24 16.376 20.3 16.984 ;
      RECT MASK 1 20.904 16.376 20.964 16.984 ;
      RECT MASK 1 21.236 16.376 21.296 16.984 ;
      RECT MASK 1 21.568 16.376 21.628 16.984 ;
      RECT MASK 1 21.9 16.376 21.96 16.984 ;
      RECT MASK 1 22.564 16.376 22.624 16.984 ;
      RECT MASK 1 22.896 16.376 22.956 16.984 ;
      RECT MASK 1 23.228 16.376 23.288 16.984 ;
      RECT MASK 1 23.56 16.376 23.62 16.984 ;
      RECT MASK 1 24.224 16.376 24.284 16.984 ;
      RECT MASK 1 24.556 16.376 24.616 16.984 ;
      RECT MASK 1 24.888 16.376 24.948 16.984 ;
      RECT MASK 1 25.22 16.376 25.28 16.984 ;
      RECT MASK 1 25.884 16.376 25.944 16.984 ;
      RECT MASK 1 26.216 16.376 26.276 16.984 ;
      RECT MASK 1 26.548 16.376 26.608 16.984 ;
      RECT MASK 1 26.88 16.376 26.94 16.984 ;
      RECT MASK 1 27.544 16.376 27.604 16.984 ;
      RECT MASK 1 27.876 16.376 27.936 16.984 ;
      RECT MASK 1 28.208 16.376 28.268 16.984 ;
      RECT MASK 1 28.54 16.376 28.6 16.984 ;
      RECT MASK 1 29.204 16.376 29.264 16.984 ;
      RECT MASK 1 29.536 16.376 29.596 16.984 ;
      RECT MASK 1 29.868 16.376 29.928 16.984 ;
      RECT MASK 1 30.2 16.376 30.26 16.984 ;
      RECT MASK 1 30.864 16.376 30.924 16.984 ;
      RECT MASK 1 31.196 16.376 31.256 16.984 ;
      RECT MASK 1 31.528 16.376 31.588 16.984 ;
      RECT MASK 1 31.86 16.376 31.92 16.984 ;
      RECT MASK 1 32.524 16.376 32.584 16.984 ;
      RECT MASK 1 32.856 16.376 32.916 16.984 ;
      RECT MASK 1 33.188 16.376 33.248 16.984 ;
      RECT MASK 1 33.52 16.376 33.58 16.984 ;
      RECT MASK 1 34.184 16.376 34.244 16.984 ;
      RECT MASK 1 34.516 16.376 34.576 16.984 ;
      RECT MASK 1 34.848 16.376 34.908 16.984 ;
      RECT MASK 1 35.18 16.376 35.24 16.984 ;
      RECT MASK 1 35.844 16.376 35.904 16.984 ;
      RECT MASK 1 36.176 16.376 36.236 16.984 ;
      RECT MASK 1 36.508 16.376 36.568 16.984 ;
      RECT MASK 1 36.84 16.376 36.9 16.984 ;
      RECT MASK 1 37.504 16.376 37.564 16.984 ;
      RECT MASK 1 37.836 16.376 37.896 16.984 ;
      RECT MASK 1 38.168 16.376 38.228 16.984 ;
      RECT MASK 1 38.5 16.376 38.56 16.984 ;
      RECT MASK 1 39.164 16.376 39.224 16.984 ;
      RECT MASK 1 39.496 16.376 39.556 16.984 ;
      RECT MASK 1 39.828 16.376 39.888 16.984 ;
      RECT MASK 1 40.16 16.376 40.22 16.984 ;
      RECT MASK 1 40.824 16.376 40.884 16.984 ;
      RECT MASK 1 41.156 16.376 41.216 16.984 ;
      RECT MASK 1 41.488 16.376 41.548 16.984 ;
      RECT MASK 1 41.82 16.376 41.88 16.984 ;
      RECT MASK 1 42.484 16.376 42.544 16.984 ;
      RECT MASK 1 42.816 16.376 42.876 16.984 ;
      RECT MASK 1 43.148 16.376 43.208 16.984 ;
      RECT MASK 1 43.48 16.376 43.54 16.984 ;
      RECT MASK 1 44.144 16.376 44.204 16.984 ;
      RECT MASK 1 44.476 16.376 44.536 16.984 ;
      RECT MASK 1 44.808 16.376 44.868 16.984 ;
      RECT MASK 1 45.14 16.376 45.2 16.984 ;
      RECT MASK 1 45.804 16.376 45.864 16.984 ;
      RECT MASK 1 46.136 16.376 46.196 16.984 ;
      RECT MASK 1 46.468 16.376 46.528 16.984 ;
      RECT MASK 1 46.8 16.376 46.86 16.984 ;
      RECT MASK 1 47.464 16.376 47.524 16.984 ;
      RECT MASK 1 47.796 16.376 47.856 16.984 ;
      RECT MASK 1 48.128 16.376 48.188 16.984 ;
      RECT MASK 1 48.46 16.376 48.52 16.984 ;
      RECT MASK 1 49.124 16.376 49.184 16.984 ;
      RECT MASK 1 49.456 16.376 49.516 16.984 ;
      RECT MASK 1 49.788 16.376 49.848 16.984 ;
      RECT MASK 1 50.12 16.376 50.18 16.984 ;
      RECT MASK 1 50.784 16.376 50.844 16.984 ;
      RECT MASK 1 51.116 16.376 51.176 16.984 ;
      RECT MASK 1 51.448 16.376 51.508 16.984 ;
      RECT MASK 1 51.78 16.376 51.84 16.984 ;
      RECT MASK 1 52.444 16.376 52.504 16.984 ;
      RECT MASK 1 52.776 16.376 52.836 16.984 ;
      RECT MASK 1 53.108 16.376 53.168 16.984 ;
      RECT MASK 1 53.44 16.376 53.5 16.984 ;
      RECT MASK 1 54.104 16.376 54.164 16.984 ;
      RECT MASK 1 54.436 16.376 54.496 16.984 ;
      RECT MASK 1 54.768 16.376 54.828 16.984 ;
      RECT MASK 1 55.1 16.376 55.16 16.984 ;
      RECT MASK 1 55.764 16.376 55.824 16.984 ;
      RECT MASK 1 56.096 16.376 56.156 16.984 ;
      RECT MASK 1 56.594 16.376 56.654 16.984 ;
      RECT MASK 1 56.926 16.376 56.986 16.984 ;
      RECT MASK 1 57.59 16.376 57.65 16.984 ;
      RECT MASK 1 57.922 16.376 57.982 16.984 ;
      RECT MASK 1 58.254 16.376 58.314 16.984 ;
      RECT MASK 1 58.586 16.376 58.646 16.984 ;
      RECT MASK 1 59.25 16.376 59.31 16.984 ;
      RECT MASK 1 59.582 16.376 59.642 16.984 ;
      RECT MASK 1 59.914 16.376 59.974 16.984 ;
      RECT MASK 1 60.246 16.376 60.306 16.984 ;
      RECT MASK 1 60.91 16.376 60.97 16.984 ;
      RECT MASK 1 61.242 16.376 61.302 16.984 ;
      RECT MASK 1 61.574 16.376 61.634 16.984 ;
      RECT MASK 1 61.906 16.376 61.966 16.984 ;
      RECT MASK 1 62.57 16.376 62.63 16.984 ;
      RECT MASK 1 62.902 16.376 62.962 16.984 ;
      RECT MASK 1 63.234 16.376 63.294 16.984 ;
      RECT MASK 1 63.566 16.376 63.626 16.984 ;
      RECT MASK 1 64.23 16.376 64.29 16.984 ;
      RECT MASK 1 64.562 16.376 64.622 16.984 ;
      RECT MASK 1 64.894 16.376 64.954 16.984 ;
      RECT MASK 1 65.226 16.376 65.286 16.984 ;
      RECT MASK 1 65.89 16.376 65.95 16.984 ;
      RECT MASK 1 66.222 16.376 66.282 16.984 ;
      RECT MASK 1 66.554 16.376 66.614 16.984 ;
      RECT MASK 1 66.886 16.376 66.946 16.984 ;
      RECT MASK 1 67.55 16.376 67.61 16.984 ;
      RECT MASK 1 67.882 16.376 67.942 16.984 ;
      RECT MASK 1 68.214 16.376 68.274 16.984 ;
      RECT MASK 1 68.546 16.376 68.606 16.984 ;
      RECT MASK 1 69.21 16.376 69.27 16.984 ;
      RECT MASK 1 69.542 16.376 69.602 16.984 ;
      RECT MASK 1 69.874 16.376 69.934 16.984 ;
      RECT MASK 1 70.206 16.376 70.266 16.984 ;
      RECT MASK 1 70.87 16.376 70.93 16.984 ;
      RECT MASK 1 71.202 16.376 71.262 16.984 ;
      RECT MASK 1 71.534 16.376 71.594 16.984 ;
      RECT MASK 1 71.866 16.376 71.926 16.984 ;
      RECT MASK 1 72.53 16.376 72.59 16.984 ;
      RECT MASK 1 72.862 16.376 72.922 16.984 ;
      RECT MASK 1 73.194 16.376 73.254 16.984 ;
      RECT MASK 1 73.526 16.376 73.586 16.984 ;
      RECT MASK 1 74.19 16.376 74.25 16.984 ;
      RECT MASK 1 74.522 16.376 74.582 16.984 ;
      RECT MASK 1 74.854 16.376 74.914 16.984 ;
      RECT MASK 1 75.186 16.376 75.246 16.984 ;
      RECT MASK 1 75.85 16.376 75.91 16.984 ;
      RECT MASK 1 76.182 16.376 76.242 16.984 ;
      RECT MASK 1 76.514 16.376 76.574 16.984 ;
      RECT MASK 1 76.846 16.376 76.906 16.984 ;
      RECT MASK 1 77.51 16.376 77.57 16.984 ;
      RECT MASK 1 77.842 16.376 77.902 16.984 ;
      RECT MASK 1 78.174 16.376 78.234 16.984 ;
      RECT MASK 1 78.506 16.376 78.566 16.984 ;
      RECT MASK 1 79.17 16.376 79.23 16.984 ;
      RECT MASK 1 79.502 16.376 79.562 16.984 ;
      RECT MASK 1 79.834 16.376 79.894 16.984 ;
      RECT MASK 1 80.166 16.376 80.226 16.984 ;
      RECT MASK 1 80.83 16.376 80.89 16.984 ;
      RECT MASK 1 81.162 16.376 81.222 16.984 ;
      RECT MASK 1 81.494 16.376 81.554 16.984 ;
      RECT MASK 1 81.826 16.376 81.886 16.984 ;
      RECT MASK 1 82.49 16.376 82.55 16.984 ;
      RECT MASK 1 82.822 16.376 82.882 16.984 ;
      RECT MASK 1 83.154 16.376 83.214 16.984 ;
      RECT MASK 1 83.486 16.376 83.546 16.984 ;
      RECT MASK 1 84.15 16.376 84.21 16.984 ;
      RECT MASK 1 84.482 16.376 84.542 16.984 ;
      RECT MASK 1 84.814 16.376 84.874 16.984 ;
      RECT MASK 1 85.146 16.376 85.206 16.984 ;
      RECT MASK 1 85.81 16.376 85.87 16.984 ;
      RECT MASK 1 86.142 16.376 86.202 16.984 ;
      RECT MASK 1 86.474 16.376 86.534 16.984 ;
      RECT MASK 1 86.806 16.376 86.866 16.984 ;
      RECT MASK 1 87.47 16.376 87.53 16.984 ;
      RECT MASK 1 87.802 16.376 87.862 16.984 ;
      RECT MASK 1 88.134 16.376 88.194 16.984 ;
      RECT MASK 1 88.466 16.376 88.526 16.984 ;
      RECT MASK 1 89.13 16.376 89.19 16.984 ;
      RECT MASK 1 89.462 16.376 89.522 16.984 ;
      RECT MASK 1 89.794 16.376 89.854 16.984 ;
      RECT MASK 1 90.126 16.376 90.186 16.984 ;
      RECT MASK 1 90.79 16.376 90.85 16.984 ;
      RECT MASK 1 91.122 16.376 91.182 16.984 ;
      RECT MASK 1 91.454 16.376 91.514 16.984 ;
      RECT MASK 1 91.786 16.376 91.846 16.984 ;
      RECT MASK 1 92.45 16.376 92.51 16.984 ;
      RECT MASK 1 92.782 16.376 92.842 16.984 ;
      RECT MASK 1 93.114 16.376 93.174 16.984 ;
      RECT MASK 1 93.446 16.376 93.506 16.984 ;
      RECT MASK 1 94.11 16.376 94.17 16.984 ;
      RECT MASK 1 94.442 16.376 94.502 16.984 ;
      RECT MASK 1 94.774 16.376 94.834 16.984 ;
      RECT MASK 1 95.106 16.376 95.166 16.984 ;
      RECT MASK 1 95.77 16.376 95.83 16.984 ;
      RECT MASK 1 96.102 16.376 96.162 16.984 ;
      RECT MASK 1 96.434 16.376 96.494 16.984 ;
      RECT MASK 1 96.766 16.376 96.826 16.984 ;
      RECT MASK 1 97.43 16.376 97.49 16.984 ;
      RECT MASK 1 97.762 16.376 97.822 16.984 ;
      RECT MASK 1 98.094 16.376 98.154 16.984 ;
      RECT MASK 1 98.426 16.376 98.486 16.984 ;
      RECT MASK 1 99.09 16.376 99.15 16.984 ;
      RECT MASK 1 99.422 16.376 99.482 16.984 ;
      RECT MASK 1 99.754 16.376 99.814 16.984 ;
      RECT MASK 1 100.086 16.376 100.146 16.984 ;
      RECT MASK 1 100.75 16.376 100.81 16.984 ;
      RECT MASK 1 101.082 16.376 101.142 16.984 ;
      RECT MASK 1 101.414 16.376 101.474 16.984 ;
      RECT MASK 1 101.746 16.376 101.806 16.984 ;
      RECT MASK 1 102.41 16.376 102.47 16.984 ;
      RECT MASK 1 102.742 16.376 102.802 16.984 ;
      RECT MASK 1 103.074 16.376 103.134 16.984 ;
      RECT MASK 1 103.406 16.376 103.466 16.984 ;
      RECT MASK 1 104.07 16.376 104.13 16.984 ;
      RECT MASK 1 104.402 16.376 104.462 16.984 ;
      RECT MASK 1 104.734 16.376 104.794 16.984 ;
      RECT MASK 1 105.066 16.376 105.126 16.984 ;
      RECT MASK 1 105.73 16.376 105.79 16.984 ;
      RECT MASK 1 106.062 16.376 106.122 16.984 ;
      RECT MASK 1 106.394 16.376 106.454 16.984 ;
      RECT MASK 1 106.726 16.376 106.786 16.984 ;
      RECT MASK 1 107.39 16.376 107.45 16.984 ;
      RECT MASK 1 107.722 16.376 107.782 16.984 ;
      RECT MASK 1 108.054 16.376 108.114 16.984 ;
      RECT MASK 1 108.386 16.376 108.446 16.984 ;
      RECT MASK 1 109.05 16.376 109.11 16.984 ;
      RECT MASK 1 109.382 16.376 109.442 16.984 ;
      RECT MASK 1 109.714 16.376 109.774 16.984 ;
      RECT MASK 1 110.046 16.376 110.106 16.984 ;
      RECT MASK 1 110.71 16.376 110.77 16.984 ;
      RECT MASK 1 111.042 16.376 111.102 16.984 ;
      RECT MASK 1 4.387 16.8425 4.447 17.76 ;
      RECT MASK 1 111.623 16.8425 111.683 17.76 ;
      RECT MASK 1 37.172 16.969 37.232 17.429 ;
      RECT MASK 1 109.548 16.9705 109.608 17.429 ;
      RECT MASK 1 42.982 16.9775 43.042 17.429 ;
      RECT MASK 1 10.612 16.981 10.672 17.429 ;
      RECT MASK 1 16.422 16.981 16.482 17.429 ;
      RECT MASK 1 22.232 16.981 22.292 17.429 ;
      RECT MASK 1 29.702 16.981 29.762 17.429 ;
      RECT MASK 1 50.452 16.981 50.512 17.429 ;
      RECT MASK 1 56.428 16.981 56.488 17.429 ;
      RECT MASK 1 63.898 16.981 63.958 17.429 ;
      RECT MASK 1 69.708 16.981 69.768 17.429 ;
      RECT MASK 1 77.178 16.981 77.238 17.429 ;
      RECT MASK 1 81.328 16.981 81.388 17.429 ;
      RECT MASK 1 82.988 16.981 83.048 17.429 ;
      RECT MASK 1 90.458 16.981 90.518 17.429 ;
      RECT MASK 1 96.268 16.981 96.328 17.429 ;
      RECT MASK 1 103.738 16.981 103.798 17.429 ;
      RECT MASK 1 67.208 17.075 67.288 17.76 ;
      RECT MASK 1 4.636 17.104 4.696 17.76 ;
      RECT MASK 1 4.802 17.104 4.862 17.76 ;
      RECT MASK 1 4.968 17.104 5.028 17.76 ;
      RECT MASK 1 5.632 17.104 5.692 17.76 ;
      RECT MASK 1 6.296 17.104 6.356 17.76 ;
      RECT MASK 1 6.462 17.104 6.522 17.76 ;
      RECT MASK 1 6.628 17.104 6.688 17.76 ;
      RECT MASK 1 7.292 17.104 7.352 17.76 ;
      RECT MASK 1 7.956 17.104 8.016 17.76 ;
      RECT MASK 1 8.122 17.104 8.182 17.76 ;
      RECT MASK 1 8.288 17.104 8.348 17.76 ;
      RECT MASK 1 8.952 17.104 9.012 17.76 ;
      RECT MASK 1 9.616 17.104 9.676 17.76 ;
      RECT MASK 1 9.782 17.104 9.842 17.76 ;
      RECT MASK 1 9.948 17.104 10.008 17.76 ;
      RECT MASK 1 11.276 17.104 11.336 17.76 ;
      RECT MASK 1 11.442 17.104 11.502 17.76 ;
      RECT MASK 1 11.608 17.104 11.668 17.76 ;
      RECT MASK 1 12.272 17.104 12.332 17.76 ;
      RECT MASK 1 12.936 17.104 12.996 17.76 ;
      RECT MASK 1 13.102 17.104 13.162 17.76 ;
      RECT MASK 1 13.268 17.104 13.328 17.76 ;
      RECT MASK 1 13.932 17.104 13.992 17.76 ;
      RECT MASK 1 14.596 17.104 14.656 17.76 ;
      RECT MASK 1 14.762 17.104 14.822 17.76 ;
      RECT MASK 1 14.928 17.104 14.988 17.76 ;
      RECT MASK 1 15.592 17.104 15.652 17.76 ;
      RECT MASK 1 16.256 17.104 16.316 17.76 ;
      RECT MASK 1 16.588 17.104 16.648 17.76 ;
      RECT MASK 1 17.252 17.104 17.312 17.76 ;
      RECT MASK 1 17.916 17.104 17.976 17.76 ;
      RECT MASK 1 18.082 17.104 18.142 17.76 ;
      RECT MASK 1 18.248 17.104 18.308 17.76 ;
      RECT MASK 1 18.912 17.104 18.972 17.76 ;
      RECT MASK 1 19.576 17.104 19.636 17.76 ;
      RECT MASK 1 19.742 17.104 19.802 17.76 ;
      RECT MASK 1 19.908 17.104 19.968 17.76 ;
      RECT MASK 1 20.572 17.104 20.632 17.76 ;
      RECT MASK 1 21.236 17.104 21.296 17.76 ;
      RECT MASK 1 21.402 17.104 21.462 17.76 ;
      RECT MASK 1 21.568 17.104 21.628 17.76 ;
      RECT MASK 1 22.896 17.104 22.956 17.76 ;
      RECT MASK 1 23.062 17.104 23.122 17.76 ;
      RECT MASK 1 23.228 17.104 23.288 17.76 ;
      RECT MASK 1 24.556 17.104 24.616 17.76 ;
      RECT MASK 1 24.722 17.104 24.782 17.76 ;
      RECT MASK 1 24.888 17.104 24.948 17.76 ;
      RECT MASK 1 25.552 17.104 25.612 17.76 ;
      RECT MASK 1 26.216 17.104 26.276 17.76 ;
      RECT MASK 1 26.382 17.104 26.442 17.76 ;
      RECT MASK 1 26.548 17.104 26.608 17.76 ;
      RECT MASK 1 27.212 17.104 27.272 17.76 ;
      RECT MASK 1 27.876 17.104 27.936 17.76 ;
      RECT MASK 1 28.042 17.104 28.102 17.76 ;
      RECT MASK 1 28.208 17.104 28.268 17.76 ;
      RECT MASK 1 28.872 17.104 28.932 17.76 ;
      RECT MASK 1 29.536 17.104 29.596 17.76 ;
      RECT MASK 1 29.868 17.104 29.928 17.76 ;
      RECT MASK 1 30.532 17.104 30.592 17.76 ;
      RECT MASK 1 31.196 17.104 31.256 17.76 ;
      RECT MASK 1 31.528 17.104 31.588 17.76 ;
      RECT MASK 1 32.192 17.104 32.252 17.76 ;
      RECT MASK 1 32.856 17.104 32.916 17.76 ;
      RECT MASK 1 33.022 17.104 33.082 17.76 ;
      RECT MASK 1 33.188 17.104 33.248 17.76 ;
      RECT MASK 1 33.852 17.104 33.912 17.76 ;
      RECT MASK 1 34.516 17.104 34.576 17.76 ;
      RECT MASK 1 34.682 17.104 34.742 17.76 ;
      RECT MASK 1 34.848 17.104 34.908 17.76 ;
      RECT MASK 1 35.512 17.104 35.572 17.76 ;
      RECT MASK 1 36.176 17.104 36.236 17.76 ;
      RECT MASK 1 36.342 17.104 36.402 17.76 ;
      RECT MASK 1 36.508 17.104 36.568 17.76 ;
      RECT MASK 1 37.836 17.104 37.896 17.76 ;
      RECT MASK 1 38.002 17.104 38.062 17.76 ;
      RECT MASK 1 38.168 17.104 38.228 17.76 ;
      RECT MASK 1 38.832 17.104 38.892 17.76 ;
      RECT MASK 1 39.496 17.104 39.556 17.76 ;
      RECT MASK 1 39.662 17.104 39.722 17.76 ;
      RECT MASK 1 39.828 17.104 39.888 17.76 ;
      RECT MASK 1 40.492 17.104 40.552 17.76 ;
      RECT MASK 1 41.156 17.104 41.216 17.76 ;
      RECT MASK 1 41.322 17.104 41.382 17.76 ;
      RECT MASK 1 41.488 17.104 41.548 17.76 ;
      RECT MASK 1 42.152 17.104 42.212 17.76 ;
      RECT MASK 1 42.816 17.104 42.876 17.76 ;
      RECT MASK 1 43.148 17.104 43.208 17.76 ;
      RECT MASK 1 43.812 17.104 43.872 17.76 ;
      RECT MASK 1 44.476 17.104 44.536 17.76 ;
      RECT MASK 1 44.642 17.104 44.702 17.76 ;
      RECT MASK 1 44.808 17.104 44.868 17.76 ;
      RECT MASK 1 45.472 17.104 45.532 17.76 ;
      RECT MASK 1 46.136 17.104 46.196 17.76 ;
      RECT MASK 1 46.302 17.104 46.362 17.76 ;
      RECT MASK 1 46.468 17.104 46.528 17.76 ;
      RECT MASK 1 47.132 17.104 47.192 17.76 ;
      RECT MASK 1 47.796 17.104 47.856 17.76 ;
      RECT MASK 1 47.962 17.104 48.022 17.76 ;
      RECT MASK 1 48.128 17.104 48.188 17.76 ;
      RECT MASK 1 48.792 17.104 48.852 17.76 ;
      RECT MASK 1 49.456 17.104 49.516 17.76 ;
      RECT MASK 1 49.622 17.104 49.682 17.76 ;
      RECT MASK 1 49.788 17.104 49.848 17.76 ;
      RECT MASK 1 51.116 17.104 51.176 17.76 ;
      RECT MASK 1 51.282 17.104 51.342 17.76 ;
      RECT MASK 1 51.448 17.104 51.508 17.76 ;
      RECT MASK 1 52.112 17.104 52.172 17.76 ;
      RECT MASK 1 52.776 17.104 52.836 17.76 ;
      RECT MASK 1 52.942 17.104 53.002 17.76 ;
      RECT MASK 1 53.108 17.104 53.168 17.76 ;
      RECT MASK 1 53.772 17.104 53.832 17.76 ;
      RECT MASK 1 54.436 17.104 54.496 17.76 ;
      RECT MASK 1 54.602 17.104 54.662 17.76 ;
      RECT MASK 1 54.768 17.104 54.828 17.76 ;
      RECT MASK 1 55.432 17.104 55.492 17.76 ;
      RECT MASK 1 56.096 17.104 56.156 17.76 ;
      RECT MASK 1 56.262 17.104 56.322 17.76 ;
      RECT MASK 1 56.594 17.104 56.654 17.76 ;
      RECT MASK 1 57.258 17.104 57.318 17.76 ;
      RECT MASK 1 57.922 17.104 57.982 17.76 ;
      RECT MASK 1 58.254 17.104 58.314 17.76 ;
      RECT MASK 1 58.918 17.104 58.978 17.76 ;
      RECT MASK 1 59.582 17.104 59.642 17.76 ;
      RECT MASK 1 59.748 17.104 59.808 17.76 ;
      RECT MASK 1 59.914 17.104 59.974 17.76 ;
      RECT MASK 1 60.578 17.104 60.638 17.76 ;
      RECT MASK 1 61.242 17.104 61.302 17.76 ;
      RECT MASK 1 61.408 17.104 61.468 17.76 ;
      RECT MASK 1 61.574 17.104 61.634 17.76 ;
      RECT MASK 1 62.238 17.104 62.298 17.76 ;
      RECT MASK 1 62.902 17.104 62.962 17.76 ;
      RECT MASK 1 63.068 17.104 63.128 17.76 ;
      RECT MASK 1 63.234 17.104 63.294 17.76 ;
      RECT MASK 1 64.562 17.104 64.622 17.76 ;
      RECT MASK 1 64.728 17.104 64.788 17.76 ;
      RECT MASK 1 64.894 17.104 64.954 17.76 ;
      RECT MASK 1 65.558 17.104 65.618 17.76 ;
      RECT MASK 1 66.212 17.104 66.292 17.76 ;
      RECT MASK 1 66.378 17.104 66.458 17.76 ;
      RECT MASK 1 66.544 17.104 66.624 17.76 ;
      RECT MASK 1 67.882 17.104 67.942 17.76 ;
      RECT MASK 1 68.048 17.104 68.108 17.76 ;
      RECT MASK 1 68.214 17.104 68.274 17.76 ;
      RECT MASK 1 68.878 17.104 68.938 17.76 ;
      RECT MASK 1 69.542 17.104 69.602 17.76 ;
      RECT MASK 1 69.874 17.104 69.934 17.76 ;
      RECT MASK 1 70.538 17.104 70.598 17.76 ;
      RECT MASK 1 71.202 17.104 71.262 17.76 ;
      RECT MASK 1 71.534 17.104 71.594 17.76 ;
      RECT MASK 1 72.198 17.104 72.258 17.76 ;
      RECT MASK 1 72.862 17.104 72.922 17.76 ;
      RECT MASK 1 73.028 17.104 73.088 17.76 ;
      RECT MASK 1 73.194 17.104 73.254 17.76 ;
      RECT MASK 1 73.858 17.104 73.918 17.76 ;
      RECT MASK 1 74.522 17.104 74.582 17.76 ;
      RECT MASK 1 74.688 17.104 74.748 17.76 ;
      RECT MASK 1 74.854 17.104 74.914 17.76 ;
      RECT MASK 1 75.518 17.104 75.578 17.76 ;
      RECT MASK 1 76.182 17.104 76.242 17.76 ;
      RECT MASK 1 76.348 17.104 76.408 17.76 ;
      RECT MASK 1 76.514 17.104 76.574 17.76 ;
      RECT MASK 1 77.842 17.104 77.902 17.76 ;
      RECT MASK 1 78.174 17.104 78.234 17.76 ;
      RECT MASK 1 78.838 17.104 78.898 17.76 ;
      RECT MASK 1 79.502 17.104 79.562 17.76 ;
      RECT MASK 1 79.668 17.104 79.728 17.76 ;
      RECT MASK 1 79.834 17.104 79.894 17.76 ;
      RECT MASK 1 80.498 17.104 80.558 17.76 ;
      RECT MASK 1 81.162 17.104 81.222 17.76 ;
      RECT MASK 1 81.494 17.104 81.554 17.76 ;
      RECT MASK 1 82.158 17.104 82.218 17.76 ;
      RECT MASK 1 82.822 17.104 82.882 17.76 ;
      RECT MASK 1 83.154 17.104 83.214 17.76 ;
      RECT MASK 1 83.818 17.104 83.878 17.76 ;
      RECT MASK 1 84.482 17.104 84.542 17.76 ;
      RECT MASK 1 84.648 17.104 84.708 17.76 ;
      RECT MASK 1 84.814 17.104 84.874 17.76 ;
      RECT MASK 1 85.478 17.104 85.538 17.76 ;
      RECT MASK 1 86.142 17.104 86.202 17.76 ;
      RECT MASK 1 86.308 17.104 86.368 17.76 ;
      RECT MASK 1 86.474 17.104 86.534 17.76 ;
      RECT MASK 1 87.138 17.104 87.198 17.76 ;
      RECT MASK 1 87.802 17.104 87.862 17.76 ;
      RECT MASK 1 87.968 17.104 88.028 17.76 ;
      RECT MASK 1 88.134 17.104 88.194 17.76 ;
      RECT MASK 1 88.798 17.104 88.858 17.76 ;
      RECT MASK 1 89.462 17.104 89.522 17.76 ;
      RECT MASK 1 89.628 17.104 89.688 17.76 ;
      RECT MASK 1 89.794 17.104 89.854 17.76 ;
      RECT MASK 1 91.122 17.104 91.182 17.76 ;
      RECT MASK 1 91.288 17.104 91.348 17.76 ;
      RECT MASK 1 91.454 17.104 91.514 17.76 ;
      RECT MASK 1 92.118 17.104 92.178 17.76 ;
      RECT MASK 1 92.782 17.104 92.842 17.76 ;
      RECT MASK 1 92.948 17.104 93.008 17.76 ;
      RECT MASK 1 93.114 17.104 93.174 17.76 ;
      RECT MASK 1 93.778 17.104 93.838 17.76 ;
      RECT MASK 1 94.442 17.104 94.502 17.76 ;
      RECT MASK 1 94.608 17.104 94.668 17.76 ;
      RECT MASK 1 94.774 17.104 94.834 17.76 ;
      RECT MASK 1 95.438 17.104 95.498 17.76 ;
      RECT MASK 1 96.102 17.104 96.162 17.76 ;
      RECT MASK 1 96.434 17.104 96.494 17.76 ;
      RECT MASK 1 97.098 17.104 97.158 17.76 ;
      RECT MASK 1 97.762 17.104 97.822 17.76 ;
      RECT MASK 1 97.928 17.104 97.988 17.76 ;
      RECT MASK 1 98.094 17.104 98.154 17.76 ;
      RECT MASK 1 98.758 17.104 98.818 17.76 ;
      RECT MASK 1 99.422 17.104 99.482 17.76 ;
      RECT MASK 1 99.588 17.104 99.648 17.76 ;
      RECT MASK 1 99.754 17.104 99.814 17.76 ;
      RECT MASK 1 100.418 17.104 100.478 17.76 ;
      RECT MASK 1 101.082 17.104 101.142 17.76 ;
      RECT MASK 1 101.248 17.104 101.308 17.76 ;
      RECT MASK 1 101.414 17.104 101.474 17.76 ;
      RECT MASK 1 102.078 17.104 102.138 17.76 ;
      RECT MASK 1 102.742 17.104 102.802 17.76 ;
      RECT MASK 1 102.908 17.104 102.968 17.76 ;
      RECT MASK 1 103.074 17.104 103.134 17.76 ;
      RECT MASK 1 104.402 17.104 104.462 17.76 ;
      RECT MASK 1 104.568 17.104 104.628 17.76 ;
      RECT MASK 1 104.734 17.104 104.794 17.76 ;
      RECT MASK 1 105.398 17.104 105.458 17.76 ;
      RECT MASK 1 106.062 17.104 106.122 17.76 ;
      RECT MASK 1 106.228 17.104 106.288 17.76 ;
      RECT MASK 1 106.394 17.104 106.454 17.76 ;
      RECT MASK 1 107.058 17.104 107.118 17.76 ;
      RECT MASK 1 107.722 17.104 107.782 17.76 ;
      RECT MASK 1 107.888 17.104 107.948 17.76 ;
      RECT MASK 1 108.054 17.104 108.114 17.76 ;
      RECT MASK 1 108.718 17.104 108.778 17.76 ;
      RECT MASK 1 109.382 17.104 109.442 17.76 ;
      RECT MASK 1 109.714 17.104 109.774 17.76 ;
      RECT MASK 1 110.378 17.104 110.438 17.76 ;
      RECT MASK 1 111.042 17.104 111.102 17.76 ;
      RECT MASK 1 111.208 17.104 111.268 17.76 ;
      RECT MASK 1 111.374 17.104 111.434 17.76 ;
      RECT MASK 1 5.466 17.279 5.526 17.76 ;
      RECT MASK 1 5.798 17.279 5.858 17.76 ;
      RECT MASK 1 7.126 17.279 7.186 17.76 ;
      RECT MASK 1 7.458 17.279 7.518 17.76 ;
      RECT MASK 1 8.786 17.279 8.846 17.76 ;
      RECT MASK 1 9.118 17.279 9.178 17.76 ;
      RECT MASK 1 10.446 17.279 10.506 17.76 ;
      RECT MASK 1 10.778 17.279 10.838 17.76 ;
      RECT MASK 1 12.106 17.279 12.166 17.76 ;
      RECT MASK 1 12.438 17.279 12.498 17.76 ;
      RECT MASK 1 13.766 17.279 13.826 17.76 ;
      RECT MASK 1 14.098 17.279 14.158 17.76 ;
      RECT MASK 1 15.426 17.279 15.486 17.76 ;
      RECT MASK 1 15.758 17.279 15.818 17.76 ;
      RECT MASK 1 17.086 17.279 17.146 17.76 ;
      RECT MASK 1 17.418 17.279 17.478 17.76 ;
      RECT MASK 1 18.746 17.279 18.806 17.76 ;
      RECT MASK 1 19.078 17.279 19.138 17.76 ;
      RECT MASK 1 20.406 17.279 20.466 17.76 ;
      RECT MASK 1 20.738 17.279 20.798 17.76 ;
      RECT MASK 1 22.066 17.279 22.126 17.76 ;
      RECT MASK 1 22.398 17.279 22.458 17.76 ;
      RECT MASK 1 23.726 17.279 23.786 17.76 ;
      RECT MASK 1 24.058 17.279 24.118 17.76 ;
      RECT MASK 1 25.386 17.279 25.446 17.76 ;
      RECT MASK 1 25.718 17.279 25.778 17.76 ;
      RECT MASK 1 27.046 17.279 27.106 17.76 ;
      RECT MASK 1 27.378 17.279 27.438 17.76 ;
      RECT MASK 1 28.706 17.279 28.766 17.76 ;
      RECT MASK 1 29.038 17.279 29.098 17.76 ;
      RECT MASK 1 30.366 17.279 30.426 17.76 ;
      RECT MASK 1 30.698 17.279 30.758 17.76 ;
      RECT MASK 1 32.026 17.279 32.086 17.76 ;
      RECT MASK 1 32.358 17.279 32.418 17.76 ;
      RECT MASK 1 33.686 17.279 33.746 17.76 ;
      RECT MASK 1 34.018 17.279 34.078 17.76 ;
      RECT MASK 1 35.346 17.279 35.406 17.76 ;
      RECT MASK 1 35.678 17.279 35.738 17.76 ;
      RECT MASK 1 37.006 17.279 37.066 17.76 ;
      RECT MASK 1 37.338 17.279 37.398 17.76 ;
      RECT MASK 1 38.666 17.279 38.726 17.76 ;
      RECT MASK 1 38.998 17.279 39.058 17.76 ;
      RECT MASK 1 40.326 17.279 40.386 17.76 ;
      RECT MASK 1 40.658 17.279 40.718 17.76 ;
      RECT MASK 1 41.986 17.279 42.046 17.76 ;
      RECT MASK 1 42.318 17.279 42.378 17.76 ;
      RECT MASK 1 43.646 17.279 43.706 17.76 ;
      RECT MASK 1 43.978 17.279 44.038 17.76 ;
      RECT MASK 1 45.306 17.279 45.366 17.76 ;
      RECT MASK 1 45.638 17.279 45.698 17.76 ;
      RECT MASK 1 46.966 17.279 47.026 17.76 ;
      RECT MASK 1 47.298 17.279 47.358 17.76 ;
      RECT MASK 1 48.626 17.279 48.686 17.76 ;
      RECT MASK 1 48.958 17.279 49.018 17.76 ;
      RECT MASK 1 50.286 17.279 50.346 17.76 ;
      RECT MASK 1 50.618 17.279 50.678 17.76 ;
      RECT MASK 1 51.946 17.279 52.006 17.76 ;
      RECT MASK 1 52.278 17.279 52.338 17.76 ;
      RECT MASK 1 53.606 17.279 53.666 17.76 ;
      RECT MASK 1 53.938 17.279 53.998 17.76 ;
      RECT MASK 1 55.266 17.279 55.326 17.76 ;
      RECT MASK 1 55.598 17.279 55.658 17.76 ;
      RECT MASK 1 57.092 17.279 57.152 17.76 ;
      RECT MASK 1 57.424 17.279 57.484 17.76 ;
      RECT MASK 1 58.752 17.279 58.812 17.76 ;
      RECT MASK 1 59.084 17.279 59.144 17.76 ;
      RECT MASK 1 60.412 17.279 60.472 17.76 ;
      RECT MASK 1 60.744 17.279 60.804 17.76 ;
      RECT MASK 1 62.072 17.279 62.132 17.76 ;
      RECT MASK 1 62.404 17.279 62.464 17.76 ;
      RECT MASK 1 63.732 17.279 63.792 17.76 ;
      RECT MASK 1 64.064 17.279 64.124 17.76 ;
      RECT MASK 1 65.392 17.279 65.452 17.76 ;
      RECT MASK 1 65.724 17.279 65.784 17.76 ;
      RECT MASK 1 67.042 17.279 67.122 17.76 ;
      RECT MASK 1 67.374 17.279 67.454 17.76 ;
      RECT MASK 1 68.712 17.279 68.772 17.76 ;
      RECT MASK 1 69.044 17.279 69.104 17.76 ;
      RECT MASK 1 70.372 17.279 70.432 17.76 ;
      RECT MASK 1 70.704 17.279 70.764 17.76 ;
      RECT MASK 1 72.032 17.279 72.092 17.76 ;
      RECT MASK 1 72.364 17.279 72.424 17.76 ;
      RECT MASK 1 73.692 17.279 73.752 17.76 ;
      RECT MASK 1 74.024 17.279 74.084 17.76 ;
      RECT MASK 1 75.352 17.279 75.412 17.76 ;
      RECT MASK 1 75.684 17.279 75.744 17.76 ;
      RECT MASK 1 77.012 17.279 77.072 17.76 ;
      RECT MASK 1 77.344 17.279 77.404 17.76 ;
      RECT MASK 1 78.672 17.279 78.732 17.76 ;
      RECT MASK 1 79.004 17.279 79.064 17.76 ;
      RECT MASK 1 80.332 17.279 80.392 17.76 ;
      RECT MASK 1 80.664 17.279 80.724 17.76 ;
      RECT MASK 1 81.992 17.279 82.052 17.76 ;
      RECT MASK 1 82.324 17.279 82.384 17.76 ;
      RECT MASK 1 83.652 17.279 83.712 17.76 ;
      RECT MASK 1 83.984 17.279 84.044 17.76 ;
      RECT MASK 1 85.312 17.279 85.372 17.76 ;
      RECT MASK 1 85.644 17.279 85.704 17.76 ;
      RECT MASK 1 86.972 17.279 87.032 17.76 ;
      RECT MASK 1 87.304 17.279 87.364 17.76 ;
      RECT MASK 1 88.632 17.279 88.692 17.76 ;
      RECT MASK 1 88.964 17.279 89.024 17.76 ;
      RECT MASK 1 90.292 17.279 90.352 17.76 ;
      RECT MASK 1 90.624 17.279 90.684 17.76 ;
      RECT MASK 1 91.952 17.279 92.012 17.76 ;
      RECT MASK 1 92.284 17.279 92.344 17.76 ;
      RECT MASK 1 93.612 17.279 93.672 17.76 ;
      RECT MASK 1 93.944 17.279 94.004 17.76 ;
      RECT MASK 1 95.272 17.279 95.332 17.76 ;
      RECT MASK 1 95.604 17.279 95.664 17.76 ;
      RECT MASK 1 96.932 17.279 96.992 17.76 ;
      RECT MASK 1 97.264 17.279 97.324 17.76 ;
      RECT MASK 1 98.592 17.279 98.652 17.76 ;
      RECT MASK 1 98.924 17.279 98.984 17.76 ;
      RECT MASK 1 100.252 17.279 100.312 17.76 ;
      RECT MASK 1 100.584 17.279 100.644 17.76 ;
      RECT MASK 1 101.912 17.279 101.972 17.76 ;
      RECT MASK 1 102.244 17.279 102.304 17.76 ;
      RECT MASK 1 103.572 17.279 103.632 17.76 ;
      RECT MASK 1 103.904 17.279 103.964 17.76 ;
      RECT MASK 1 105.232 17.279 105.292 17.76 ;
      RECT MASK 1 105.564 17.279 105.624 17.76 ;
      RECT MASK 1 106.892 17.279 106.952 17.76 ;
      RECT MASK 1 107.224 17.279 107.284 17.76 ;
      RECT MASK 1 108.552 17.279 108.612 17.76 ;
      RECT MASK 1 108.884 17.279 108.944 17.76 ;
      RECT MASK 1 110.212 17.279 110.272 17.76 ;
      RECT MASK 1 110.544 17.279 110.604 17.76 ;
      RECT MASK 1 8.072 17.905 8.132 18.719 ;
      RECT MASK 1 8.404 17.905 8.464 18.473 ;
      RECT MASK 1 14.69 17.905 14.75 18.719 ;
      RECT MASK 1 15.022 17.905 15.082 18.473 ;
      RECT MASK 1 21.308 17.905 21.368 18.719 ;
      RECT MASK 1 21.64 17.905 21.7 18.473 ;
      RECT MASK 1 27.926 17.905 27.986 18.719 ;
      RECT MASK 1 28.258 17.905 28.318 18.473 ;
      RECT MASK 1 34.544 17.905 34.604 18.719 ;
      RECT MASK 1 34.876 17.905 34.936 18.473 ;
      RECT MASK 1 41.162 17.905 41.222 18.719 ;
      RECT MASK 1 41.494 17.905 41.554 18.473 ;
      RECT MASK 1 47.78 17.905 47.84 18.719 ;
      RECT MASK 1 48.112 17.905 48.172 18.473 ;
      RECT MASK 1 54.398 17.905 54.458 18.719 ;
      RECT MASK 1 54.73 17.905 54.79 18.473 ;
      RECT MASK 1 61.016 17.905 61.076 18.719 ;
      RECT MASK 1 61.348 17.905 61.408 18.473 ;
      RECT MASK 1 67.634 17.905 67.694 18.719 ;
      RECT MASK 1 67.966 17.905 68.026 18.473 ;
      RECT MASK 1 74.252 17.905 74.312 18.719 ;
      RECT MASK 1 74.584 17.905 74.644 18.473 ;
      RECT MASK 1 80.87 17.905 80.93 18.719 ;
      RECT MASK 1 81.202 17.905 81.262 18.473 ;
      RECT MASK 1 87.488 17.905 87.548 18.719 ;
      RECT MASK 1 87.82 17.905 87.88 18.473 ;
      RECT MASK 1 94.106 17.905 94.166 18.719 ;
      RECT MASK 1 94.438 17.905 94.498 18.473 ;
      RECT MASK 1 100.724 17.905 100.784 18.719 ;
      RECT MASK 1 101.056 17.905 101.116 18.473 ;
      RECT MASK 1 107.342 17.905 107.402 18.719 ;
      RECT MASK 1 107.674 17.905 107.734 18.473 ;
      RECT MASK 1 5.167 17.906 5.227 19.672 ;
      RECT MASK 1 5.4575 17.906 5.5175 18.474 ;
      RECT MASK 1 5.748 17.906 5.808 18.719 ;
      RECT MASK 1 6.08 17.906 6.14 18.474 ;
      RECT MASK 1 6.412 17.906 6.472 18.719 ;
      RECT MASK 1 6.6575 17.906 6.7175 18.474 ;
      RECT MASK 1 6.91 17.906 6.97 18.719 ;
      RECT MASK 1 7.242 17.906 7.302 18.474 ;
      RECT MASK 1 7.574 17.906 7.634 18.719 ;
      RECT MASK 1 8.736 17.906 8.796 18.719 ;
      RECT MASK 1 9.234 17.906 9.294 18.719 ;
      RECT MASK 1 9.566 17.906 9.626 18.474 ;
      RECT MASK 1 9.898 17.906 9.958 18.719 ;
      RECT MASK 1 10.23 17.906 10.29 18.474 ;
      RECT MASK 1 10.479 17.906 10.539 19.672 ;
      RECT MASK 1 11.785 17.906 11.845 19.672 ;
      RECT MASK 1 12.0755 17.906 12.1355 18.474 ;
      RECT MASK 1 12.366 17.906 12.426 18.719 ;
      RECT MASK 1 12.698 17.906 12.758 18.474 ;
      RECT MASK 1 13.03 17.906 13.09 18.719 ;
      RECT MASK 1 13.2755 17.906 13.3355 18.474 ;
      RECT MASK 1 13.528 17.906 13.588 18.719 ;
      RECT MASK 1 13.86 17.906 13.92 18.474 ;
      RECT MASK 1 14.192 17.906 14.252 18.719 ;
      RECT MASK 1 15.354 17.906 15.414 18.719 ;
      RECT MASK 1 15.852 17.906 15.912 18.719 ;
      RECT MASK 1 16.184 17.906 16.244 18.474 ;
      RECT MASK 1 16.516 17.906 16.576 18.719 ;
      RECT MASK 1 16.848 17.906 16.908 18.474 ;
      RECT MASK 1 17.097 17.906 17.157 19.672 ;
      RECT MASK 1 18.403 17.906 18.463 19.672 ;
      RECT MASK 1 18.6935 17.906 18.7535 18.474 ;
      RECT MASK 1 18.984 17.906 19.044 18.719 ;
      RECT MASK 1 19.316 17.906 19.376 18.474 ;
      RECT MASK 1 19.648 17.906 19.708 18.719 ;
      RECT MASK 1 19.8935 17.906 19.9535 18.474 ;
      RECT MASK 1 20.146 17.906 20.206 18.719 ;
      RECT MASK 1 20.478 17.906 20.538 18.474 ;
      RECT MASK 1 20.81 17.906 20.87 18.719 ;
      RECT MASK 1 21.972 17.906 22.032 18.719 ;
      RECT MASK 1 22.47 17.906 22.53 18.719 ;
      RECT MASK 1 22.802 17.906 22.862 18.474 ;
      RECT MASK 1 23.134 17.906 23.194 18.719 ;
      RECT MASK 1 23.466 17.906 23.526 18.474 ;
      RECT MASK 1 23.715 17.906 23.775 19.672 ;
      RECT MASK 1 25.021 17.906 25.081 19.672 ;
      RECT MASK 1 25.3115 17.906 25.3715 18.474 ;
      RECT MASK 1 25.602 17.906 25.662 18.719 ;
      RECT MASK 1 25.934 17.906 25.994 18.474 ;
      RECT MASK 1 26.266 17.906 26.326 18.719 ;
      RECT MASK 1 26.5115 17.906 26.5715 18.474 ;
      RECT MASK 1 26.764 17.906 26.824 18.719 ;
      RECT MASK 1 27.096 17.906 27.156 18.474 ;
      RECT MASK 1 27.428 17.906 27.488 18.719 ;
      RECT MASK 1 28.59 17.906 28.65 18.719 ;
      RECT MASK 1 29.088 17.906 29.148 18.719 ;
      RECT MASK 1 29.42 17.906 29.48 18.474 ;
      RECT MASK 1 29.752 17.906 29.812 18.719 ;
      RECT MASK 1 30.084 17.906 30.144 18.474 ;
      RECT MASK 1 30.333 17.906 30.393 19.672 ;
      RECT MASK 1 31.639 17.906 31.699 19.672 ;
      RECT MASK 1 31.9295 17.906 31.9895 18.474 ;
      RECT MASK 1 32.22 17.906 32.28 18.719 ;
      RECT MASK 1 32.552 17.906 32.612 18.474 ;
      RECT MASK 1 32.884 17.906 32.944 18.719 ;
      RECT MASK 1 33.1295 17.906 33.1895 18.474 ;
      RECT MASK 1 33.382 17.906 33.442 18.719 ;
      RECT MASK 1 33.714 17.906 33.774 18.474 ;
      RECT MASK 1 34.046 17.906 34.106 18.719 ;
      RECT MASK 1 35.208 17.906 35.268 18.719 ;
      RECT MASK 1 35.706 17.906 35.766 18.719 ;
      RECT MASK 1 36.038 17.906 36.098 18.474 ;
      RECT MASK 1 36.37 17.906 36.43 18.719 ;
      RECT MASK 1 36.702 17.906 36.762 18.474 ;
      RECT MASK 1 36.951 17.906 37.011 19.672 ;
      RECT MASK 1 38.257 17.906 38.317 19.672 ;
      RECT MASK 1 38.5475 17.906 38.6075 18.474 ;
      RECT MASK 1 38.838 17.906 38.898 18.719 ;
      RECT MASK 1 39.17 17.906 39.23 18.474 ;
      RECT MASK 1 39.502 17.906 39.562 18.719 ;
      RECT MASK 1 39.7475 17.906 39.8075 18.474 ;
      RECT MASK 1 40 17.906 40.06 18.719 ;
      RECT MASK 1 40.332 17.906 40.392 18.474 ;
      RECT MASK 1 40.664 17.906 40.724 18.719 ;
      RECT MASK 1 41.826 17.906 41.886 18.719 ;
      RECT MASK 1 42.324 17.906 42.384 18.719 ;
      RECT MASK 1 42.656 17.906 42.716 18.474 ;
      RECT MASK 1 42.988 17.906 43.048 18.719 ;
      RECT MASK 1 43.32 17.906 43.38 18.474 ;
      RECT MASK 1 43.569 17.906 43.629 19.672 ;
      RECT MASK 1 44.875 17.906 44.935 19.672 ;
      RECT MASK 1 45.1655 17.906 45.2255 18.474 ;
      RECT MASK 1 45.456 17.906 45.516 18.719 ;
      RECT MASK 1 45.788 17.906 45.848 18.474 ;
      RECT MASK 1 46.12 17.906 46.18 18.719 ;
      RECT MASK 1 46.3655 17.906 46.4255 18.474 ;
      RECT MASK 1 46.618 17.906 46.678 18.719 ;
      RECT MASK 1 46.95 17.906 47.01 18.474 ;
      RECT MASK 1 47.282 17.906 47.342 18.719 ;
      RECT MASK 1 48.444 17.906 48.504 18.719 ;
      RECT MASK 1 48.942 17.906 49.002 18.719 ;
      RECT MASK 1 49.274 17.906 49.334 18.474 ;
      RECT MASK 1 49.606 17.906 49.666 18.719 ;
      RECT MASK 1 49.938 17.906 49.998 18.474 ;
      RECT MASK 1 50.187 17.906 50.247 19.672 ;
      RECT MASK 1 51.493 17.906 51.553 19.672 ;
      RECT MASK 1 51.7835 17.906 51.8435 18.474 ;
      RECT MASK 1 52.074 17.906 52.134 18.719 ;
      RECT MASK 1 52.406 17.906 52.466 18.474 ;
      RECT MASK 1 52.738 17.906 52.798 18.719 ;
      RECT MASK 1 52.9835 17.906 53.0435 18.474 ;
      RECT MASK 1 53.236 17.906 53.296 18.719 ;
      RECT MASK 1 53.568 17.906 53.628 18.474 ;
      RECT MASK 1 53.9 17.906 53.96 18.719 ;
      RECT MASK 1 55.062 17.906 55.122 18.719 ;
      RECT MASK 1 55.56 17.906 55.62 18.719 ;
      RECT MASK 1 55.892 17.906 55.952 18.474 ;
      RECT MASK 1 56.224 17.906 56.284 18.719 ;
      RECT MASK 1 56.556 17.906 56.616 18.474 ;
      RECT MASK 1 56.805 17.906 56.865 19.672 ;
      RECT MASK 1 58.111 17.906 58.171 19.672 ;
      RECT MASK 1 58.4015 17.906 58.4615 18.474 ;
      RECT MASK 1 58.692 17.906 58.752 18.719 ;
      RECT MASK 1 59.024 17.906 59.084 18.474 ;
      RECT MASK 1 59.356 17.906 59.416 18.719 ;
      RECT MASK 1 59.6015 17.906 59.6615 18.474 ;
      RECT MASK 1 59.854 17.906 59.914 18.719 ;
      RECT MASK 1 60.186 17.906 60.246 18.474 ;
      RECT MASK 1 60.518 17.906 60.578 18.719 ;
      RECT MASK 1 61.68 17.906 61.74 18.719 ;
      RECT MASK 1 62.178 17.906 62.238 18.719 ;
      RECT MASK 1 62.51 17.906 62.57 18.474 ;
      RECT MASK 1 62.842 17.906 62.902 18.719 ;
      RECT MASK 1 63.174 17.906 63.234 18.474 ;
      RECT MASK 1 63.423 17.906 63.483 19.672 ;
      RECT MASK 1 64.729 17.906 64.789 19.672 ;
      RECT MASK 1 65.0195 17.906 65.0795 18.474 ;
      RECT MASK 1 65.31 17.906 65.37 18.719 ;
      RECT MASK 1 65.642 17.906 65.702 18.474 ;
      RECT MASK 1 65.974 17.906 66.034 18.719 ;
      RECT MASK 1 66.2195 17.906 66.2795 18.474 ;
      RECT MASK 1 66.472 17.906 66.532 18.719 ;
      RECT MASK 1 66.804 17.906 66.864 18.474 ;
      RECT MASK 1 67.136 17.906 67.196 18.719 ;
      RECT MASK 1 68.298 17.906 68.358 18.719 ;
      RECT MASK 1 68.796 17.906 68.856 18.719 ;
      RECT MASK 1 69.128 17.906 69.188 18.474 ;
      RECT MASK 1 69.46 17.906 69.52 18.719 ;
      RECT MASK 1 69.792 17.906 69.852 18.474 ;
      RECT MASK 1 70.041 17.906 70.101 19.672 ;
      RECT MASK 1 71.347 17.906 71.407 19.672 ;
      RECT MASK 1 71.6375 17.906 71.6975 18.474 ;
      RECT MASK 1 71.928 17.906 71.988 18.719 ;
      RECT MASK 1 72.26 17.906 72.32 18.474 ;
      RECT MASK 1 72.592 17.906 72.652 18.719 ;
      RECT MASK 1 72.8375 17.906 72.8975 18.474 ;
      RECT MASK 1 73.09 17.906 73.15 18.719 ;
      RECT MASK 1 73.422 17.906 73.482 18.474 ;
      RECT MASK 1 73.754 17.906 73.814 18.719 ;
      RECT MASK 1 74.916 17.906 74.976 18.719 ;
      RECT MASK 1 75.414 17.906 75.474 18.719 ;
      RECT MASK 1 75.746 17.906 75.806 18.474 ;
      RECT MASK 1 76.078 17.906 76.138 18.719 ;
      RECT MASK 1 76.41 17.906 76.47 18.474 ;
      RECT MASK 1 76.659 17.906 76.719 19.672 ;
      RECT MASK 1 77.965 17.906 78.025 19.672 ;
      RECT MASK 1 78.2555 17.906 78.3155 18.474 ;
      RECT MASK 1 78.546 17.906 78.606 18.719 ;
      RECT MASK 1 78.878 17.906 78.938 18.474 ;
      RECT MASK 1 79.21 17.906 79.27 18.719 ;
      RECT MASK 1 79.4555 17.906 79.5155 18.474 ;
      RECT MASK 1 79.708 17.906 79.768 18.719 ;
      RECT MASK 1 80.04 17.906 80.1 18.474 ;
      RECT MASK 1 80.372 17.906 80.432 18.719 ;
      RECT MASK 1 81.534 17.906 81.594 18.719 ;
      RECT MASK 1 82.032 17.906 82.092 18.719 ;
      RECT MASK 1 82.364 17.906 82.424 18.474 ;
      RECT MASK 1 82.696 17.906 82.756 18.719 ;
      RECT MASK 1 83.028 17.906 83.088 18.474 ;
      RECT MASK 1 83.277 17.906 83.337 19.672 ;
      RECT MASK 1 84.583 17.906 84.643 19.672 ;
      RECT MASK 1 84.8735 17.906 84.9335 18.474 ;
      RECT MASK 1 85.164 17.906 85.224 18.719 ;
      RECT MASK 1 85.496 17.906 85.556 18.474 ;
      RECT MASK 1 85.828 17.906 85.888 18.719 ;
      RECT MASK 1 86.0735 17.906 86.1335 18.474 ;
      RECT MASK 1 86.326 17.906 86.386 18.719 ;
      RECT MASK 1 86.658 17.906 86.718 18.474 ;
      RECT MASK 1 86.99 17.906 87.05 18.719 ;
      RECT MASK 1 88.152 17.906 88.212 18.719 ;
      RECT MASK 1 88.65 17.906 88.71 18.719 ;
      RECT MASK 1 88.982 17.906 89.042 18.474 ;
      RECT MASK 1 89.314 17.906 89.374 18.719 ;
      RECT MASK 1 89.646 17.906 89.706 18.474 ;
      RECT MASK 1 89.895 17.906 89.955 19.672 ;
      RECT MASK 1 91.201 17.906 91.261 19.672 ;
      RECT MASK 1 91.4915 17.906 91.5515 18.474 ;
      RECT MASK 1 91.782 17.906 91.842 18.719 ;
      RECT MASK 1 92.114 17.906 92.174 18.474 ;
      RECT MASK 1 92.446 17.906 92.506 18.719 ;
      RECT MASK 1 92.6915 17.906 92.7515 18.474 ;
      RECT MASK 1 92.944 17.906 93.004 18.719 ;
      RECT MASK 1 93.276 17.906 93.336 18.474 ;
      RECT MASK 1 93.608 17.906 93.668 18.719 ;
      RECT MASK 1 94.77 17.906 94.83 18.719 ;
      RECT MASK 1 95.268 17.906 95.328 18.719 ;
      RECT MASK 1 95.6 17.906 95.66 18.474 ;
      RECT MASK 1 95.932 17.906 95.992 18.719 ;
      RECT MASK 1 96.264 17.906 96.324 18.474 ;
      RECT MASK 1 96.513 17.906 96.573 19.672 ;
      RECT MASK 1 97.819 17.906 97.879 19.672 ;
      RECT MASK 1 98.1095 17.906 98.1695 18.474 ;
      RECT MASK 1 98.4 17.906 98.46 18.719 ;
      RECT MASK 1 98.732 17.906 98.792 18.474 ;
      RECT MASK 1 99.064 17.906 99.124 18.719 ;
      RECT MASK 1 99.3095 17.906 99.3695 18.474 ;
      RECT MASK 1 99.562 17.906 99.622 18.719 ;
      RECT MASK 1 99.894 17.906 99.954 18.474 ;
      RECT MASK 1 100.226 17.906 100.286 18.719 ;
      RECT MASK 1 101.388 17.906 101.448 18.719 ;
      RECT MASK 1 101.886 17.906 101.946 18.719 ;
      RECT MASK 1 102.218 17.906 102.278 18.474 ;
      RECT MASK 1 102.55 17.906 102.61 18.719 ;
      RECT MASK 1 102.882 17.906 102.942 18.474 ;
      RECT MASK 1 103.131 17.906 103.191 19.672 ;
      RECT MASK 1 104.437 17.906 104.497 19.672 ;
      RECT MASK 1 104.7275 17.906 104.7875 18.474 ;
      RECT MASK 1 105.018 17.906 105.078 18.719 ;
      RECT MASK 1 105.35 17.906 105.41 18.474 ;
      RECT MASK 1 105.682 17.906 105.742 18.719 ;
      RECT MASK 1 105.9275 17.906 105.9875 18.474 ;
      RECT MASK 1 106.18 17.906 106.24 18.719 ;
      RECT MASK 1 106.512 17.906 106.572 18.474 ;
      RECT MASK 1 106.844 17.906 106.904 18.719 ;
      RECT MASK 1 108.006 17.906 108.066 18.719 ;
      RECT MASK 1 108.504 17.906 108.564 18.719 ;
      RECT MASK 1 108.836 17.906 108.896 18.474 ;
      RECT MASK 1 109.168 17.906 109.228 18.719 ;
      RECT MASK 1 109.5 17.906 109.56 18.474 ;
      RECT MASK 1 109.749 17.906 109.809 19.672 ;
      RECT MASK 1 5.748 18.839 5.808 20.671 ;
      RECT MASK 1 6.412 18.839 6.472 20.671 ;
      RECT MASK 1 6.91 18.839 6.97 20.671 ;
      RECT MASK 1 7.574 18.839 7.634 20.671 ;
      RECT MASK 1 8.072 18.839 8.132 20.671 ;
      RECT MASK 1 8.736 18.839 8.796 20.671 ;
      RECT MASK 1 9.234 18.839 9.294 20.671 ;
      RECT MASK 1 9.898 18.839 9.958 20.671 ;
      RECT MASK 1 12.366 18.839 12.426 20.671 ;
      RECT MASK 1 13.03 18.839 13.09 20.671 ;
      RECT MASK 1 13.528 18.839 13.588 20.671 ;
      RECT MASK 1 14.192 18.839 14.252 20.671 ;
      RECT MASK 1 14.69 18.839 14.75 20.671 ;
      RECT MASK 1 15.354 18.839 15.414 20.671 ;
      RECT MASK 1 15.852 18.839 15.912 20.671 ;
      RECT MASK 1 16.516 18.839 16.576 20.671 ;
      RECT MASK 1 18.984 18.839 19.044 20.671 ;
      RECT MASK 1 19.648 18.839 19.708 20.671 ;
      RECT MASK 1 20.146 18.839 20.206 20.671 ;
      RECT MASK 1 20.81 18.839 20.87 20.671 ;
      RECT MASK 1 21.308 18.839 21.368 20.671 ;
      RECT MASK 1 21.972 18.839 22.032 20.671 ;
      RECT MASK 1 22.47 18.839 22.53 20.671 ;
      RECT MASK 1 23.134 18.839 23.194 20.671 ;
      RECT MASK 1 25.602 18.839 25.662 20.671 ;
      RECT MASK 1 26.266 18.839 26.326 20.671 ;
      RECT MASK 1 26.764 18.839 26.824 20.671 ;
      RECT MASK 1 27.428 18.839 27.488 20.671 ;
      RECT MASK 1 27.926 18.839 27.986 20.671 ;
      RECT MASK 1 28.59 18.839 28.65 20.671 ;
      RECT MASK 1 29.088 18.839 29.148 20.671 ;
      RECT MASK 1 29.752 18.839 29.812 20.671 ;
      RECT MASK 1 32.22 18.839 32.28 20.671 ;
      RECT MASK 1 32.884 18.839 32.944 20.671 ;
      RECT MASK 1 33.382 18.839 33.442 20.671 ;
      RECT MASK 1 34.046 18.839 34.106 20.671 ;
      RECT MASK 1 34.544 18.839 34.604 20.671 ;
      RECT MASK 1 35.208 18.839 35.268 20.671 ;
      RECT MASK 1 35.706 18.839 35.766 20.671 ;
      RECT MASK 1 36.37 18.839 36.43 20.671 ;
      RECT MASK 1 38.838 18.839 38.898 20.671 ;
      RECT MASK 1 39.502 18.839 39.562 20.671 ;
      RECT MASK 1 40 18.839 40.06 20.671 ;
      RECT MASK 1 40.664 18.839 40.724 20.671 ;
      RECT MASK 1 41.162 18.839 41.222 20.671 ;
      RECT MASK 1 41.826 18.839 41.886 20.671 ;
      RECT MASK 1 42.324 18.839 42.384 20.671 ;
      RECT MASK 1 42.988 18.839 43.048 20.671 ;
      RECT MASK 1 45.456 18.839 45.516 20.671 ;
      RECT MASK 1 46.12 18.839 46.18 20.671 ;
      RECT MASK 1 46.618 18.839 46.678 20.671 ;
      RECT MASK 1 47.282 18.839 47.342 20.671 ;
      RECT MASK 1 47.78 18.839 47.84 20.671 ;
      RECT MASK 1 48.444 18.839 48.504 20.671 ;
      RECT MASK 1 48.942 18.839 49.002 20.671 ;
      RECT MASK 1 49.606 18.839 49.666 20.671 ;
      RECT MASK 1 52.074 18.839 52.134 20.671 ;
      RECT MASK 1 52.738 18.839 52.798 20.671 ;
      RECT MASK 1 53.236 18.839 53.296 20.671 ;
      RECT MASK 1 53.9 18.839 53.96 20.671 ;
      RECT MASK 1 54.398 18.839 54.458 20.671 ;
      RECT MASK 1 55.062 18.839 55.122 20.671 ;
      RECT MASK 1 55.56 18.839 55.62 20.671 ;
      RECT MASK 1 56.224 18.839 56.284 20.671 ;
      RECT MASK 1 58.692 18.839 58.752 20.671 ;
      RECT MASK 1 59.356 18.839 59.416 20.671 ;
      RECT MASK 1 59.854 18.839 59.914 20.671 ;
      RECT MASK 1 60.518 18.839 60.578 20.671 ;
      RECT MASK 1 61.016 18.839 61.076 20.671 ;
      RECT MASK 1 61.68 18.839 61.74 20.671 ;
      RECT MASK 1 62.178 18.839 62.238 20.671 ;
      RECT MASK 1 62.842 18.839 62.902 20.671 ;
      RECT MASK 1 65.31 18.839 65.37 20.671 ;
      RECT MASK 1 65.974 18.839 66.034 20.671 ;
      RECT MASK 1 66.472 18.839 66.532 20.671 ;
      RECT MASK 1 67.136 18.839 67.196 20.671 ;
      RECT MASK 1 67.634 18.839 67.694 20.671 ;
      RECT MASK 1 68.298 18.839 68.358 20.671 ;
      RECT MASK 1 68.796 18.839 68.856 20.671 ;
      RECT MASK 1 69.46 18.839 69.52 20.671 ;
      RECT MASK 1 71.928 18.839 71.988 20.671 ;
      RECT MASK 1 72.592 18.839 72.652 20.671 ;
      RECT MASK 1 73.09 18.839 73.15 20.671 ;
      RECT MASK 1 73.754 18.839 73.814 20.671 ;
      RECT MASK 1 74.252 18.839 74.312 20.671 ;
      RECT MASK 1 74.916 18.839 74.976 20.671 ;
      RECT MASK 1 75.414 18.839 75.474 20.671 ;
      RECT MASK 1 76.078 18.839 76.138 20.671 ;
      RECT MASK 1 78.546 18.839 78.606 20.671 ;
      RECT MASK 1 79.21 18.839 79.27 20.671 ;
      RECT MASK 1 79.708 18.839 79.768 20.671 ;
      RECT MASK 1 80.372 18.839 80.432 20.671 ;
      RECT MASK 1 80.87 18.839 80.93 20.671 ;
      RECT MASK 1 81.534 18.839 81.594 20.671 ;
      RECT MASK 1 82.032 18.839 82.092 20.671 ;
      RECT MASK 1 82.696 18.839 82.756 20.671 ;
      RECT MASK 1 85.164 18.839 85.224 20.671 ;
      RECT MASK 1 85.828 18.839 85.888 20.671 ;
      RECT MASK 1 86.326 18.839 86.386 20.671 ;
      RECT MASK 1 86.99 18.839 87.05 20.671 ;
      RECT MASK 1 87.488 18.839 87.548 20.671 ;
      RECT MASK 1 88.152 18.839 88.212 20.671 ;
      RECT MASK 1 88.65 18.839 88.71 20.671 ;
      RECT MASK 1 89.314 18.839 89.374 20.671 ;
      RECT MASK 1 91.782 18.839 91.842 20.671 ;
      RECT MASK 1 92.446 18.839 92.506 20.671 ;
      RECT MASK 1 92.944 18.839 93.004 20.671 ;
      RECT MASK 1 93.608 18.839 93.668 20.671 ;
      RECT MASK 1 94.106 18.839 94.166 20.671 ;
      RECT MASK 1 94.77 18.839 94.83 20.671 ;
      RECT MASK 1 95.268 18.839 95.328 20.671 ;
      RECT MASK 1 95.932 18.839 95.992 20.671 ;
      RECT MASK 1 98.4 18.839 98.46 20.671 ;
      RECT MASK 1 99.064 18.839 99.124 20.671 ;
      RECT MASK 1 99.562 18.839 99.622 20.671 ;
      RECT MASK 1 100.226 18.839 100.286 20.671 ;
      RECT MASK 1 100.724 18.839 100.784 20.671 ;
      RECT MASK 1 101.388 18.839 101.448 20.671 ;
      RECT MASK 1 101.886 18.839 101.946 20.671 ;
      RECT MASK 1 102.55 18.839 102.61 20.671 ;
      RECT MASK 1 105.018 18.839 105.078 20.671 ;
      RECT MASK 1 105.682 18.839 105.742 20.671 ;
      RECT MASK 1 106.18 18.839 106.24 20.671 ;
      RECT MASK 1 106.844 18.839 106.904 20.671 ;
      RECT MASK 1 107.342 18.839 107.402 20.671 ;
      RECT MASK 1 108.006 18.839 108.066 20.671 ;
      RECT MASK 1 108.504 18.839 108.564 20.671 ;
      RECT MASK 1 109.168 18.839 109.228 20.671 ;
      RECT MASK 1 1.421 18.95 1.521 24.951 ;
      RECT MASK 1 4.575 18.95 4.675 24.951 ;
      RECT MASK 1 2.225 19.56 2.285 24.422 ;
      RECT MASK 1 2.499 19.56 2.559 24.53 ;
      RECT MASK 1 2.773 19.56 2.833 24.53 ;
      RECT MASK 1 3.047 19.56 3.107 24.53 ;
      RECT MASK 1 3.321 19.56 3.381 24.53 ;
      RECT MASK 1 3.595 19.56 3.655 24.53 ;
      RECT MASK 1 3.869 19.56 3.929 24.422 ;
      RECT MASK 1 58.111 19.798 58.171 23.55 ;
      RECT MASK 1 5.167 19.816 5.227 23.545 ;
      RECT MASK 1 10.479 19.816 10.539 21.21 ;
      RECT MASK 1 11.785 19.816 11.845 21.21 ;
      RECT MASK 1 17.097 19.816 17.157 21.21 ;
      RECT MASK 1 18.403 19.816 18.463 21.21 ;
      RECT MASK 1 23.715 19.816 23.775 21.21 ;
      RECT MASK 1 25.021 19.816 25.081 21.21 ;
      RECT MASK 1 30.333 19.816 30.393 21.21 ;
      RECT MASK 1 31.639 19.816 31.699 21.21 ;
      RECT MASK 1 36.951 19.816 37.011 21.21 ;
      RECT MASK 1 38.257 19.816 38.317 21.21 ;
      RECT MASK 1 43.569 19.816 43.629 21.21 ;
      RECT MASK 1 44.875 19.816 44.935 21.21 ;
      RECT MASK 1 50.187 19.816 50.247 21.21 ;
      RECT MASK 1 51.493 19.816 51.553 21.21 ;
      RECT MASK 1 56.805 19.816 56.865 23.545 ;
      RECT MASK 1 63.423 19.816 63.483 21.21 ;
      RECT MASK 1 64.729 19.816 64.789 21.21 ;
      RECT MASK 1 70.041 19.816 70.101 21.21 ;
      RECT MASK 1 71.347 19.816 71.407 21.21 ;
      RECT MASK 1 76.659 19.816 76.719 21.21 ;
      RECT MASK 1 77.965 19.816 78.025 21.21 ;
      RECT MASK 1 83.277 19.816 83.337 21.21 ;
      RECT MASK 1 84.583 19.816 84.643 21.21 ;
      RECT MASK 1 89.895 19.816 89.955 21.21 ;
      RECT MASK 1 91.201 19.816 91.261 21.21 ;
      RECT MASK 1 96.513 19.816 96.573 21.21 ;
      RECT MASK 1 97.819 19.816 97.879 21.21 ;
      RECT MASK 1 103.131 19.816 103.191 21.21 ;
      RECT MASK 1 104.437 19.816 104.497 21.21 ;
      RECT MASK 1 109.749 19.816 109.809 21.21 ;
      RECT MASK 1 57.225 20.387 57.285 21.9635 ;
      RECT MASK 1 57.557 20.387 57.617 21.9635 ;
      RECT MASK 1 57.889 20.387 57.949 21.9635 ;
      RECT MASK 1 58.277 20.387 58.337 21.9635 ;
      RECT MASK 1 59.024 20.7735 59.084 21.6 ;
      RECT MASK 1 5.748 20.791 5.808 21.085 ;
      RECT MASK 1 6.412 20.791 6.472 21.085 ;
      RECT MASK 1 6.91 20.791 6.97 21.085 ;
      RECT MASK 1 7.574 20.791 7.634 21.085 ;
      RECT MASK 1 8.072 20.791 8.132 21.085 ;
      RECT MASK 1 8.736 20.791 8.796 21.085 ;
      RECT MASK 1 9.234 20.791 9.294 21.085 ;
      RECT MASK 1 9.898 20.791 9.958 21.085 ;
      RECT MASK 1 12.366 20.791 12.426 21.085 ;
      RECT MASK 1 13.03 20.791 13.09 21.085 ;
      RECT MASK 1 13.528 20.791 13.588 21.085 ;
      RECT MASK 1 14.192 20.791 14.252 21.085 ;
      RECT MASK 1 14.69 20.791 14.75 21.085 ;
      RECT MASK 1 15.354 20.791 15.414 21.085 ;
      RECT MASK 1 15.852 20.791 15.912 21.085 ;
      RECT MASK 1 16.516 20.791 16.576 21.085 ;
      RECT MASK 1 18.984 20.791 19.044 21.085 ;
      RECT MASK 1 19.648 20.791 19.708 21.085 ;
      RECT MASK 1 20.146 20.791 20.206 21.085 ;
      RECT MASK 1 20.81 20.791 20.87 21.085 ;
      RECT MASK 1 21.308 20.791 21.368 21.085 ;
      RECT MASK 1 21.972 20.791 22.032 21.085 ;
      RECT MASK 1 22.47 20.791 22.53 21.085 ;
      RECT MASK 1 23.134 20.791 23.194 21.085 ;
      RECT MASK 1 25.602 20.791 25.662 21.085 ;
      RECT MASK 1 26.266 20.791 26.326 21.085 ;
      RECT MASK 1 26.764 20.791 26.824 21.085 ;
      RECT MASK 1 27.428 20.791 27.488 21.085 ;
      RECT MASK 1 27.926 20.791 27.986 21.085 ;
      RECT MASK 1 28.59 20.791 28.65 21.085 ;
      RECT MASK 1 29.088 20.791 29.148 21.085 ;
      RECT MASK 1 29.752 20.791 29.812 21.085 ;
      RECT MASK 1 32.22 20.791 32.28 21.085 ;
      RECT MASK 1 32.884 20.791 32.944 21.085 ;
      RECT MASK 1 33.382 20.791 33.442 21.085 ;
      RECT MASK 1 34.046 20.791 34.106 21.085 ;
      RECT MASK 1 34.544 20.791 34.604 21.085 ;
      RECT MASK 1 35.208 20.791 35.268 21.085 ;
      RECT MASK 1 35.706 20.791 35.766 21.085 ;
      RECT MASK 1 36.37 20.791 36.43 21.085 ;
      RECT MASK 1 38.838 20.791 38.898 21.085 ;
      RECT MASK 1 39.502 20.791 39.562 21.085 ;
      RECT MASK 1 40 20.791 40.06 21.085 ;
      RECT MASK 1 40.664 20.791 40.724 21.085 ;
      RECT MASK 1 41.162 20.791 41.222 21.085 ;
      RECT MASK 1 41.826 20.791 41.886 21.085 ;
      RECT MASK 1 42.324 20.791 42.384 21.085 ;
      RECT MASK 1 42.988 20.791 43.048 21.085 ;
      RECT MASK 1 45.456 20.791 45.516 21.085 ;
      RECT MASK 1 46.12 20.791 46.18 21.085 ;
      RECT MASK 1 46.618 20.791 46.678 21.085 ;
      RECT MASK 1 47.282 20.791 47.342 21.085 ;
      RECT MASK 1 47.78 20.791 47.84 21.085 ;
      RECT MASK 1 48.444 20.791 48.504 21.085 ;
      RECT MASK 1 48.942 20.791 49.002 21.085 ;
      RECT MASK 1 49.606 20.791 49.666 21.085 ;
      RECT MASK 1 52.074 20.791 52.134 21.085 ;
      RECT MASK 1 52.738 20.791 52.798 21.085 ;
      RECT MASK 1 53.236 20.791 53.296 21.085 ;
      RECT MASK 1 53.9 20.791 53.96 21.085 ;
      RECT MASK 1 54.398 20.791 54.458 21.085 ;
      RECT MASK 1 55.062 20.791 55.122 21.085 ;
      RECT MASK 1 55.56 20.791 55.62 21.085 ;
      RECT MASK 1 56.224 20.791 56.284 21.085 ;
      RECT MASK 1 58.692 20.791 58.752 21.085 ;
      RECT MASK 1 59.356 20.791 59.416 21.085 ;
      RECT MASK 1 59.854 20.791 59.914 21.085 ;
      RECT MASK 1 60.518 20.791 60.578 21.085 ;
      RECT MASK 1 61.016 20.791 61.076 21.085 ;
      RECT MASK 1 61.68 20.791 61.74 21.085 ;
      RECT MASK 1 62.178 20.791 62.238 21.085 ;
      RECT MASK 1 62.842 20.791 62.902 21.085 ;
      RECT MASK 1 65.31 20.791 65.37 21.085 ;
      RECT MASK 1 65.974 20.791 66.034 21.085 ;
      RECT MASK 1 66.472 20.791 66.532 21.085 ;
      RECT MASK 1 67.136 20.791 67.196 21.085 ;
      RECT MASK 1 67.634 20.791 67.694 21.085 ;
      RECT MASK 1 68.298 20.791 68.358 21.085 ;
      RECT MASK 1 68.796 20.791 68.856 21.085 ;
      RECT MASK 1 69.46 20.791 69.52 21.085 ;
      RECT MASK 1 71.928 20.791 71.988 21.085 ;
      RECT MASK 1 72.592 20.791 72.652 21.085 ;
      RECT MASK 1 73.09 20.791 73.15 21.085 ;
      RECT MASK 1 73.754 20.791 73.814 21.085 ;
      RECT MASK 1 74.252 20.791 74.312 21.085 ;
      RECT MASK 1 74.916 20.791 74.976 21.085 ;
      RECT MASK 1 75.414 20.791 75.474 21.085 ;
      RECT MASK 1 76.078 20.791 76.138 21.085 ;
      RECT MASK 1 78.546 20.791 78.606 21.085 ;
      RECT MASK 1 79.21 20.791 79.27 21.085 ;
      RECT MASK 1 79.708 20.791 79.768 21.085 ;
      RECT MASK 1 80.372 20.791 80.432 21.085 ;
      RECT MASK 1 80.87 20.791 80.93 21.085 ;
      RECT MASK 1 81.534 20.791 81.594 21.085 ;
      RECT MASK 1 82.032 20.791 82.092 21.085 ;
      RECT MASK 1 82.696 20.791 82.756 21.085 ;
      RECT MASK 1 85.164 20.791 85.224 21.085 ;
      RECT MASK 1 85.828 20.791 85.888 21.085 ;
      RECT MASK 1 86.326 20.791 86.386 21.085 ;
      RECT MASK 1 86.99 20.791 87.05 21.085 ;
      RECT MASK 1 87.488 20.791 87.548 21.085 ;
      RECT MASK 1 88.152 20.791 88.212 21.085 ;
      RECT MASK 1 88.65 20.791 88.71 21.085 ;
      RECT MASK 1 89.314 20.791 89.374 21.085 ;
      RECT MASK 1 91.782 20.791 91.842 21.085 ;
      RECT MASK 1 92.446 20.791 92.506 21.085 ;
      RECT MASK 1 92.944 20.791 93.004 21.085 ;
      RECT MASK 1 93.608 20.791 93.668 21.085 ;
      RECT MASK 1 94.106 20.791 94.166 21.085 ;
      RECT MASK 1 94.77 20.791 94.83 21.085 ;
      RECT MASK 1 95.268 20.791 95.328 21.085 ;
      RECT MASK 1 95.932 20.791 95.992 21.085 ;
      RECT MASK 1 98.4 20.791 98.46 21.085 ;
      RECT MASK 1 99.064 20.791 99.124 21.085 ;
      RECT MASK 1 99.562 20.791 99.622 21.085 ;
      RECT MASK 1 100.226 20.791 100.286 21.085 ;
      RECT MASK 1 100.724 20.791 100.784 21.085 ;
      RECT MASK 1 101.388 20.791 101.448 21.085 ;
      RECT MASK 1 101.886 20.791 101.946 21.085 ;
      RECT MASK 1 102.55 20.791 102.61 21.085 ;
      RECT MASK 1 105.018 20.791 105.078 21.085 ;
      RECT MASK 1 105.682 20.791 105.742 21.085 ;
      RECT MASK 1 106.18 20.791 106.24 21.085 ;
      RECT MASK 1 106.844 20.791 106.904 21.085 ;
      RECT MASK 1 107.342 20.791 107.402 21.085 ;
      RECT MASK 1 108.006 20.791 108.066 21.085 ;
      RECT MASK 1 108.504 20.791 108.564 21.085 ;
      RECT MASK 1 109.168 20.791 109.228 21.085 ;
      RECT MASK 1 103.645 21.064 103.705 22.61 ;
      RECT MASK 1 5.665 21.33 5.725 21.6 ;
      RECT MASK 1 6.827 21.33 6.887 21.6 ;
      RECT MASK 1 7.989 21.33 8.049 21.6 ;
      RECT MASK 1 9.151 21.33 9.211 21.6 ;
      RECT MASK 1 12.283 21.33 12.343 21.6 ;
      RECT MASK 1 13.445 21.33 13.505 21.6 ;
      RECT MASK 1 14.607 21.33 14.667 21.6 ;
      RECT MASK 1 15.769 21.33 15.829 21.6 ;
      RECT MASK 1 18.901 21.33 18.961 21.6 ;
      RECT MASK 1 20.063 21.33 20.123 21.6 ;
      RECT MASK 1 21.225 21.33 21.285 21.6 ;
      RECT MASK 1 22.387 21.33 22.447 21.6 ;
      RECT MASK 1 25.519 21.33 25.579 21.6 ;
      RECT MASK 1 26.681 21.33 26.741 21.6 ;
      RECT MASK 1 27.843 21.33 27.903 21.6 ;
      RECT MASK 1 29.005 21.33 29.065 21.6 ;
      RECT MASK 1 32.137 21.33 32.197 21.6 ;
      RECT MASK 1 33.299 21.33 33.359 21.6 ;
      RECT MASK 1 34.461 21.33 34.521 21.6 ;
      RECT MASK 1 35.623 21.33 35.683 21.6 ;
      RECT MASK 1 38.755 21.33 38.815 21.6 ;
      RECT MASK 1 39.917 21.33 39.977 21.6 ;
      RECT MASK 1 41.079 21.33 41.139 21.6 ;
      RECT MASK 1 42.241 21.33 42.301 21.6 ;
      RECT MASK 1 45.373 21.33 45.433 21.6 ;
      RECT MASK 1 46.535 21.33 46.595 21.6 ;
      RECT MASK 1 47.697 21.33 47.757 21.6 ;
      RECT MASK 1 48.859 21.33 48.919 21.6 ;
      RECT MASK 1 51.991 21.33 52.051 21.6 ;
      RECT MASK 1 53.153 21.33 53.213 21.6 ;
      RECT MASK 1 54.315 21.33 54.375 21.6 ;
      RECT MASK 1 55.477 21.33 55.537 21.6 ;
      RECT MASK 1 58.609 21.33 58.669 21.9635 ;
      RECT MASK 1 58.753 21.33 58.793 21.9635 ;
      RECT MASK 1 59.771 21.33 59.831 21.6 ;
      RECT MASK 1 60.933 21.33 60.993 21.6 ;
      RECT MASK 1 62.095 21.33 62.155 21.6 ;
      RECT MASK 1 65.227 21.33 65.287 21.6 ;
      RECT MASK 1 66.389 21.33 66.449 21.6 ;
      RECT MASK 1 67.551 21.33 67.611 21.6 ;
      RECT MASK 1 68.713 21.33 68.773 21.6 ;
      RECT MASK 1 71.845 21.33 71.905 21.6 ;
      RECT MASK 1 73.007 21.33 73.067 21.6 ;
      RECT MASK 1 74.169 21.33 74.229 21.6 ;
      RECT MASK 1 75.331 21.33 75.391 21.6 ;
      RECT MASK 1 78.463 21.33 78.523 21.6 ;
      RECT MASK 1 79.625 21.33 79.685 21.6 ;
      RECT MASK 1 80.787 21.33 80.847 21.6 ;
      RECT MASK 1 81.949 21.33 82.009 21.6 ;
      RECT MASK 1 85.081 21.33 85.141 21.6 ;
      RECT MASK 1 86.243 21.33 86.303 21.6 ;
      RECT MASK 1 87.405 21.33 87.465 21.6 ;
      RECT MASK 1 88.567 21.33 88.627 21.6 ;
      RECT MASK 1 91.699 21.33 91.759 21.6 ;
      RECT MASK 1 92.861 21.33 92.921 21.6 ;
      RECT MASK 1 94.023 21.33 94.083 21.6 ;
      RECT MASK 1 95.185 21.33 95.245 21.6 ;
      RECT MASK 1 98.317 21.33 98.377 21.6 ;
      RECT MASK 1 99.479 21.33 99.539 21.6 ;
      RECT MASK 1 100.641 21.33 100.701 21.6 ;
      RECT MASK 1 101.803 21.33 101.863 21.6 ;
      RECT MASK 1 104.935 21.33 104.995 21.6 ;
      RECT MASK 1 106.097 21.33 106.157 21.6 ;
      RECT MASK 1 107.259 21.33 107.319 21.6 ;
      RECT MASK 1 108.421 21.33 108.481 21.6 ;
      RECT MASK 1 10.479 21.335 10.539 23.545 ;
      RECT MASK 1 11.785 21.335 11.845 23.545 ;
      RECT MASK 1 23.715 21.335 23.775 23.545 ;
      RECT MASK 1 25.021 21.335 25.081 23.545 ;
      RECT MASK 1 30.333 21.335 30.393 23.545 ;
      RECT MASK 1 31.639 21.335 31.699 23.545 ;
      RECT MASK 1 36.951 21.335 37.011 23.545 ;
      RECT MASK 1 38.257 21.335 38.317 23.545 ;
      RECT MASK 1 43.569 21.335 43.629 23.545 ;
      RECT MASK 1 44.875 21.335 44.935 23.545 ;
      RECT MASK 1 50.187 21.335 50.247 23.545 ;
      RECT MASK 1 51.493 21.335 51.553 23.545 ;
      RECT MASK 1 63.423 21.335 63.483 23.545 ;
      RECT MASK 1 64.729 21.335 64.789 23.545 ;
      RECT MASK 1 70.041 21.335 70.101 23.545 ;
      RECT MASK 1 71.347 21.335 71.407 23.545 ;
      RECT MASK 1 76.659 21.335 76.719 23.545 ;
      RECT MASK 1 77.965 21.335 78.025 23.545 ;
      RECT MASK 1 83.277 21.335 83.337 23.545 ;
      RECT MASK 1 84.583 21.335 84.643 23.545 ;
      RECT MASK 1 89.895 21.335 89.955 23.545 ;
      RECT MASK 1 91.201 21.335 91.261 23.545 ;
      RECT MASK 1 96.513 21.335 96.573 23.545 ;
      RECT MASK 1 97.819 21.335 97.879 23.545 ;
      RECT MASK 1 103.131 21.335 103.191 23.545 ;
      RECT MASK 1 104.437 21.335 104.497 23.545 ;
      RECT MASK 1 109.749 21.335 109.809 23.545 ;
      RECT MASK 1 6.495 21.64 6.555 24.999 ;
      RECT MASK 1 7.657 21.64 7.717 24.999 ;
      RECT MASK 1 8.819 21.64 8.879 24.999 ;
      RECT MASK 1 9.981 21.64 10.041 24.999 ;
      RECT MASK 1 13.113 21.64 13.173 24.999 ;
      RECT MASK 1 14.275 21.64 14.335 24.999 ;
      RECT MASK 1 15.437 21.64 15.497 24.999 ;
      RECT MASK 1 16.599 21.64 16.659 24.999 ;
      RECT MASK 1 19.731 21.64 19.791 24.999 ;
      RECT MASK 1 20.893 21.64 20.953 24.999 ;
      RECT MASK 1 22.055 21.64 22.115 24.999 ;
      RECT MASK 1 23.217 21.64 23.277 24.999 ;
      RECT MASK 1 26.349 21.64 26.409 24.999 ;
      RECT MASK 1 27.511 21.64 27.571 24.999 ;
      RECT MASK 1 28.673 21.64 28.733 24.999 ;
      RECT MASK 1 29.835 21.64 29.895 24.999 ;
      RECT MASK 1 32.967 21.64 33.027 24.999 ;
      RECT MASK 1 34.129 21.64 34.189 24.999 ;
      RECT MASK 1 35.291 21.64 35.351 24.999 ;
      RECT MASK 1 36.453 21.64 36.513 24.999 ;
      RECT MASK 1 39.585 21.64 39.645 24.999 ;
      RECT MASK 1 40.747 21.64 40.807 24.999 ;
      RECT MASK 1 41.909 21.64 41.969 24.999 ;
      RECT MASK 1 43.071 21.64 43.131 24.999 ;
      RECT MASK 1 46.203 21.64 46.263 24.999 ;
      RECT MASK 1 47.365 21.64 47.425 24.999 ;
      RECT MASK 1 48.527 21.64 48.587 24.999 ;
      RECT MASK 1 49.689 21.64 49.749 24.999 ;
      RECT MASK 1 52.821 21.64 52.881 24.999 ;
      RECT MASK 1 53.983 21.64 54.043 24.999 ;
      RECT MASK 1 55.145 21.64 55.205 24.999 ;
      RECT MASK 1 56.307 21.64 56.367 24.999 ;
      RECT MASK 1 59.439 21.64 59.499 24.999 ;
      RECT MASK 1 60.601 21.64 60.661 24.999 ;
      RECT MASK 1 61.763 21.64 61.823 24.999 ;
      RECT MASK 1 62.925 21.64 62.985 24.999 ;
      RECT MASK 1 66.057 21.64 66.117 24.999 ;
      RECT MASK 1 67.219 21.64 67.279 24.999 ;
      RECT MASK 1 68.381 21.64 68.441 24.999 ;
      RECT MASK 1 69.543 21.64 69.603 24.999 ;
      RECT MASK 1 72.675 21.64 72.735 24.999 ;
      RECT MASK 1 73.837 21.64 73.897 24.999 ;
      RECT MASK 1 74.999 21.64 75.059 24.999 ;
      RECT MASK 1 76.161 21.64 76.221 24.999 ;
      RECT MASK 1 79.293 21.64 79.353 24.999 ;
      RECT MASK 1 80.455 21.64 80.515 24.999 ;
      RECT MASK 1 81.617 21.64 81.677 24.999 ;
      RECT MASK 1 82.779 21.64 82.839 24.999 ;
      RECT MASK 1 85.911 21.64 85.971 24.999 ;
      RECT MASK 1 87.073 21.64 87.133 24.999 ;
      RECT MASK 1 88.235 21.64 88.295 24.999 ;
      RECT MASK 1 89.397 21.64 89.457 24.999 ;
      RECT MASK 1 92.529 21.64 92.589 24.999 ;
      RECT MASK 1 93.691 21.64 93.751 24.999 ;
      RECT MASK 1 94.853 21.64 94.913 24.999 ;
      RECT MASK 1 96.015 21.64 96.075 24.999 ;
      RECT MASK 1 99.147 21.64 99.207 24.999 ;
      RECT MASK 1 100.309 21.64 100.369 24.999 ;
      RECT MASK 1 101.471 21.64 101.531 24.999 ;
      RECT MASK 1 102.633 21.64 102.693 24.999 ;
      RECT MASK 1 105.765 21.64 105.825 24.999 ;
      RECT MASK 1 106.927 21.64 106.987 24.999 ;
      RECT MASK 1 108.089 21.64 108.149 24.999 ;
      RECT MASK 1 109.251 21.64 109.311 24.999 ;
      RECT MASK 1 5.821 22.0915 5.901 25.394 ;
      RECT MASK 1 6.153 22.0915 6.233 25.394 ;
      RECT MASK 1 6.983 22.0915 7.063 25.394 ;
      RECT MASK 1 7.315 22.0915 7.395 25.394 ;
      RECT MASK 1 8.145 22.0915 8.225 25.394 ;
      RECT MASK 1 8.477 22.0915 8.557 25.394 ;
      RECT MASK 1 9.307 22.0915 9.387 25.394 ;
      RECT MASK 1 9.639 22.0915 9.719 25.394 ;
      RECT MASK 1 12.439 22.0915 12.519 25.394 ;
      RECT MASK 1 12.771 22.0915 12.851 25.394 ;
      RECT MASK 1 13.601 22.0915 13.681 25.394 ;
      RECT MASK 1 13.933 22.0915 14.013 25.394 ;
      RECT MASK 1 14.763 22.0915 14.843 25.394 ;
      RECT MASK 1 15.095 22.0915 15.175 25.394 ;
      RECT MASK 1 15.925 22.0915 16.005 25.394 ;
      RECT MASK 1 16.257 22.0915 16.337 25.394 ;
      RECT MASK 1 19.057 22.0915 19.137 25.394 ;
      RECT MASK 1 19.389 22.0915 19.469 25.394 ;
      RECT MASK 1 20.219 22.0915 20.299 25.394 ;
      RECT MASK 1 20.551 22.0915 20.631 25.394 ;
      RECT MASK 1 21.381 22.0915 21.461 25.394 ;
      RECT MASK 1 21.713 22.0915 21.793 25.394 ;
      RECT MASK 1 22.543 22.0915 22.623 25.394 ;
      RECT MASK 1 22.875 22.0915 22.955 25.394 ;
      RECT MASK 1 25.675 22.0915 25.755 25.394 ;
      RECT MASK 1 26.007 22.0915 26.087 25.394 ;
      RECT MASK 1 26.837 22.0915 26.917 25.394 ;
      RECT MASK 1 27.169 22.0915 27.249 25.394 ;
      RECT MASK 1 27.999 22.0915 28.079 25.394 ;
      RECT MASK 1 28.331 22.0915 28.411 25.394 ;
      RECT MASK 1 29.161 22.0915 29.241 25.394 ;
      RECT MASK 1 29.493 22.0915 29.573 25.394 ;
      RECT MASK 1 32.293 22.0915 32.373 25.394 ;
      RECT MASK 1 32.625 22.0915 32.705 25.394 ;
      RECT MASK 1 33.455 22.0915 33.535 25.394 ;
      RECT MASK 1 33.787 22.0915 33.867 25.394 ;
      RECT MASK 1 34.617 22.0915 34.697 25.394 ;
      RECT MASK 1 34.949 22.0915 35.029 25.394 ;
      RECT MASK 1 35.779 22.0915 35.859 25.394 ;
      RECT MASK 1 36.111 22.0915 36.191 25.394 ;
      RECT MASK 1 38.911 22.0915 38.991 25.394 ;
      RECT MASK 1 39.243 22.0915 39.323 25.394 ;
      RECT MASK 1 40.073 22.0915 40.153 25.394 ;
      RECT MASK 1 40.405 22.0915 40.485 25.394 ;
      RECT MASK 1 41.235 22.0915 41.315 25.394 ;
      RECT MASK 1 41.567 22.0915 41.647 25.394 ;
      RECT MASK 1 42.397 22.0915 42.477 25.394 ;
      RECT MASK 1 42.729 22.0915 42.809 25.394 ;
      RECT MASK 1 45.529 22.0915 45.609 25.394 ;
      RECT MASK 1 45.861 22.0915 45.941 25.394 ;
      RECT MASK 1 46.691 22.0915 46.771 25.394 ;
      RECT MASK 1 47.023 22.0915 47.103 25.394 ;
      RECT MASK 1 47.853 22.0915 47.933 25.394 ;
      RECT MASK 1 48.185 22.0915 48.265 25.394 ;
      RECT MASK 1 49.015 22.0915 49.095 25.394 ;
      RECT MASK 1 49.347 22.0915 49.427 25.394 ;
      RECT MASK 1 52.147 22.0915 52.227 25.394 ;
      RECT MASK 1 52.479 22.0915 52.559 25.394 ;
      RECT MASK 1 53.309 22.0915 53.389 25.394 ;
      RECT MASK 1 53.641 22.0915 53.721 25.394 ;
      RECT MASK 1 54.471 22.0915 54.551 25.394 ;
      RECT MASK 1 54.803 22.0915 54.883 25.394 ;
      RECT MASK 1 55.633 22.0915 55.713 25.394 ;
      RECT MASK 1 55.965 22.0915 56.045 25.394 ;
      RECT MASK 1 58.765 22.0915 58.845 25.394 ;
      RECT MASK 1 59.097 22.0915 59.177 25.394 ;
      RECT MASK 1 59.927 22.0915 60.007 25.394 ;
      RECT MASK 1 60.259 22.0915 60.339 25.394 ;
      RECT MASK 1 61.089 22.0915 61.169 25.394 ;
      RECT MASK 1 61.421 22.0915 61.501 25.394 ;
      RECT MASK 1 62.251 22.0915 62.331 25.394 ;
      RECT MASK 1 62.583 22.0915 62.663 25.394 ;
      RECT MASK 1 65.383 22.0915 65.463 25.394 ;
      RECT MASK 1 65.715 22.0915 65.795 25.394 ;
      RECT MASK 1 66.545 22.0915 66.625 25.394 ;
      RECT MASK 1 66.877 22.0915 66.957 25.394 ;
      RECT MASK 1 67.707 22.0915 67.787 25.394 ;
      RECT MASK 1 68.039 22.0915 68.119 25.394 ;
      RECT MASK 1 68.869 22.0915 68.949 25.394 ;
      RECT MASK 1 69.201 22.0915 69.281 25.394 ;
      RECT MASK 1 72.001 22.0915 72.081 25.394 ;
      RECT MASK 1 72.333 22.0915 72.413 25.394 ;
      RECT MASK 1 73.163 22.0915 73.243 25.394 ;
      RECT MASK 1 73.495 22.0915 73.575 25.394 ;
      RECT MASK 1 74.325 22.0915 74.405 25.394 ;
      RECT MASK 1 74.657 22.0915 74.737 25.394 ;
      RECT MASK 1 75.487 22.0915 75.567 25.394 ;
      RECT MASK 1 75.819 22.0915 75.899 25.394 ;
      RECT MASK 1 78.619 22.0915 78.699 25.394 ;
      RECT MASK 1 78.951 22.0915 79.031 25.394 ;
      RECT MASK 1 79.781 22.0915 79.861 25.394 ;
      RECT MASK 1 80.113 22.0915 80.193 25.394 ;
      RECT MASK 1 80.943 22.0915 81.023 25.394 ;
      RECT MASK 1 81.275 22.0915 81.355 25.394 ;
      RECT MASK 1 82.105 22.0915 82.185 25.394 ;
      RECT MASK 1 82.437 22.0915 82.517 25.394 ;
      RECT MASK 1 85.237 22.0915 85.317 25.394 ;
      RECT MASK 1 85.569 22.0915 85.649 25.394 ;
      RECT MASK 1 86.399 22.0915 86.479 25.394 ;
      RECT MASK 1 86.731 22.0915 86.811 25.394 ;
      RECT MASK 1 87.561 22.0915 87.641 25.394 ;
      RECT MASK 1 87.893 22.0915 87.973 25.394 ;
      RECT MASK 1 88.723 22.0915 88.803 25.394 ;
      RECT MASK 1 89.055 22.0915 89.135 25.394 ;
      RECT MASK 1 91.855 22.0915 91.935 25.394 ;
      RECT MASK 1 92.187 22.0915 92.267 25.394 ;
      RECT MASK 1 93.017 22.0915 93.097 25.394 ;
      RECT MASK 1 93.349 22.0915 93.429 25.394 ;
      RECT MASK 1 94.179 22.0915 94.259 25.394 ;
      RECT MASK 1 94.511 22.0915 94.591 25.394 ;
      RECT MASK 1 95.341 22.0915 95.421 25.394 ;
      RECT MASK 1 95.673 22.0915 95.753 25.394 ;
      RECT MASK 1 98.473 22.0915 98.553 25.394 ;
      RECT MASK 1 98.805 22.0915 98.885 25.394 ;
      RECT MASK 1 99.635 22.0915 99.715 25.394 ;
      RECT MASK 1 99.967 22.0915 100.047 25.394 ;
      RECT MASK 1 100.797 22.0915 100.877 25.394 ;
      RECT MASK 1 101.129 22.0915 101.209 25.394 ;
      RECT MASK 1 101.959 22.0915 102.039 25.394 ;
      RECT MASK 1 102.291 22.0915 102.371 25.394 ;
      RECT MASK 1 105.091 22.0915 105.171 25.394 ;
      RECT MASK 1 105.423 22.0915 105.503 25.394 ;
      RECT MASK 1 106.253 22.0915 106.333 25.394 ;
      RECT MASK 1 106.585 22.0915 106.665 25.394 ;
      RECT MASK 1 107.415 22.0915 107.495 25.394 ;
      RECT MASK 1 107.747 22.0915 107.827 25.394 ;
      RECT MASK 1 108.577 22.0915 108.657 25.394 ;
      RECT MASK 1 108.909 22.0915 108.989 25.394 ;
      RECT MASK 1 10.23 22.466 10.29 22.686 ;
      RECT MASK 1 12.034 22.466 12.094 22.686 ;
      RECT MASK 1 16.848 22.466 16.908 22.686 ;
      RECT MASK 1 18.652 22.466 18.712 22.686 ;
      RECT MASK 1 23.466 22.466 23.526 22.686 ;
      RECT MASK 1 25.27 22.466 25.33 22.686 ;
      RECT MASK 1 30.084 22.466 30.144 22.686 ;
      RECT MASK 1 31.888 22.466 31.948 22.686 ;
      RECT MASK 1 36.702 22.466 36.762 22.686 ;
      RECT MASK 1 38.506 22.466 38.566 22.686 ;
      RECT MASK 1 43.32 22.466 43.38 22.686 ;
      RECT MASK 1 45.124 22.466 45.184 22.686 ;
      RECT MASK 1 49.938 22.466 49.998 22.686 ;
      RECT MASK 1 51.742 22.466 51.802 22.686 ;
      RECT MASK 1 56.556 22.466 56.616 22.686 ;
      RECT MASK 1 58.36 22.466 58.42 22.686 ;
      RECT MASK 1 63.174 22.466 63.234 22.686 ;
      RECT MASK 1 64.978 22.466 65.038 22.686 ;
      RECT MASK 1 69.792 22.466 69.852 22.686 ;
      RECT MASK 1 71.596 22.466 71.656 22.686 ;
      RECT MASK 1 76.41 22.466 76.47 22.686 ;
      RECT MASK 1 78.214 22.466 78.274 22.686 ;
      RECT MASK 1 83.028 22.466 83.088 22.686 ;
      RECT MASK 1 84.832 22.466 84.892 22.686 ;
      RECT MASK 1 89.646 22.466 89.706 22.686 ;
      RECT MASK 1 91.45 22.466 91.51 22.686 ;
      RECT MASK 1 96.264 22.466 96.324 22.686 ;
      RECT MASK 1 98.068 22.466 98.128 22.686 ;
      RECT MASK 1 102.882 22.466 102.942 22.686 ;
      RECT MASK 1 104.686 22.466 104.746 22.686 ;
      RECT MASK 1 109.5 22.466 109.56 22.686 ;
      RECT MASK 1 5.167 23.731 5.227 25.966 ;
      RECT MASK 1 10.479 23.731 10.539 25.966 ;
      RECT MASK 1 11.785 23.731 11.845 25.966 ;
      RECT MASK 1 17.097 23.731 17.157 25.966 ;
      RECT MASK 1 18.403 23.731 18.463 25.966 ;
      RECT MASK 1 23.715 23.735 23.775 25.945 ;
      RECT MASK 1 25.021 23.735 25.081 25.945 ;
      RECT MASK 1 30.333 23.735 30.393 25.945 ;
      RECT MASK 1 31.639 23.735 31.699 25.945 ;
      RECT MASK 1 36.951 23.735 37.011 25.945 ;
      RECT MASK 1 38.257 23.735 38.317 25.945 ;
      RECT MASK 1 43.569 23.735 43.629 25.945 ;
      RECT MASK 1 44.875 23.735 44.935 25.945 ;
      RECT MASK 1 50.187 23.735 50.247 25.945 ;
      RECT MASK 1 51.493 23.735 51.553 25.945 ;
      RECT MASK 1 56.805 23.735 56.865 25.945 ;
      RECT MASK 1 58.111 23.735 58.171 25.945 ;
      RECT MASK 1 63.423 23.735 63.483 25.945 ;
      RECT MASK 1 64.729 23.735 64.789 25.945 ;
      RECT MASK 1 70.041 23.735 70.101 25.945 ;
      RECT MASK 1 71.347 23.735 71.407 25.945 ;
      RECT MASK 1 76.659 23.735 76.719 25.945 ;
      RECT MASK 1 77.965 23.735 78.025 25.945 ;
      RECT MASK 1 83.277 23.735 83.337 25.945 ;
      RECT MASK 1 84.583 23.735 84.643 25.945 ;
      RECT MASK 1 89.895 23.735 89.955 25.945 ;
      RECT MASK 1 91.201 23.735 91.261 25.945 ;
      RECT MASK 1 96.513 23.735 96.573 25.945 ;
      RECT MASK 1 97.819 23.735 97.879 25.945 ;
      RECT MASK 1 103.131 23.735 103.191 25.945 ;
      RECT MASK 1 104.437 23.735 104.497 25.945 ;
      RECT MASK 1 109.749 23.735 109.809 25.945 ;
      RECT MASK 1 10.23 24.19 10.29 24.41 ;
      RECT MASK 1 12.034 24.19 12.094 24.41 ;
      RECT MASK 1 16.848 24.19 16.908 24.41 ;
      RECT MASK 1 18.652 24.19 18.712 24.41 ;
      RECT MASK 1 23.466 24.19 23.526 24.41 ;
      RECT MASK 1 25.27 24.19 25.33 24.41 ;
      RECT MASK 1 30.084 24.19 30.144 24.41 ;
      RECT MASK 1 31.888 24.19 31.948 24.41 ;
      RECT MASK 1 36.702 24.19 36.762 24.41 ;
      RECT MASK 1 38.506 24.19 38.566 24.41 ;
      RECT MASK 1 43.32 24.19 43.38 24.41 ;
      RECT MASK 1 45.124 24.19 45.184 24.41 ;
      RECT MASK 1 49.938 24.19 49.998 24.41 ;
      RECT MASK 1 51.742 24.19 51.802 24.41 ;
      RECT MASK 1 56.556 24.19 56.616 24.41 ;
      RECT MASK 1 58.36 24.19 58.42 24.41 ;
      RECT MASK 1 63.174 24.19 63.234 24.41 ;
      RECT MASK 1 64.978 24.19 65.038 24.41 ;
      RECT MASK 1 69.792 24.19 69.852 24.41 ;
      RECT MASK 1 71.596 24.19 71.656 24.41 ;
      RECT MASK 1 76.41 24.19 76.47 24.41 ;
      RECT MASK 1 78.214 24.19 78.274 24.41 ;
      RECT MASK 1 83.028 24.19 83.088 24.41 ;
      RECT MASK 1 84.832 24.19 84.892 24.41 ;
      RECT MASK 1 89.646 24.19 89.706 24.41 ;
      RECT MASK 1 91.45 24.19 91.51 24.41 ;
      RECT MASK 1 96.264 24.19 96.324 24.41 ;
      RECT MASK 1 98.068 24.19 98.128 24.41 ;
      RECT MASK 1 102.882 24.19 102.942 24.41 ;
      RECT MASK 1 104.686 24.19 104.746 24.41 ;
      RECT MASK 1 109.5 24.19 109.56 24.41 ;
      RECT MASK 1 5.831 25.68 5.891 25.95 ;
      RECT MASK 1 6.163 25.68 6.223 25.95 ;
      RECT MASK 1 6.495 25.68 6.555 25.95 ;
      RECT MASK 1 6.993 25.68 7.053 25.95 ;
      RECT MASK 1 7.325 25.68 7.385 25.95 ;
      RECT MASK 1 7.657 25.68 7.717 25.95 ;
      RECT MASK 1 8.155 25.68 8.215 25.95 ;
      RECT MASK 1 8.487 25.68 8.547 25.95 ;
      RECT MASK 1 8.819 25.68 8.879 25.95 ;
      RECT MASK 1 9.317 25.68 9.377 25.95 ;
      RECT MASK 1 9.649 25.68 9.709 25.95 ;
      RECT MASK 1 9.981 25.68 10.041 25.95 ;
      RECT MASK 1 12.449 25.68 12.509 25.95 ;
      RECT MASK 1 12.781 25.68 12.841 25.95 ;
      RECT MASK 1 13.113 25.68 13.173 25.95 ;
      RECT MASK 1 13.611 25.68 13.671 25.95 ;
      RECT MASK 1 13.943 25.68 14.003 25.95 ;
      RECT MASK 1 14.275 25.68 14.335 25.95 ;
      RECT MASK 1 14.773 25.68 14.833 25.95 ;
      RECT MASK 1 15.105 25.68 15.165 25.95 ;
      RECT MASK 1 15.437 25.68 15.497 25.95 ;
      RECT MASK 1 15.935 25.68 15.995 25.95 ;
      RECT MASK 1 16.267 25.68 16.327 25.95 ;
      RECT MASK 1 16.599 25.68 16.659 25.95 ;
      RECT MASK 1 19.067 25.68 19.127 25.95 ;
      RECT MASK 1 19.399 25.68 19.459 25.95 ;
      RECT MASK 1 19.731 25.68 19.791 25.95 ;
      RECT MASK 1 20.229 25.68 20.289 25.95 ;
      RECT MASK 1 20.561 25.68 20.621 25.95 ;
      RECT MASK 1 20.893 25.68 20.953 25.95 ;
      RECT MASK 1 21.391 25.68 21.451 25.95 ;
      RECT MASK 1 21.723 25.68 21.783 25.95 ;
      RECT MASK 1 22.055 25.68 22.115 25.95 ;
      RECT MASK 1 22.553 25.68 22.613 25.95 ;
      RECT MASK 1 22.885 25.68 22.945 25.95 ;
      RECT MASK 1 23.217 25.68 23.277 25.95 ;
      RECT MASK 1 25.685 25.68 25.745 25.95 ;
      RECT MASK 1 26.017 25.68 26.077 25.95 ;
      RECT MASK 1 26.349 25.68 26.409 25.95 ;
      RECT MASK 1 26.847 25.68 26.907 25.95 ;
      RECT MASK 1 27.179 25.68 27.239 25.95 ;
      RECT MASK 1 27.511 25.68 27.571 25.95 ;
      RECT MASK 1 28.009 25.68 28.069 25.95 ;
      RECT MASK 1 28.341 25.68 28.401 25.95 ;
      RECT MASK 1 28.673 25.68 28.733 25.95 ;
      RECT MASK 1 29.171 25.68 29.231 25.95 ;
      RECT MASK 1 29.503 25.68 29.563 25.95 ;
      RECT MASK 1 29.835 25.68 29.895 25.95 ;
      RECT MASK 1 32.303 25.68 32.363 25.95 ;
      RECT MASK 1 32.635 25.68 32.695 25.95 ;
      RECT MASK 1 32.967 25.68 33.027 25.95 ;
      RECT MASK 1 33.465 25.68 33.525 25.95 ;
      RECT MASK 1 33.797 25.68 33.857 25.95 ;
      RECT MASK 1 34.129 25.68 34.189 25.95 ;
      RECT MASK 1 34.627 25.68 34.687 25.95 ;
      RECT MASK 1 34.959 25.68 35.019 25.95 ;
      RECT MASK 1 35.291 25.68 35.351 25.95 ;
      RECT MASK 1 35.789 25.68 35.849 25.95 ;
      RECT MASK 1 36.121 25.68 36.181 25.95 ;
      RECT MASK 1 36.453 25.68 36.513 25.95 ;
      RECT MASK 1 38.921 25.68 38.981 25.95 ;
      RECT MASK 1 39.253 25.68 39.313 25.95 ;
      RECT MASK 1 39.585 25.68 39.645 25.95 ;
      RECT MASK 1 40.083 25.68 40.143 25.95 ;
      RECT MASK 1 40.415 25.68 40.475 25.95 ;
      RECT MASK 1 40.747 25.68 40.807 25.95 ;
      RECT MASK 1 41.245 25.68 41.305 25.95 ;
      RECT MASK 1 41.577 25.68 41.637 25.95 ;
      RECT MASK 1 41.909 25.68 41.969 25.95 ;
      RECT MASK 1 42.407 25.68 42.467 25.95 ;
      RECT MASK 1 42.739 25.68 42.799 25.95 ;
      RECT MASK 1 43.071 25.68 43.131 25.95 ;
      RECT MASK 1 45.539 25.68 45.599 25.95 ;
      RECT MASK 1 45.871 25.68 45.931 25.95 ;
      RECT MASK 1 46.203 25.68 46.263 25.95 ;
      RECT MASK 1 46.701 25.68 46.761 25.95 ;
      RECT MASK 1 47.033 25.68 47.093 25.95 ;
      RECT MASK 1 47.365 25.68 47.425 25.95 ;
      RECT MASK 1 47.863 25.68 47.923 25.95 ;
      RECT MASK 1 48.195 25.68 48.255 25.95 ;
      RECT MASK 1 48.527 25.68 48.587 25.95 ;
      RECT MASK 1 49.025 25.68 49.085 25.95 ;
      RECT MASK 1 49.357 25.68 49.417 25.95 ;
      RECT MASK 1 49.689 25.68 49.749 25.95 ;
      RECT MASK 1 52.157 25.68 52.217 25.95 ;
      RECT MASK 1 52.489 25.68 52.549 25.95 ;
      RECT MASK 1 52.821 25.68 52.881 25.95 ;
      RECT MASK 1 53.319 25.68 53.379 25.95 ;
      RECT MASK 1 53.651 25.68 53.711 25.95 ;
      RECT MASK 1 53.983 25.68 54.043 25.95 ;
      RECT MASK 1 54.481 25.68 54.541 25.95 ;
      RECT MASK 1 54.813 25.68 54.873 25.95 ;
      RECT MASK 1 55.145 25.68 55.205 25.95 ;
      RECT MASK 1 55.643 25.68 55.703 25.95 ;
      RECT MASK 1 55.975 25.68 56.035 25.95 ;
      RECT MASK 1 56.307 25.68 56.367 25.95 ;
      RECT MASK 1 58.775 25.68 58.835 25.95 ;
      RECT MASK 1 59.107 25.68 59.167 25.95 ;
      RECT MASK 1 59.439 25.68 59.499 25.95 ;
      RECT MASK 1 59.937 25.68 59.997 25.95 ;
      RECT MASK 1 60.269 25.68 60.329 25.95 ;
      RECT MASK 1 60.601 25.68 60.661 25.95 ;
      RECT MASK 1 61.099 25.68 61.159 25.95 ;
      RECT MASK 1 61.431 25.68 61.491 25.95 ;
      RECT MASK 1 61.763 25.68 61.823 25.95 ;
      RECT MASK 1 62.261 25.68 62.321 25.95 ;
      RECT MASK 1 62.593 25.68 62.653 25.95 ;
      RECT MASK 1 62.925 25.68 62.985 25.95 ;
      RECT MASK 1 65.393 25.68 65.453 25.95 ;
      RECT MASK 1 65.725 25.68 65.785 25.95 ;
      RECT MASK 1 66.057 25.68 66.117 25.95 ;
      RECT MASK 1 66.555 25.68 66.615 25.95 ;
      RECT MASK 1 66.887 25.68 66.947 25.95 ;
      RECT MASK 1 67.219 25.68 67.279 25.95 ;
      RECT MASK 1 67.717 25.68 67.777 25.95 ;
      RECT MASK 1 68.049 25.68 68.109 25.95 ;
      RECT MASK 1 68.381 25.68 68.441 25.95 ;
      RECT MASK 1 68.879 25.68 68.939 25.95 ;
      RECT MASK 1 69.211 25.68 69.271 25.95 ;
      RECT MASK 1 69.543 25.68 69.603 25.95 ;
      RECT MASK 1 72.011 25.68 72.071 25.95 ;
      RECT MASK 1 72.343 25.68 72.403 25.95 ;
      RECT MASK 1 72.675 25.68 72.735 25.95 ;
      RECT MASK 1 73.173 25.68 73.233 25.95 ;
      RECT MASK 1 73.505 25.68 73.565 25.95 ;
      RECT MASK 1 73.837 25.68 73.897 25.95 ;
      RECT MASK 1 74.335 25.68 74.395 25.95 ;
      RECT MASK 1 74.667 25.68 74.727 25.95 ;
      RECT MASK 1 74.999 25.68 75.059 25.95 ;
      RECT MASK 1 75.497 25.68 75.557 25.95 ;
      RECT MASK 1 75.829 25.68 75.889 25.95 ;
      RECT MASK 1 76.161 25.68 76.221 25.95 ;
      RECT MASK 1 78.629 25.68 78.689 25.95 ;
      RECT MASK 1 78.961 25.68 79.021 25.95 ;
      RECT MASK 1 79.293 25.68 79.353 25.95 ;
      RECT MASK 1 79.791 25.68 79.851 25.95 ;
      RECT MASK 1 80.123 25.68 80.183 25.95 ;
      RECT MASK 1 80.455 25.68 80.515 25.95 ;
      RECT MASK 1 80.953 25.68 81.013 25.95 ;
      RECT MASK 1 81.285 25.68 81.345 25.95 ;
      RECT MASK 1 81.617 25.68 81.677 25.95 ;
      RECT MASK 1 82.115 25.68 82.175 25.95 ;
      RECT MASK 1 82.447 25.68 82.507 25.95 ;
      RECT MASK 1 82.779 25.68 82.839 25.95 ;
      RECT MASK 1 85.247 25.68 85.307 25.95 ;
      RECT MASK 1 85.579 25.68 85.639 25.95 ;
      RECT MASK 1 85.911 25.68 85.971 25.95 ;
      RECT MASK 1 86.409 25.68 86.469 25.95 ;
      RECT MASK 1 86.741 25.68 86.801 25.95 ;
      RECT MASK 1 87.073 25.68 87.133 25.95 ;
      RECT MASK 1 87.571 25.68 87.631 25.95 ;
      RECT MASK 1 87.903 25.68 87.963 25.95 ;
      RECT MASK 1 88.235 25.68 88.295 25.95 ;
      RECT MASK 1 88.733 25.68 88.793 25.95 ;
      RECT MASK 1 89.065 25.68 89.125 25.95 ;
      RECT MASK 1 89.397 25.68 89.457 25.95 ;
      RECT MASK 1 91.865 25.68 91.925 25.95 ;
      RECT MASK 1 92.197 25.68 92.257 25.95 ;
      RECT MASK 1 92.529 25.68 92.589 25.95 ;
      RECT MASK 1 93.027 25.68 93.087 25.95 ;
      RECT MASK 1 93.359 25.68 93.419 25.95 ;
      RECT MASK 1 93.691 25.68 93.751 25.95 ;
      RECT MASK 1 94.189 25.68 94.249 25.95 ;
      RECT MASK 1 94.521 25.68 94.581 25.95 ;
      RECT MASK 1 94.853 25.68 94.913 25.95 ;
      RECT MASK 1 95.351 25.68 95.411 25.95 ;
      RECT MASK 1 95.683 25.68 95.743 25.95 ;
      RECT MASK 1 96.015 25.68 96.075 25.95 ;
      RECT MASK 1 98.483 25.68 98.543 25.95 ;
      RECT MASK 1 98.815 25.68 98.875 25.95 ;
      RECT MASK 1 99.147 25.68 99.207 25.95 ;
      RECT MASK 1 99.645 25.68 99.705 25.95 ;
      RECT MASK 1 99.977 25.68 100.037 25.95 ;
      RECT MASK 1 100.309 25.68 100.369 25.95 ;
      RECT MASK 1 100.807 25.68 100.867 25.95 ;
      RECT MASK 1 101.139 25.68 101.199 25.95 ;
      RECT MASK 1 101.471 25.68 101.531 25.95 ;
      RECT MASK 1 101.969 25.68 102.029 25.95 ;
      RECT MASK 1 102.301 25.68 102.361 25.95 ;
      RECT MASK 1 102.633 25.68 102.693 25.95 ;
      RECT MASK 1 105.101 25.68 105.161 25.95 ;
      RECT MASK 1 105.433 25.68 105.493 25.95 ;
      RECT MASK 1 105.765 25.68 105.825 25.95 ;
      RECT MASK 1 106.263 25.68 106.323 25.95 ;
      RECT MASK 1 106.595 25.68 106.655 25.95 ;
      RECT MASK 1 106.927 25.68 106.987 25.95 ;
      RECT MASK 1 107.425 25.68 107.485 25.95 ;
      RECT MASK 1 107.757 25.68 107.817 25.95 ;
      RECT MASK 1 108.089 25.68 108.149 25.95 ;
      RECT MASK 1 108.587 25.68 108.647 25.95 ;
      RECT MASK 1 108.919 25.68 108.979 25.95 ;
      RECT MASK 1 109.251 25.68 109.311 25.95 ;
      RECT MASK 1 3.589 26.1 3.889 77.8205 ;
      RECT MASK 1 2.005 26.156 2.085 26.476 ;
      RECT MASK 1 2.337 26.156 2.417 26.476 ;
      RECT MASK 1 2.669 26.156 2.749 26.476 ;
      RECT MASK 1 4.329 26.156 4.409 26.476 ;
      RECT MASK 1 4.661 26.156 4.741 26.476 ;
      RECT MASK 1 4.993 26.156 5.073 26.476 ;
      RECT MASK 1 5.325 26.156 5.405 26.476 ;
      RECT MASK 1 5.657 26.156 5.737 26.476 ;
      RECT MASK 1 5.989 26.156 6.069 26.476 ;
      RECT MASK 1 6.321 26.156 6.401 26.476 ;
      RECT MASK 1 6.653 26.156 6.733 26.476 ;
      RECT MASK 1 6.985 26.156 7.065 26.476 ;
      RECT MASK 1 7.317 26.156 7.397 26.476 ;
      RECT MASK 1 7.649 26.156 7.729 26.476 ;
      RECT MASK 1 7.981 26.156 8.061 26.476 ;
      RECT MASK 1 8.313 26.156 8.393 26.476 ;
      RECT MASK 1 8.645 26.156 8.725 26.476 ;
      RECT MASK 1 8.977 26.156 9.057 26.476 ;
      RECT MASK 1 9.309 26.156 9.389 26.476 ;
      RECT MASK 1 9.641 26.156 9.721 26.476 ;
      RECT MASK 1 9.973 26.156 10.053 26.476 ;
      RECT MASK 1 10.305 26.156 10.385 26.476 ;
      RECT MASK 1 10.637 26.156 10.717 26.476 ;
      RECT MASK 1 10.969 26.156 11.049 26.476 ;
      RECT MASK 1 11.301 26.156 11.381 26.476 ;
      RECT MASK 1 11.633 26.156 11.713 26.476 ;
      RECT MASK 1 11.965 26.156 12.045 26.476 ;
      RECT MASK 1 12.297 26.156 12.377 26.476 ;
      RECT MASK 1 12.629 26.156 12.709 26.476 ;
      RECT MASK 1 12.961 26.156 13.041 26.476 ;
      RECT MASK 1 13.293 26.156 13.373 26.476 ;
      RECT MASK 1 13.625 26.156 13.705 26.476 ;
      RECT MASK 1 13.957 26.156 14.037 26.476 ;
      RECT MASK 1 14.289 26.156 14.369 26.476 ;
      RECT MASK 1 14.621 26.156 14.701 26.476 ;
      RECT MASK 1 14.953 26.156 15.033 26.476 ;
      RECT MASK 1 15.285 26.156 15.365 26.476 ;
      RECT MASK 1 15.617 26.156 15.697 26.476 ;
      RECT MASK 1 15.949 26.156 16.029 26.476 ;
      RECT MASK 1 16.281 26.156 16.361 26.476 ;
      RECT MASK 1 16.613 26.156 16.693 26.476 ;
      RECT MASK 1 16.945 26.156 17.025 26.476 ;
      RECT MASK 1 17.277 26.156 17.357 26.476 ;
      RECT MASK 1 17.609 26.156 17.689 26.476 ;
      RECT MASK 1 17.941 26.156 18.021 26.476 ;
      RECT MASK 1 18.273 26.156 18.353 26.476 ;
      RECT MASK 1 18.605 26.156 18.685 26.476 ;
      RECT MASK 1 18.937 26.156 19.017 26.476 ;
      RECT MASK 1 19.269 26.156 19.349 26.476 ;
      RECT MASK 1 19.601 26.156 19.681 26.476 ;
      RECT MASK 1 19.933 26.156 20.013 26.476 ;
      RECT MASK 1 20.265 26.156 20.345 26.476 ;
      RECT MASK 1 20.597 26.156 20.677 26.476 ;
      RECT MASK 1 20.929 26.156 21.009 26.476 ;
      RECT MASK 1 21.261 26.156 21.341 26.476 ;
      RECT MASK 1 21.593 26.156 21.673 26.476 ;
      RECT MASK 1 21.925 26.156 22.005 26.476 ;
      RECT MASK 1 22.257 26.156 22.337 26.476 ;
      RECT MASK 1 22.589 26.156 22.669 26.476 ;
      RECT MASK 1 22.921 26.156 23.001 26.476 ;
      RECT MASK 1 23.253 26.156 23.333 26.476 ;
      RECT MASK 1 23.585 26.156 23.665 26.476 ;
      RECT MASK 1 23.917 26.156 23.997 26.476 ;
      RECT MASK 1 24.249 26.156 24.329 26.476 ;
      RECT MASK 1 24.581 26.156 24.661 26.476 ;
      RECT MASK 1 24.913 26.156 24.993 26.476 ;
      RECT MASK 1 25.245 26.156 25.325 26.476 ;
      RECT MASK 1 25.577 26.156 25.657 26.476 ;
      RECT MASK 1 25.909 26.156 25.989 26.476 ;
      RECT MASK 1 26.241 26.156 26.321 26.476 ;
      RECT MASK 1 26.573 26.156 26.653 26.476 ;
      RECT MASK 1 26.905 26.156 26.985 26.476 ;
      RECT MASK 1 27.237 26.156 27.317 26.476 ;
      RECT MASK 1 27.569 26.156 27.649 26.476 ;
      RECT MASK 1 27.901 26.156 27.981 26.476 ;
      RECT MASK 1 28.233 26.156 28.313 26.476 ;
      RECT MASK 1 28.565 26.156 28.645 26.476 ;
      RECT MASK 1 28.897 26.156 28.977 26.476 ;
      RECT MASK 1 29.229 26.156 29.309 26.476 ;
      RECT MASK 1 29.561 26.156 29.641 26.476 ;
      RECT MASK 1 29.893 26.156 29.973 26.476 ;
      RECT MASK 1 30.225 26.156 30.305 26.476 ;
      RECT MASK 1 30.557 26.156 30.637 26.476 ;
      RECT MASK 1 30.889 26.156 30.969 26.476 ;
      RECT MASK 1 31.221 26.156 31.301 26.476 ;
      RECT MASK 1 31.553 26.156 31.633 26.476 ;
      RECT MASK 1 31.885 26.156 31.965 26.476 ;
      RECT MASK 1 32.217 26.156 32.297 26.476 ;
      RECT MASK 1 32.549 26.156 32.629 26.476 ;
      RECT MASK 1 32.881 26.156 32.961 26.476 ;
      RECT MASK 1 33.213 26.156 33.293 26.476 ;
      RECT MASK 1 33.545 26.156 33.625 26.476 ;
      RECT MASK 1 33.877 26.156 33.957 26.476 ;
      RECT MASK 1 34.209 26.156 34.289 26.476 ;
      RECT MASK 1 34.541 26.156 34.621 26.476 ;
      RECT MASK 1 34.873 26.156 34.953 26.476 ;
      RECT MASK 1 35.205 26.156 35.285 26.476 ;
      RECT MASK 1 35.537 26.156 35.617 26.476 ;
      RECT MASK 1 35.869 26.156 35.949 26.476 ;
      RECT MASK 1 36.201 26.156 36.281 26.476 ;
      RECT MASK 1 36.533 26.156 36.613 26.476 ;
      RECT MASK 1 36.865 26.156 36.945 26.476 ;
      RECT MASK 1 37.197 26.156 37.277 26.476 ;
      RECT MASK 1 37.529 26.156 37.609 26.476 ;
      RECT MASK 1 37.861 26.156 37.941 26.476 ;
      RECT MASK 1 38.193 26.156 38.273 26.476 ;
      RECT MASK 1 38.525 26.156 38.605 26.476 ;
      RECT MASK 1 38.857 26.156 38.937 26.476 ;
      RECT MASK 1 39.189 26.156 39.269 26.476 ;
      RECT MASK 1 39.521 26.156 39.601 26.476 ;
      RECT MASK 1 39.853 26.156 39.933 26.476 ;
      RECT MASK 1 40.185 26.156 40.265 26.476 ;
      RECT MASK 1 40.517 26.156 40.597 26.476 ;
      RECT MASK 1 40.849 26.156 40.929 26.476 ;
      RECT MASK 1 41.181 26.156 41.261 26.476 ;
      RECT MASK 1 41.513 26.156 41.593 26.476 ;
      RECT MASK 1 41.845 26.156 41.925 26.476 ;
      RECT MASK 1 42.177 26.156 42.257 26.476 ;
      RECT MASK 1 42.509 26.156 42.589 26.476 ;
      RECT MASK 1 42.841 26.156 42.921 26.476 ;
      RECT MASK 1 43.173 26.156 43.253 26.476 ;
      RECT MASK 1 43.505 26.156 43.585 26.476 ;
      RECT MASK 1 43.837 26.156 43.917 26.476 ;
      RECT MASK 1 44.169 26.156 44.249 26.476 ;
      RECT MASK 1 44.501 26.156 44.581 26.476 ;
      RECT MASK 1 44.833 26.156 44.913 26.476 ;
      RECT MASK 1 45.165 26.156 45.245 26.476 ;
      RECT MASK 1 45.497 26.156 45.577 26.476 ;
      RECT MASK 1 45.829 26.156 45.909 26.476 ;
      RECT MASK 1 46.161 26.156 46.241 26.476 ;
      RECT MASK 1 46.493 26.156 46.573 26.476 ;
      RECT MASK 1 46.825 26.156 46.905 26.476 ;
      RECT MASK 1 47.157 26.156 47.237 26.476 ;
      RECT MASK 1 47.489 26.156 47.569 26.476 ;
      RECT MASK 1 47.821 26.156 47.901 26.476 ;
      RECT MASK 1 48.153 26.156 48.233 26.476 ;
      RECT MASK 1 48.485 26.156 48.565 26.476 ;
      RECT MASK 1 48.817 26.156 48.897 26.476 ;
      RECT MASK 1 49.149 26.156 49.229 26.476 ;
      RECT MASK 1 49.481 26.156 49.561 26.476 ;
      RECT MASK 1 49.813 26.156 49.893 26.476 ;
      RECT MASK 1 50.145 26.156 50.225 26.476 ;
      RECT MASK 1 50.477 26.156 50.557 26.476 ;
      RECT MASK 1 50.809 26.156 50.889 26.476 ;
      RECT MASK 1 51.141 26.156 51.221 26.476 ;
      RECT MASK 1 51.473 26.156 51.553 26.476 ;
      RECT MASK 1 51.805 26.156 51.885 26.476 ;
      RECT MASK 1 52.137 26.156 52.217 26.476 ;
      RECT MASK 1 52.469 26.156 52.549 26.476 ;
      RECT MASK 1 52.801 26.156 52.881 26.476 ;
      RECT MASK 1 53.133 26.156 53.213 26.476 ;
      RECT MASK 1 53.465 26.156 53.545 26.476 ;
      RECT MASK 1 53.797 26.156 53.877 26.476 ;
      RECT MASK 1 54.129 26.156 54.209 26.476 ;
      RECT MASK 1 54.461 26.156 54.541 26.476 ;
      RECT MASK 1 54.793 26.156 54.873 26.476 ;
      RECT MASK 1 55.125 26.156 55.205 26.476 ;
      RECT MASK 1 55.457 26.156 55.537 26.476 ;
      RECT MASK 1 55.789 26.156 55.869 26.476 ;
      RECT MASK 1 56.121 26.156 56.201 26.476 ;
      RECT MASK 1 56.453 26.156 56.533 26.476 ;
      RECT MASK 1 56.785 26.156 56.865 26.476 ;
      RECT MASK 1 57.117 26.156 57.197 26.476 ;
      RECT MASK 1 57.449 26.156 57.529 26.476 ;
      RECT MASK 1 57.781 26.156 57.861 26.476 ;
      RECT MASK 1 58.113 26.156 58.193 26.476 ;
      RECT MASK 1 58.445 26.156 58.525 26.476 ;
      RECT MASK 1 58.777 26.156 58.857 26.476 ;
      RECT MASK 1 59.109 26.156 59.189 26.476 ;
      RECT MASK 1 59.441 26.156 59.521 26.476 ;
      RECT MASK 1 59.773 26.156 59.853 26.476 ;
      RECT MASK 1 60.105 26.156 60.185 26.476 ;
      RECT MASK 1 60.437 26.156 60.517 26.476 ;
      RECT MASK 1 60.769 26.156 60.849 26.476 ;
      RECT MASK 1 61.101 26.156 61.181 26.476 ;
      RECT MASK 1 61.433 26.156 61.513 26.476 ;
      RECT MASK 1 61.765 26.156 61.845 26.476 ;
      RECT MASK 1 62.097 26.156 62.177 26.476 ;
      RECT MASK 1 62.429 26.156 62.509 26.476 ;
      RECT MASK 1 62.761 26.156 62.841 26.476 ;
      RECT MASK 1 63.093 26.156 63.173 26.476 ;
      RECT MASK 1 63.425 26.156 63.505 26.476 ;
      RECT MASK 1 63.757 26.156 63.837 26.476 ;
      RECT MASK 1 64.089 26.156 64.169 26.476 ;
      RECT MASK 1 64.421 26.156 64.501 26.476 ;
      RECT MASK 1 64.753 26.156 64.833 26.476 ;
      RECT MASK 1 65.085 26.156 65.165 26.476 ;
      RECT MASK 1 65.417 26.156 65.497 26.476 ;
      RECT MASK 1 65.749 26.156 65.829 26.476 ;
      RECT MASK 1 66.081 26.156 66.161 26.476 ;
      RECT MASK 1 66.413 26.156 66.493 26.476 ;
      RECT MASK 1 66.745 26.156 66.825 26.476 ;
      RECT MASK 1 67.077 26.156 67.157 26.476 ;
      RECT MASK 1 67.409 26.156 67.489 26.476 ;
      RECT MASK 1 67.741 26.156 67.821 26.476 ;
      RECT MASK 1 68.073 26.156 68.153 26.476 ;
      RECT MASK 1 68.405 26.156 68.485 26.476 ;
      RECT MASK 1 68.737 26.156 68.817 26.476 ;
      RECT MASK 1 69.069 26.156 69.149 26.476 ;
      RECT MASK 1 69.401 26.156 69.481 26.476 ;
      RECT MASK 1 69.733 26.156 69.813 26.476 ;
      RECT MASK 1 70.065 26.156 70.145 26.476 ;
      RECT MASK 1 70.397 26.156 70.477 26.476 ;
      RECT MASK 1 70.729 26.156 70.809 26.476 ;
      RECT MASK 1 71.061 26.156 71.141 26.476 ;
      RECT MASK 1 71.393 26.156 71.473 26.476 ;
      RECT MASK 1 71.725 26.156 71.805 26.476 ;
      RECT MASK 1 72.057 26.156 72.137 26.476 ;
      RECT MASK 1 72.389 26.156 72.469 26.476 ;
      RECT MASK 1 72.721 26.156 72.801 26.476 ;
      RECT MASK 1 73.053 26.156 73.133 26.476 ;
      RECT MASK 1 73.385 26.156 73.465 26.476 ;
      RECT MASK 1 73.717 26.156 73.797 26.476 ;
      RECT MASK 1 74.049 26.156 74.129 26.476 ;
      RECT MASK 1 74.381 26.156 74.461 26.476 ;
      RECT MASK 1 74.713 26.156 74.793 26.476 ;
      RECT MASK 1 75.045 26.156 75.125 26.476 ;
      RECT MASK 1 75.377 26.156 75.457 26.476 ;
      RECT MASK 1 75.709 26.156 75.789 26.476 ;
      RECT MASK 1 76.041 26.156 76.121 26.476 ;
      RECT MASK 1 76.373 26.156 76.453 26.476 ;
      RECT MASK 1 76.705 26.156 76.785 26.476 ;
      RECT MASK 1 77.037 26.156 77.117 26.476 ;
      RECT MASK 1 77.369 26.156 77.449 26.476 ;
      RECT MASK 1 77.701 26.156 77.781 26.476 ;
      RECT MASK 1 78.033 26.156 78.113 26.476 ;
      RECT MASK 1 78.365 26.156 78.445 26.476 ;
      RECT MASK 1 78.697 26.156 78.777 26.476 ;
      RECT MASK 1 79.029 26.156 79.109 26.476 ;
      RECT MASK 1 79.361 26.156 79.441 26.476 ;
      RECT MASK 1 79.693 26.156 79.773 26.476 ;
      RECT MASK 1 80.025 26.156 80.105 26.476 ;
      RECT MASK 1 80.357 26.156 80.437 26.476 ;
      RECT MASK 1 80.689 26.156 80.769 26.476 ;
      RECT MASK 1 81.021 26.156 81.101 26.476 ;
      RECT MASK 1 81.353 26.156 81.433 26.476 ;
      RECT MASK 1 81.685 26.156 81.765 26.476 ;
      RECT MASK 1 82.017 26.156 82.097 26.476 ;
      RECT MASK 1 82.349 26.156 82.429 26.476 ;
      RECT MASK 1 82.681 26.156 82.761 26.476 ;
      RECT MASK 1 83.013 26.156 83.093 26.476 ;
      RECT MASK 1 83.345 26.156 83.425 26.476 ;
      RECT MASK 1 83.677 26.156 83.757 26.476 ;
      RECT MASK 1 84.009 26.156 84.089 26.476 ;
      RECT MASK 1 84.341 26.156 84.421 26.476 ;
      RECT MASK 1 84.673 26.156 84.753 26.476 ;
      RECT MASK 1 85.005 26.156 85.085 26.476 ;
      RECT MASK 1 85.337 26.156 85.417 26.476 ;
      RECT MASK 1 85.669 26.156 85.749 26.476 ;
      RECT MASK 1 86.001 26.156 86.081 26.476 ;
      RECT MASK 1 86.333 26.156 86.413 26.476 ;
      RECT MASK 1 86.665 26.156 86.745 26.476 ;
      RECT MASK 1 86.997 26.156 87.077 26.476 ;
      RECT MASK 1 87.329 26.156 87.409 26.476 ;
      RECT MASK 1 87.661 26.156 87.741 26.476 ;
      RECT MASK 1 87.993 26.156 88.073 26.476 ;
      RECT MASK 1 88.325 26.156 88.405 26.476 ;
      RECT MASK 1 88.657 26.156 88.737 26.476 ;
      RECT MASK 1 88.989 26.156 89.069 26.476 ;
      RECT MASK 1 89.321 26.156 89.401 26.476 ;
      RECT MASK 1 89.653 26.156 89.733 26.476 ;
      RECT MASK 1 89.985 26.156 90.065 26.476 ;
      RECT MASK 1 90.317 26.156 90.397 26.476 ;
      RECT MASK 1 90.649 26.156 90.729 26.476 ;
      RECT MASK 1 90.981 26.156 91.061 26.476 ;
      RECT MASK 1 91.313 26.156 91.393 26.476 ;
      RECT MASK 1 91.645 26.156 91.725 26.476 ;
      RECT MASK 1 91.977 26.156 92.057 26.476 ;
      RECT MASK 1 92.309 26.156 92.389 26.476 ;
      RECT MASK 1 92.641 26.156 92.721 26.476 ;
      RECT MASK 1 92.973 26.156 93.053 26.476 ;
      RECT MASK 1 93.305 26.156 93.385 26.476 ;
      RECT MASK 1 93.637 26.156 93.717 26.476 ;
      RECT MASK 1 93.969 26.156 94.049 26.476 ;
      RECT MASK 1 94.301 26.156 94.381 26.476 ;
      RECT MASK 1 94.633 26.156 94.713 26.476 ;
      RECT MASK 1 94.965 26.156 95.045 26.476 ;
      RECT MASK 1 95.297 26.156 95.377 26.476 ;
      RECT MASK 1 95.629 26.156 95.709 26.476 ;
      RECT MASK 1 95.961 26.156 96.041 26.476 ;
      RECT MASK 1 96.293 26.156 96.373 26.476 ;
      RECT MASK 1 96.625 26.156 96.705 26.476 ;
      RECT MASK 1 96.957 26.156 97.037 26.476 ;
      RECT MASK 1 97.289 26.156 97.369 26.476 ;
      RECT MASK 1 97.621 26.156 97.701 26.476 ;
      RECT MASK 1 97.953 26.156 98.033 26.476 ;
      RECT MASK 1 98.285 26.156 98.365 26.476 ;
      RECT MASK 1 98.617 26.156 98.697 26.476 ;
      RECT MASK 1 98.949 26.156 99.029 26.476 ;
      RECT MASK 1 99.281 26.156 99.361 26.476 ;
      RECT MASK 1 99.613 26.156 99.693 26.476 ;
      RECT MASK 1 99.945 26.156 100.025 26.476 ;
      RECT MASK 1 100.277 26.156 100.357 26.476 ;
      RECT MASK 1 100.609 26.156 100.689 26.476 ;
      RECT MASK 1 100.941 26.156 101.021 26.476 ;
      RECT MASK 1 101.273 26.156 101.353 26.476 ;
      RECT MASK 1 101.605 26.156 101.685 26.476 ;
      RECT MASK 1 101.937 26.156 102.017 26.476 ;
      RECT MASK 1 102.269 26.156 102.349 26.476 ;
      RECT MASK 1 102.601 26.156 102.681 26.476 ;
      RECT MASK 1 102.933 26.156 103.013 26.476 ;
      RECT MASK 1 103.265 26.156 103.345 26.476 ;
      RECT MASK 1 103.597 26.156 103.677 26.476 ;
      RECT MASK 1 103.929 26.156 104.009 26.476 ;
      RECT MASK 1 104.261 26.156 104.341 26.476 ;
      RECT MASK 1 104.593 26.156 104.673 26.476 ;
      RECT MASK 1 104.925 26.156 105.005 26.476 ;
      RECT MASK 1 105.257 26.156 105.337 26.476 ;
      RECT MASK 1 105.589 26.156 105.669 26.476 ;
      RECT MASK 1 105.921 26.156 106.001 26.476 ;
      RECT MASK 1 106.253 26.156 106.333 26.476 ;
      RECT MASK 1 106.585 26.156 106.665 26.476 ;
      RECT MASK 1 106.917 26.156 106.997 26.476 ;
      RECT MASK 1 107.249 26.156 107.329 26.476 ;
      RECT MASK 1 107.581 26.156 107.661 26.476 ;
      RECT MASK 1 107.913 26.156 107.993 26.476 ;
      RECT MASK 1 108.245 26.156 108.325 26.476 ;
      RECT MASK 1 108.577 26.156 108.657 26.476 ;
      RECT MASK 1 108.909 26.156 108.989 26.476 ;
      RECT MASK 1 109.241 26.156 109.321 26.476 ;
      RECT MASK 1 109.573 26.156 109.653 26.476 ;
      RECT MASK 1 109.905 26.156 109.985 26.476 ;
      RECT MASK 1 110.237 26.156 110.317 26.476 ;
      RECT MASK 1 110.569 26.156 110.649 26.476 ;
      RECT MASK 1 110.901 26.156 110.981 26.476 ;
      RECT MASK 1 111.233 26.156 111.313 77.818 ;
      RECT MASK 1 111.565 26.156 111.645 77.818 ;
      RECT MASK 1 111.897 26.156 111.977 77.818 ;
      RECT MASK 1 112.229 26.156 112.309 26.476 ;
      RECT MASK 1 112.561 26.156 112.641 26.476 ;
      RECT MASK 1 112.893 26.156 112.973 26.476 ;
      RECT MASK 1 113.225 26.156 113.305 26.476 ;
      RECT MASK 1 113.557 26.156 113.637 26.476 ;
      RECT MASK 1 113.869 26.175 113.989 31.468 ;
      RECT MASK 1 115.539 26.426 115.659 30.511 ;
      RECT MASK 1 116.261 26.426 116.341 26.728 ;
      RECT MASK 1 116.593 26.426 116.673 26.728 ;
      RECT MASK 1 116.925 26.426 117.005 26.728 ;
      RECT MASK 1 117.257 26.426 117.337 26.728 ;
      RECT MASK 1 117.589 26.426 117.669 26.728 ;
      RECT MASK 1 117.921 26.426 118.001 26.728 ;
      RECT MASK 1 118.253 26.426 118.333 26.728 ;
      RECT MASK 1 118.585 26.426 118.665 26.728 ;
      RECT MASK 1 118.917 26.426 118.997 26.728 ;
      RECT MASK 1 119.249 26.426 119.329 26.728 ;
      RECT MASK 1 119.581 26.426 119.661 26.728 ;
      RECT MASK 1 119.913 26.426 119.993 26.728 ;
      RECT MASK 1 120.245 26.426 120.325 26.728 ;
      RECT MASK 1 120.577 26.426 120.657 26.728 ;
      RECT MASK 1 120.909 26.426 120.989 26.728 ;
      RECT MASK 1 121.241 26.426 121.321 26.728 ;
      RECT MASK 1 121.573 26.426 121.653 26.728 ;
      RECT MASK 1 121.905 26.426 121.985 26.728 ;
      RECT MASK 1 122.237 26.426 122.317 26.728 ;
      RECT MASK 1 122.569 26.426 122.649 26.728 ;
      RECT MASK 1 122.901 26.426 122.981 26.728 ;
      RECT MASK 1 123.233 26.426 123.313 26.728 ;
      RECT MASK 1 123.565 26.426 123.645 26.728 ;
      RECT MASK 1 123.897 26.426 123.977 26.728 ;
      RECT MASK 1 124.229 26.426 124.309 26.728 ;
      RECT MASK 1 124.561 26.426 124.641 26.728 ;
      RECT MASK 1 124.893 26.426 124.973 26.728 ;
      RECT MASK 1 125.225 26.426 125.305 26.728 ;
      RECT MASK 1 125.557 26.426 125.637 26.728 ;
      RECT MASK 1 125.889 26.426 125.969 26.728 ;
      RECT MASK 1 126.221 26.426 126.301 26.728 ;
      RECT MASK 1 126.827 26.426 126.947 30.51 ;
      RECT MASK 1 116.261 27.155 116.341 28.237 ;
      RECT MASK 1 116.593 27.155 116.673 28.237 ;
      RECT MASK 1 116.925 27.155 117.005 28.237 ;
      RECT MASK 1 117.257 27.155 117.337 28.237 ;
      RECT MASK 1 117.589 27.155 117.669 28.237 ;
      RECT MASK 1 117.921 27.155 118.001 28.237 ;
      RECT MASK 1 118.253 27.155 118.333 28.237 ;
      RECT MASK 1 118.585 27.155 118.665 28.237 ;
      RECT MASK 1 118.917 27.155 118.997 28.237 ;
      RECT MASK 1 119.249 27.155 119.329 28.237 ;
      RECT MASK 1 119.581 27.155 119.661 28.237 ;
      RECT MASK 1 119.913 27.155 119.993 28.237 ;
      RECT MASK 1 120.245 27.155 120.325 28.237 ;
      RECT MASK 1 120.577 27.155 120.657 28.237 ;
      RECT MASK 1 120.909 27.155 120.989 28.237 ;
      RECT MASK 1 121.241 27.155 121.321 28.237 ;
      RECT MASK 1 121.573 27.155 121.653 28.237 ;
      RECT MASK 1 121.905 27.155 121.985 28.237 ;
      RECT MASK 1 122.237 27.155 122.317 28.237 ;
      RECT MASK 1 122.569 27.155 122.649 28.237 ;
      RECT MASK 1 122.901 27.155 122.981 28.237 ;
      RECT MASK 1 123.233 27.155 123.313 28.237 ;
      RECT MASK 1 123.565 27.155 123.645 28.237 ;
      RECT MASK 1 123.897 27.155 123.977 28.237 ;
      RECT MASK 1 124.229 27.155 124.309 28.237 ;
      RECT MASK 1 124.561 27.155 124.641 28.237 ;
      RECT MASK 1 124.893 27.155 124.973 28.237 ;
      RECT MASK 1 125.225 27.155 125.305 28.237 ;
      RECT MASK 1 125.557 27.155 125.637 28.237 ;
      RECT MASK 1 125.889 27.155 125.969 28.237 ;
      RECT MASK 1 126.221 27.155 126.301 28.396 ;
      RECT MASK 1 4.681 28.009 4.801 39.191 ;
      RECT MASK 1 5.121 28.009 5.241 39.191 ;
      RECT MASK 1 5.561 28.009 5.681 39.191 ;
      RECT MASK 1 6.001 28.009 6.121 39.191 ;
      RECT MASK 1 6.441 28.009 6.561 39.191 ;
      RECT MASK 1 6.881 28.009 7.001 39.191 ;
      RECT MASK 1 7.321 28.009 7.441 39.191 ;
      RECT MASK 1 7.761 28.009 7.881 39.191 ;
      RECT MASK 1 8.201 28.009 8.321 39.191 ;
      RECT MASK 1 8.641 28.009 8.761 39.191 ;
      RECT MASK 1 9.081 28.009 9.201 39.191 ;
      RECT MASK 1 9.521 28.009 9.641 39.191 ;
      RECT MASK 1 9.961 28.009 10.081 39.191 ;
      RECT MASK 1 10.401 28.009 10.521 39.191 ;
      RECT MASK 1 10.841 28.009 10.961 39.191 ;
      RECT MASK 1 11.299 28.009 11.419 39.191 ;
      RECT MASK 1 11.739 28.009 11.859 39.191 ;
      RECT MASK 1 12.179 28.009 12.299 39.191 ;
      RECT MASK 1 12.619 28.009 12.739 39.191 ;
      RECT MASK 1 13.059 28.009 13.179 39.191 ;
      RECT MASK 1 13.499 28.009 13.619 39.191 ;
      RECT MASK 1 13.939 28.009 14.059 39.191 ;
      RECT MASK 1 14.379 28.009 14.499 39.191 ;
      RECT MASK 1 14.819 28.009 14.939 39.191 ;
      RECT MASK 1 15.259 28.009 15.379 39.191 ;
      RECT MASK 1 15.699 28.009 15.819 39.191 ;
      RECT MASK 1 16.139 28.009 16.259 39.191 ;
      RECT MASK 1 16.579 28.009 16.699 39.191 ;
      RECT MASK 1 17.019 28.009 17.139 39.191 ;
      RECT MASK 1 17.459 28.009 17.579 39.191 ;
      RECT MASK 1 17.917 28.009 18.037 39.191 ;
      RECT MASK 1 18.357 28.009 18.477 39.191 ;
      RECT MASK 1 18.797 28.009 18.917 39.191 ;
      RECT MASK 1 19.237 28.009 19.357 39.191 ;
      RECT MASK 1 19.677 28.009 19.797 39.191 ;
      RECT MASK 1 20.117 28.009 20.237 39.191 ;
      RECT MASK 1 20.557 28.009 20.677 39.191 ;
      RECT MASK 1 20.997 28.009 21.117 39.191 ;
      RECT MASK 1 21.437 28.009 21.557 39.191 ;
      RECT MASK 1 21.877 28.009 21.997 39.191 ;
      RECT MASK 1 22.317 28.009 22.437 39.191 ;
      RECT MASK 1 22.757 28.009 22.877 39.191 ;
      RECT MASK 1 23.197 28.009 23.317 39.191 ;
      RECT MASK 1 23.637 28.009 23.757 39.191 ;
      RECT MASK 1 24.077 28.009 24.197 39.191 ;
      RECT MASK 1 24.535 28.009 24.655 39.191 ;
      RECT MASK 1 24.975 28.009 25.095 39.191 ;
      RECT MASK 1 25.415 28.009 25.535 39.191 ;
      RECT MASK 1 25.855 28.009 25.975 39.191 ;
      RECT MASK 1 26.295 28.009 26.415 39.191 ;
      RECT MASK 1 26.735 28.009 26.855 39.191 ;
      RECT MASK 1 27.175 28.009 27.295 39.191 ;
      RECT MASK 1 27.615 28.009 27.735 39.191 ;
      RECT MASK 1 28.055 28.009 28.175 39.191 ;
      RECT MASK 1 28.495 28.009 28.615 39.191 ;
      RECT MASK 1 28.935 28.009 29.055 39.191 ;
      RECT MASK 1 29.375 28.009 29.495 39.191 ;
      RECT MASK 1 29.815 28.009 29.935 39.191 ;
      RECT MASK 1 30.255 28.009 30.375 39.191 ;
      RECT MASK 1 30.695 28.009 30.815 39.191 ;
      RECT MASK 1 31.153 28.009 31.273 39.191 ;
      RECT MASK 1 31.593 28.009 31.713 39.191 ;
      RECT MASK 1 32.033 28.009 32.153 39.191 ;
      RECT MASK 1 32.473 28.009 32.593 39.191 ;
      RECT MASK 1 32.913 28.009 33.033 39.191 ;
      RECT MASK 1 33.353 28.009 33.473 39.191 ;
      RECT MASK 1 33.793 28.009 33.913 39.191 ;
      RECT MASK 1 34.233 28.009 34.353 39.191 ;
      RECT MASK 1 34.673 28.009 34.793 39.191 ;
      RECT MASK 1 35.113 28.009 35.233 39.191 ;
      RECT MASK 1 35.553 28.009 35.673 39.191 ;
      RECT MASK 1 35.993 28.009 36.113 39.191 ;
      RECT MASK 1 36.433 28.009 36.553 39.191 ;
      RECT MASK 1 36.873 28.009 36.993 39.191 ;
      RECT MASK 1 37.313 28.009 37.433 39.191 ;
      RECT MASK 1 37.771 28.009 37.891 39.191 ;
      RECT MASK 1 38.211 28.009 38.331 39.191 ;
      RECT MASK 1 38.651 28.009 38.771 39.191 ;
      RECT MASK 1 39.091 28.009 39.211 39.191 ;
      RECT MASK 1 39.531 28.009 39.651 39.191 ;
      RECT MASK 1 39.971 28.009 40.091 39.191 ;
      RECT MASK 1 40.411 28.009 40.531 39.191 ;
      RECT MASK 1 40.851 28.009 40.971 39.191 ;
      RECT MASK 1 41.291 28.009 41.411 39.191 ;
      RECT MASK 1 41.731 28.009 41.851 39.191 ;
      RECT MASK 1 42.171 28.009 42.291 39.191 ;
      RECT MASK 1 42.611 28.009 42.731 39.191 ;
      RECT MASK 1 43.051 28.009 43.171 39.191 ;
      RECT MASK 1 43.491 28.009 43.611 39.191 ;
      RECT MASK 1 43.931 28.009 44.051 39.191 ;
      RECT MASK 1 44.389 28.009 44.509 39.191 ;
      RECT MASK 1 44.829 28.009 44.949 39.191 ;
      RECT MASK 1 45.269 28.009 45.389 39.191 ;
      RECT MASK 1 45.709 28.009 45.829 39.191 ;
      RECT MASK 1 46.149 28.009 46.269 39.191 ;
      RECT MASK 1 46.589 28.009 46.709 39.191 ;
      RECT MASK 1 47.029 28.009 47.149 39.191 ;
      RECT MASK 1 47.469 28.009 47.589 39.191 ;
      RECT MASK 1 47.909 28.009 48.029 39.191 ;
      RECT MASK 1 48.349 28.009 48.469 39.191 ;
      RECT MASK 1 48.789 28.009 48.909 39.191 ;
      RECT MASK 1 49.229 28.009 49.349 39.191 ;
      RECT MASK 1 49.669 28.009 49.789 39.191 ;
      RECT MASK 1 50.109 28.009 50.229 39.191 ;
      RECT MASK 1 50.549 28.009 50.669 39.191 ;
      RECT MASK 1 51.007 28.009 51.127 39.191 ;
      RECT MASK 1 51.447 28.009 51.567 39.191 ;
      RECT MASK 1 51.887 28.009 52.007 39.191 ;
      RECT MASK 1 52.327 28.009 52.447 39.191 ;
      RECT MASK 1 52.767 28.009 52.887 39.191 ;
      RECT MASK 1 53.207 28.009 53.327 39.191 ;
      RECT MASK 1 53.647 28.009 53.767 39.191 ;
      RECT MASK 1 54.087 28.009 54.207 39.191 ;
      RECT MASK 1 54.527 28.009 54.647 39.191 ;
      RECT MASK 1 54.967 28.009 55.087 39.191 ;
      RECT MASK 1 55.407 28.009 55.527 39.191 ;
      RECT MASK 1 55.847 28.009 55.967 39.191 ;
      RECT MASK 1 56.287 28.009 56.407 39.191 ;
      RECT MASK 1 56.727 28.009 56.847 39.191 ;
      RECT MASK 1 57.167 28.009 57.287 39.191 ;
      RECT MASK 1 57.625 28.009 57.745 39.191 ;
      RECT MASK 1 58.065 28.009 58.185 39.191 ;
      RECT MASK 1 58.505 28.009 58.625 39.191 ;
      RECT MASK 1 58.945 28.009 59.065 39.191 ;
      RECT MASK 1 59.385 28.009 59.505 39.191 ;
      RECT MASK 1 59.825 28.009 59.945 39.191 ;
      RECT MASK 1 60.265 28.009 60.385 39.191 ;
      RECT MASK 1 60.705 28.009 60.825 39.191 ;
      RECT MASK 1 61.145 28.009 61.265 39.191 ;
      RECT MASK 1 61.585 28.009 61.705 39.191 ;
      RECT MASK 1 62.025 28.009 62.145 39.191 ;
      RECT MASK 1 62.465 28.009 62.585 39.191 ;
      RECT MASK 1 62.905 28.009 63.025 39.191 ;
      RECT MASK 1 63.345 28.009 63.465 39.191 ;
      RECT MASK 1 63.785 28.009 63.905 39.191 ;
      RECT MASK 1 64.243 28.009 64.363 39.191 ;
      RECT MASK 1 64.683 28.009 64.803 39.191 ;
      RECT MASK 1 65.123 28.009 65.243 39.191 ;
      RECT MASK 1 65.563 28.009 65.683 39.191 ;
      RECT MASK 1 66.003 28.009 66.123 39.191 ;
      RECT MASK 1 66.443 28.009 66.563 39.191 ;
      RECT MASK 1 66.883 28.009 67.003 39.191 ;
      RECT MASK 1 67.323 28.009 67.443 39.191 ;
      RECT MASK 1 67.763 28.009 67.883 39.191 ;
      RECT MASK 1 68.203 28.009 68.323 39.191 ;
      RECT MASK 1 68.643 28.009 68.763 39.191 ;
      RECT MASK 1 69.083 28.009 69.203 39.191 ;
      RECT MASK 1 69.523 28.009 69.643 39.191 ;
      RECT MASK 1 69.963 28.009 70.083 39.191 ;
      RECT MASK 1 70.403 28.009 70.523 39.191 ;
      RECT MASK 1 70.861 28.009 70.981 39.191 ;
      RECT MASK 1 71.301 28.009 71.421 39.191 ;
      RECT MASK 1 71.741 28.009 71.861 39.191 ;
      RECT MASK 1 72.181 28.009 72.301 39.191 ;
      RECT MASK 1 72.621 28.009 72.741 39.191 ;
      RECT MASK 1 73.061 28.009 73.181 39.191 ;
      RECT MASK 1 73.501 28.009 73.621 39.191 ;
      RECT MASK 1 73.941 28.009 74.061 39.191 ;
      RECT MASK 1 74.381 28.009 74.501 39.191 ;
      RECT MASK 1 74.821 28.009 74.941 39.191 ;
      RECT MASK 1 75.261 28.009 75.381 39.191 ;
      RECT MASK 1 75.701 28.009 75.821 39.191 ;
      RECT MASK 1 76.141 28.009 76.261 39.191 ;
      RECT MASK 1 76.581 28.009 76.701 39.191 ;
      RECT MASK 1 77.021 28.009 77.141 39.191 ;
      RECT MASK 1 77.479 28.009 77.599 39.191 ;
      RECT MASK 1 77.919 28.009 78.039 39.191 ;
      RECT MASK 1 78.359 28.009 78.479 39.191 ;
      RECT MASK 1 78.799 28.009 78.919 39.191 ;
      RECT MASK 1 79.239 28.009 79.359 39.191 ;
      RECT MASK 1 79.679 28.009 79.799 39.191 ;
      RECT MASK 1 80.119 28.009 80.239 39.191 ;
      RECT MASK 1 80.559 28.009 80.679 39.191 ;
      RECT MASK 1 80.999 28.009 81.119 39.191 ;
      RECT MASK 1 81.439 28.009 81.559 39.191 ;
      RECT MASK 1 81.879 28.009 81.999 39.191 ;
      RECT MASK 1 82.319 28.009 82.439 39.191 ;
      RECT MASK 1 82.759 28.009 82.879 39.191 ;
      RECT MASK 1 83.199 28.009 83.319 39.191 ;
      RECT MASK 1 83.639 28.009 83.759 39.191 ;
      RECT MASK 1 84.097 28.009 84.217 39.191 ;
      RECT MASK 1 84.537 28.009 84.657 39.191 ;
      RECT MASK 1 84.977 28.009 85.097 39.191 ;
      RECT MASK 1 85.417 28.009 85.537 39.191 ;
      RECT MASK 1 85.857 28.009 85.977 39.191 ;
      RECT MASK 1 86.297 28.009 86.417 39.191 ;
      RECT MASK 1 86.737 28.009 86.857 39.191 ;
      RECT MASK 1 87.177 28.009 87.297 39.191 ;
      RECT MASK 1 87.617 28.009 87.737 39.191 ;
      RECT MASK 1 88.057 28.009 88.177 39.191 ;
      RECT MASK 1 88.497 28.009 88.617 39.191 ;
      RECT MASK 1 88.937 28.009 89.057 39.191 ;
      RECT MASK 1 89.377 28.009 89.497 39.191 ;
      RECT MASK 1 89.817 28.009 89.937 39.191 ;
      RECT MASK 1 90.257 28.009 90.377 39.191 ;
      RECT MASK 1 90.715 28.009 90.835 39.191 ;
      RECT MASK 1 91.155 28.009 91.275 39.191 ;
      RECT MASK 1 91.595 28.009 91.715 39.191 ;
      RECT MASK 1 92.035 28.009 92.155 39.191 ;
      RECT MASK 1 92.475 28.009 92.595 39.191 ;
      RECT MASK 1 92.915 28.009 93.035 39.191 ;
      RECT MASK 1 93.355 28.009 93.475 39.191 ;
      RECT MASK 1 93.795 28.009 93.915 39.191 ;
      RECT MASK 1 94.235 28.009 94.355 39.191 ;
      RECT MASK 1 94.675 28.009 94.795 39.191 ;
      RECT MASK 1 95.115 28.009 95.235 39.191 ;
      RECT MASK 1 95.555 28.009 95.675 39.191 ;
      RECT MASK 1 95.995 28.009 96.115 39.191 ;
      RECT MASK 1 96.435 28.009 96.555 39.191 ;
      RECT MASK 1 96.875 28.009 96.995 39.191 ;
      RECT MASK 1 97.333 28.009 97.453 39.191 ;
      RECT MASK 1 97.773 28.009 97.893 39.191 ;
      RECT MASK 1 98.213 28.009 98.333 39.191 ;
      RECT MASK 1 98.653 28.009 98.773 39.191 ;
      RECT MASK 1 99.093 28.009 99.213 39.191 ;
      RECT MASK 1 99.533 28.009 99.653 39.191 ;
      RECT MASK 1 99.973 28.009 100.093 39.191 ;
      RECT MASK 1 100.413 28.009 100.533 39.191 ;
      RECT MASK 1 100.853 28.009 100.973 39.191 ;
      RECT MASK 1 101.293 28.009 101.413 39.191 ;
      RECT MASK 1 101.733 28.009 101.853 39.191 ;
      RECT MASK 1 102.173 28.009 102.293 39.191 ;
      RECT MASK 1 102.613 28.009 102.733 39.191 ;
      RECT MASK 1 103.053 28.009 103.173 39.191 ;
      RECT MASK 1 103.493 28.009 103.613 39.191 ;
      RECT MASK 1 103.951 28.009 104.071 39.191 ;
      RECT MASK 1 104.391 28.009 104.511 39.191 ;
      RECT MASK 1 104.831 28.009 104.951 39.191 ;
      RECT MASK 1 105.271 28.009 105.391 39.191 ;
      RECT MASK 1 105.711 28.009 105.831 39.191 ;
      RECT MASK 1 106.151 28.009 106.271 39.191 ;
      RECT MASK 1 106.591 28.009 106.711 39.191 ;
      RECT MASK 1 107.031 28.009 107.151 39.191 ;
      RECT MASK 1 107.471 28.009 107.591 39.191 ;
      RECT MASK 1 107.911 28.009 108.031 39.191 ;
      RECT MASK 1 108.351 28.009 108.471 39.191 ;
      RECT MASK 1 108.791 28.009 108.911 39.191 ;
      RECT MASK 1 109.231 28.009 109.351 39.191 ;
      RECT MASK 1 109.671 28.009 109.791 39.191 ;
      RECT MASK 1 110.111 28.009 110.231 39.191 ;
      RECT MASK 1 116.261 28.715 116.341 29.797 ;
      RECT MASK 1 116.593 28.715 116.673 29.797 ;
      RECT MASK 1 116.925 28.715 117.005 29.797 ;
      RECT MASK 1 117.257 28.715 117.337 29.797 ;
      RECT MASK 1 117.589 28.715 117.669 29.797 ;
      RECT MASK 1 117.921 28.715 118.001 29.797 ;
      RECT MASK 1 118.253 28.715 118.333 29.797 ;
      RECT MASK 1 118.585 28.715 118.665 29.797 ;
      RECT MASK 1 118.917 28.715 118.997 29.797 ;
      RECT MASK 1 119.249 28.715 119.329 29.797 ;
      RECT MASK 1 119.581 28.715 119.661 29.797 ;
      RECT MASK 1 119.913 28.715 119.993 29.797 ;
      RECT MASK 1 120.245 28.715 120.325 29.797 ;
      RECT MASK 1 120.577 28.715 120.657 29.797 ;
      RECT MASK 1 120.909 28.715 120.989 29.797 ;
      RECT MASK 1 121.241 28.715 121.321 29.797 ;
      RECT MASK 1 121.573 28.715 121.653 29.797 ;
      RECT MASK 1 121.905 28.715 121.985 29.797 ;
      RECT MASK 1 122.237 28.715 122.317 29.797 ;
      RECT MASK 1 122.569 28.715 122.649 29.797 ;
      RECT MASK 1 122.901 28.715 122.981 29.797 ;
      RECT MASK 1 123.233 28.715 123.313 29.797 ;
      RECT MASK 1 123.565 28.715 123.645 29.797 ;
      RECT MASK 1 123.897 28.715 123.977 29.797 ;
      RECT MASK 1 124.229 28.715 124.309 29.797 ;
      RECT MASK 1 124.561 28.715 124.641 29.797 ;
      RECT MASK 1 124.893 28.715 124.973 29.797 ;
      RECT MASK 1 125.225 28.715 125.305 29.797 ;
      RECT MASK 1 125.557 28.715 125.637 29.797 ;
      RECT MASK 1 125.889 28.715 125.969 29.797 ;
      RECT MASK 1 126.221 28.715 126.301 29.797 ;
      RECT MASK 1 116.261 30.206 116.341 30.51 ;
      RECT MASK 1 116.593 30.206 116.673 30.51 ;
      RECT MASK 1 116.925 30.206 117.005 30.51 ;
      RECT MASK 1 117.257 30.206 117.337 30.51 ;
      RECT MASK 1 117.589 30.206 117.669 30.51 ;
      RECT MASK 1 117.921 30.206 118.001 30.51 ;
      RECT MASK 1 118.253 30.206 118.333 30.51 ;
      RECT MASK 1 118.585 30.206 118.665 30.51 ;
      RECT MASK 1 118.917 30.206 118.997 30.51 ;
      RECT MASK 1 119.249 30.206 119.329 30.51 ;
      RECT MASK 1 119.581 30.206 119.661 30.51 ;
      RECT MASK 1 119.913 30.206 119.993 30.51 ;
      RECT MASK 1 120.245 30.206 120.325 30.51 ;
      RECT MASK 1 120.577 30.206 120.657 30.51 ;
      RECT MASK 1 120.909 30.206 120.989 30.51 ;
      RECT MASK 1 121.241 30.206 121.321 30.51 ;
      RECT MASK 1 121.573 30.206 121.653 30.51 ;
      RECT MASK 1 121.905 30.206 121.985 30.51 ;
      RECT MASK 1 122.237 30.206 122.317 30.51 ;
      RECT MASK 1 122.569 30.206 122.649 30.51 ;
      RECT MASK 1 122.901 30.206 122.981 30.51 ;
      RECT MASK 1 123.233 30.206 123.313 30.51 ;
      RECT MASK 1 123.565 30.206 123.645 30.51 ;
      RECT MASK 1 123.897 30.206 123.977 30.51 ;
      RECT MASK 1 124.229 30.206 124.309 30.51 ;
      RECT MASK 1 124.561 30.206 124.641 30.51 ;
      RECT MASK 1 124.893 30.206 124.973 30.51 ;
      RECT MASK 1 125.225 30.206 125.305 30.51 ;
      RECT MASK 1 125.557 30.206 125.637 30.51 ;
      RECT MASK 1 125.889 30.206 125.969 30.51 ;
      RECT MASK 1 126.221 30.206 126.301 30.51 ;
      RECT MASK 1 114.387 31.136 114.467 31.468 ;
      RECT MASK 1 114.719 31.136 114.799 31.468 ;
      RECT MASK 1 115.051 31.136 115.131 31.468 ;
      RECT MASK 1 115.383 31.136 115.463 31.468 ;
      RECT MASK 1 115.549 31.136 115.629 31.468 ;
      RECT MASK 1 115.715 31.136 115.795 31.468 ;
      RECT MASK 1 116.047 31.136 116.127 31.468 ;
      RECT MASK 1 116.213 31.136 116.293 31.468 ;
      RECT MASK 1 116.379 31.136 116.459 31.468 ;
      RECT MASK 1 116.711 31.136 116.791 31.468 ;
      RECT MASK 1 117.043 31.136 117.123 31.468 ;
      RECT MASK 1 117.375 31.136 117.455 31.468 ;
      RECT MASK 1 117.707 31.136 117.787 31.468 ;
      RECT MASK 1 117.873 31.136 117.953 31.468 ;
      RECT MASK 1 118.039 31.136 118.119 31.468 ;
      RECT MASK 1 118.371 31.136 118.451 31.468 ;
      RECT MASK 1 118.537 31.136 118.617 31.468 ;
      RECT MASK 1 118.703 31.136 118.783 31.468 ;
      RECT MASK 1 119.035 31.136 119.115 31.468 ;
      RECT MASK 1 119.367 31.136 119.447 31.468 ;
      RECT MASK 1 119.699 31.136 119.779 31.468 ;
      RECT MASK 1 119.865 31.136 119.945 31.468 ;
      RECT MASK 1 120.031 31.136 120.111 31.468 ;
      RECT MASK 1 120.363 31.136 120.443 31.468 ;
      RECT MASK 1 120.529 31.136 120.609 31.468 ;
      RECT MASK 1 120.695 31.136 120.775 31.468 ;
      RECT MASK 1 121.027 31.136 121.107 31.468 ;
      RECT MASK 1 121.359 31.136 121.439 31.468 ;
      RECT MASK 1 121.691 31.136 121.771 31.468 ;
      RECT MASK 1 122.023 31.136 122.103 31.468 ;
      RECT MASK 1 122.189 31.136 122.269 31.468 ;
      RECT MASK 1 122.355 31.136 122.435 31.468 ;
      RECT MASK 1 122.687 31.136 122.767 31.468 ;
      RECT MASK 1 122.853 31.136 122.933 31.468 ;
      RECT MASK 1 123.019 31.136 123.099 31.468 ;
      RECT MASK 1 123.351 31.136 123.431 31.468 ;
      RECT MASK 1 123.683 31.136 123.763 31.468 ;
      RECT MASK 1 124.015 31.136 124.095 31.468 ;
      RECT MASK 1 124.181 31.136 124.261 31.468 ;
      RECT MASK 1 124.347 31.136 124.427 31.468 ;
      RECT MASK 1 124.513 31.136 124.593 31.468 ;
      RECT MASK 1 124.679 31.136 124.759 31.468 ;
      RECT MASK 1 124.845 31.136 124.925 31.468 ;
      RECT MASK 1 125.011 31.136 125.091 31.468 ;
      RECT MASK 1 125.177 31.136 125.257 31.468 ;
      RECT MASK 1 125.343 31.136 125.423 31.468 ;
      RECT MASK 1 125.675 31.136 125.755 31.468 ;
      RECT MASK 1 126.007 31.136 126.087 31.468 ;
      RECT MASK 1 126.339 31.136 126.419 31.468 ;
      RECT MASK 1 126.505 31.136 126.585 31.468 ;
      RECT MASK 1 126.671 31.136 126.751 31.468 ;
      RECT MASK 1 127.003 31.136 127.083 31.468 ;
      RECT MASK 1 127.169 31.136 127.249 31.468 ;
      RECT MASK 1 127.335 31.136 127.415 31.468 ;
      RECT MASK 1 127.667 31.136 127.747 31.468 ;
      RECT MASK 1 127.999 31.136 128.079 31.468 ;
      RECT MASK 1 128.331 31.136 128.411 31.468 ;
      RECT MASK 1 128.663 31.136 128.743 31.468 ;
      RECT MASK 1 113.2465 32.117 113.3665 32.576 ;
      RECT MASK 1 113.6865 32.117 113.8065 32.576 ;
      RECT MASK 1 114.1265 32.117 114.2465 32.576 ;
      RECT MASK 1 124.3715 32.16 124.4515 71.973 ;
      RECT MASK 1 124.7035 32.16 124.7835 71.973 ;
      RECT MASK 1 125.0355 32.16 125.1155 71.973 ;
      RECT MASK 1 125.3675 32.16 125.4475 71.973 ;
      RECT MASK 1 125.6995 32.16 125.7795 71.973 ;
      RECT MASK 1 126.0315 32.16 126.1115 71.973 ;
      RECT MASK 1 126.3635 32.16 126.4435 71.973 ;
      RECT MASK 1 126.6955 32.16 126.7755 71.973 ;
      RECT MASK 1 127.0275 32.16 127.1075 71.973 ;
      RECT MASK 1 127.3595 32.16 127.4395 71.973 ;
      RECT MASK 1 127.6915 32.16 127.7715 71.973 ;
      RECT MASK 1 112.8065 32.749 112.9265 34.469 ;
      RECT MASK 1 114.5665 32.749 114.6865 34.469 ;
      RECT MASK 1 115.0065 32.749 115.1265 34.469 ;
      RECT MASK 1 115.4465 32.749 115.5665 34.469 ;
      RECT MASK 1 115.8865 32.749 116.0065 34.469 ;
      RECT MASK 1 116.3265 32.749 116.4465 34.469 ;
      RECT MASK 1 117.6465 32.749 117.7665 34.469 ;
      RECT MASK 1 118.0865 32.749 118.2065 34.469 ;
      RECT MASK 1 118.5265 32.749 118.6465 34.469 ;
      RECT MASK 1 118.9665 32.749 119.0865 34.469 ;
      RECT MASK 1 119.4065 32.749 119.5265 34.469 ;
      RECT MASK 1 119.8465 32.749 119.9665 34.469 ;
      RECT MASK 1 120.2865 32.749 120.4065 34.469 ;
      RECT MASK 1 120.7265 32.749 120.8465 34.469 ;
      RECT MASK 1 121.1665 32.749 121.2865 34.469 ;
      RECT MASK 1 121.6065 32.749 121.7265 34.469 ;
      RECT MASK 1 122.0465 32.749 122.1665 34.469 ;
      RECT MASK 1 122.4865 32.749 122.6065 34.469 ;
      RECT MASK 1 122.9265 32.749 123.0465 34.469 ;
      RECT MASK 1 123.3665 32.749 123.4865 34.469 ;
      RECT MASK 1 123.8065 32.749 123.9265 34.469 ;
      RECT MASK 1 112.8065 34.729 112.9265 35.819 ;
      RECT MASK 1 113.2465 34.729 113.3665 35.819 ;
      RECT MASK 1 113.6865 34.729 113.8065 35.819 ;
      RECT MASK 1 114.1265 34.729 114.2465 35.819 ;
      RECT MASK 1 114.5665 34.729 114.6865 35.819 ;
      RECT MASK 1 115.0065 34.729 115.1265 35.819 ;
      RECT MASK 1 115.4465 34.729 115.5665 35.819 ;
      RECT MASK 1 115.8865 34.729 116.0065 35.819 ;
      RECT MASK 1 116.3265 34.729 116.4465 35.819 ;
      RECT MASK 1 117.6465 34.729 117.7665 35.819 ;
      RECT MASK 1 118.0865 34.729 118.2065 35.819 ;
      RECT MASK 1 118.5265 34.729 118.6465 35.819 ;
      RECT MASK 1 118.9665 34.729 119.0865 35.819 ;
      RECT MASK 1 119.4065 34.729 119.5265 35.819 ;
      RECT MASK 1 119.8465 34.729 119.9665 35.819 ;
      RECT MASK 1 120.2865 34.729 120.4065 35.819 ;
      RECT MASK 1 120.7265 34.729 120.8465 35.819 ;
      RECT MASK 1 121.1665 34.729 121.2865 35.819 ;
      RECT MASK 1 121.6065 34.729 121.7265 35.819 ;
      RECT MASK 1 122.0465 34.729 122.1665 35.819 ;
      RECT MASK 1 122.4865 34.729 122.6065 35.819 ;
      RECT MASK 1 122.9265 34.729 123.0465 35.819 ;
      RECT MASK 1 123.3665 34.729 123.4865 35.819 ;
      RECT MASK 1 123.8065 34.729 123.9265 35.819 ;
      RECT MASK 1 112.8065 36.079 112.9265 37.169 ;
      RECT MASK 1 113.2465 36.079 113.3665 37.169 ;
      RECT MASK 1 113.6865 36.079 113.8065 37.169 ;
      RECT MASK 1 114.1265 36.079 114.2465 37.169 ;
      RECT MASK 1 114.5665 36.079 114.6865 37.169 ;
      RECT MASK 1 115.0065 36.079 115.1265 37.169 ;
      RECT MASK 1 115.4465 36.079 115.5665 37.169 ;
      RECT MASK 1 115.8865 36.079 116.0065 37.169 ;
      RECT MASK 1 116.3265 36.079 116.4465 37.169 ;
      RECT MASK 1 117.6465 36.079 117.7665 37.169 ;
      RECT MASK 1 118.0865 36.079 118.2065 37.169 ;
      RECT MASK 1 118.5265 36.079 118.6465 37.169 ;
      RECT MASK 1 118.9665 36.079 119.0865 37.169 ;
      RECT MASK 1 119.4065 36.079 119.5265 37.169 ;
      RECT MASK 1 119.8465 36.079 119.9665 37.169 ;
      RECT MASK 1 120.2865 36.079 120.4065 37.169 ;
      RECT MASK 1 120.7265 36.079 120.8465 37.169 ;
      RECT MASK 1 121.1665 36.079 121.2865 37.169 ;
      RECT MASK 1 121.6065 36.079 121.7265 37.169 ;
      RECT MASK 1 122.0465 36.079 122.1665 37.169 ;
      RECT MASK 1 122.4865 36.079 122.6065 37.169 ;
      RECT MASK 1 122.9265 36.079 123.0465 37.169 ;
      RECT MASK 1 123.3665 36.079 123.4865 37.169 ;
      RECT MASK 1 123.8065 36.079 123.9265 37.169 ;
      RECT MASK 1 112.8065 37.429 112.9265 38.519 ;
      RECT MASK 1 113.2465 37.429 113.3665 38.519 ;
      RECT MASK 1 113.6865 37.429 113.8065 38.519 ;
      RECT MASK 1 114.1265 37.429 114.2465 38.519 ;
      RECT MASK 1 114.5665 37.429 114.6865 38.519 ;
      RECT MASK 1 115.0065 37.429 115.1265 38.519 ;
      RECT MASK 1 115.4465 37.429 115.5665 38.519 ;
      RECT MASK 1 115.8865 37.429 116.0065 38.519 ;
      RECT MASK 1 116.3265 37.429 116.4465 38.519 ;
      RECT MASK 1 117.6465 37.429 117.7665 38.519 ;
      RECT MASK 1 118.0865 37.429 118.2065 38.519 ;
      RECT MASK 1 118.5265 37.429 118.6465 38.519 ;
      RECT MASK 1 118.9665 37.429 119.0865 38.519 ;
      RECT MASK 1 119.4065 37.429 119.5265 38.519 ;
      RECT MASK 1 119.8465 37.429 119.9665 38.519 ;
      RECT MASK 1 120.2865 37.429 120.4065 38.519 ;
      RECT MASK 1 120.7265 37.429 120.8465 38.519 ;
      RECT MASK 1 121.1665 37.429 121.2865 38.519 ;
      RECT MASK 1 121.6065 37.429 121.7265 38.519 ;
      RECT MASK 1 122.0465 37.429 122.1665 38.519 ;
      RECT MASK 1 122.4865 37.429 122.6065 38.519 ;
      RECT MASK 1 122.9265 37.429 123.0465 38.519 ;
      RECT MASK 1 123.3665 37.429 123.4865 38.519 ;
      RECT MASK 1 123.8065 37.429 123.9265 38.519 ;
      RECT MASK 1 112.8065 38.779 112.9265 40.619 ;
      RECT MASK 1 113.2465 38.779 113.3665 40.619 ;
      RECT MASK 1 113.6865 38.779 113.8065 40.619 ;
      RECT MASK 1 114.1265 38.779 114.2465 40.619 ;
      RECT MASK 1 114.5665 38.779 114.6865 40.619 ;
      RECT MASK 1 115.0065 38.779 115.1265 40.619 ;
      RECT MASK 1 115.4465 38.779 115.5665 40.619 ;
      RECT MASK 1 115.8865 38.779 116.0065 40.619 ;
      RECT MASK 1 116.3265 38.779 116.4465 40.619 ;
      RECT MASK 1 117.6465 38.779 117.7665 40.619 ;
      RECT MASK 1 118.0865 38.779 118.2065 40.619 ;
      RECT MASK 1 118.5265 38.779 118.6465 40.619 ;
      RECT MASK 1 118.9665 38.779 119.0865 40.619 ;
      RECT MASK 1 119.4065 38.779 119.5265 40.619 ;
      RECT MASK 1 119.8465 38.779 119.9665 40.619 ;
      RECT MASK 1 120.2865 38.779 120.4065 40.619 ;
      RECT MASK 1 120.7265 38.779 120.8465 40.619 ;
      RECT MASK 1 121.1665 38.779 121.2865 40.619 ;
      RECT MASK 1 121.6065 38.779 121.7265 40.619 ;
      RECT MASK 1 122.0465 38.779 122.1665 40.619 ;
      RECT MASK 1 122.4865 38.779 122.6065 40.619 ;
      RECT MASK 1 122.9265 38.779 123.0465 40.619 ;
      RECT MASK 1 123.3665 38.779 123.4865 40.619 ;
      RECT MASK 1 123.8065 38.779 123.9265 40.619 ;
      RECT MASK 1 4.711 39.36 4.771 39.6 ;
      RECT MASK 1 5.151 39.36 5.211 39.6 ;
      RECT MASK 1 5.591 39.36 5.651 39.6 ;
      RECT MASK 1 6.031 39.36 6.091 39.6 ;
      RECT MASK 1 6.471 39.36 6.531 39.6 ;
      RECT MASK 1 6.911 39.36 6.971 39.6 ;
      RECT MASK 1 7.351 39.36 7.411 39.6 ;
      RECT MASK 1 7.791 39.36 7.851 39.6 ;
      RECT MASK 1 8.231 39.36 8.291 39.6 ;
      RECT MASK 1 8.671 39.36 8.731 39.6 ;
      RECT MASK 1 9.111 39.36 9.171 39.6 ;
      RECT MASK 1 9.551 39.36 9.611 39.6 ;
      RECT MASK 1 9.991 39.36 10.051 39.6 ;
      RECT MASK 1 10.431 39.36 10.491 39.6 ;
      RECT MASK 1 10.871 39.36 10.931 39.6 ;
      RECT MASK 1 11.329 39.36 11.389 39.6 ;
      RECT MASK 1 11.769 39.36 11.829 39.6 ;
      RECT MASK 1 12.209 39.36 12.269 39.6 ;
      RECT MASK 1 12.649 39.36 12.709 39.6 ;
      RECT MASK 1 13.089 39.36 13.149 39.6 ;
      RECT MASK 1 13.529 39.36 13.589 39.6 ;
      RECT MASK 1 13.969 39.36 14.029 39.6 ;
      RECT MASK 1 14.409 39.36 14.469 39.6 ;
      RECT MASK 1 14.849 39.36 14.909 39.6 ;
      RECT MASK 1 15.289 39.36 15.349 39.6 ;
      RECT MASK 1 15.729 39.36 15.789 39.6 ;
      RECT MASK 1 16.169 39.36 16.229 39.6 ;
      RECT MASK 1 16.609 39.36 16.669 39.6 ;
      RECT MASK 1 17.049 39.36 17.109 39.6 ;
      RECT MASK 1 17.489 39.36 17.549 39.6 ;
      RECT MASK 1 17.947 39.36 18.007 39.6 ;
      RECT MASK 1 18.387 39.36 18.447 39.6 ;
      RECT MASK 1 18.827 39.36 18.887 39.6 ;
      RECT MASK 1 19.267 39.36 19.327 39.6 ;
      RECT MASK 1 19.707 39.36 19.767 39.6 ;
      RECT MASK 1 20.147 39.36 20.207 39.6 ;
      RECT MASK 1 20.587 39.36 20.647 39.6 ;
      RECT MASK 1 21.027 39.36 21.087 39.6 ;
      RECT MASK 1 21.467 39.36 21.527 39.6 ;
      RECT MASK 1 21.907 39.36 21.967 39.6 ;
      RECT MASK 1 22.347 39.36 22.407 39.6 ;
      RECT MASK 1 22.787 39.36 22.847 39.6 ;
      RECT MASK 1 23.227 39.36 23.287 39.6 ;
      RECT MASK 1 23.667 39.36 23.727 39.6 ;
      RECT MASK 1 24.107 39.36 24.167 39.6 ;
      RECT MASK 1 24.565 39.36 24.625 39.6 ;
      RECT MASK 1 25.005 39.36 25.065 39.6 ;
      RECT MASK 1 25.445 39.36 25.505 39.6 ;
      RECT MASK 1 25.885 39.36 25.945 39.6 ;
      RECT MASK 1 26.325 39.36 26.385 39.6 ;
      RECT MASK 1 26.765 39.36 26.825 39.6 ;
      RECT MASK 1 27.205 39.36 27.265 39.6 ;
      RECT MASK 1 27.645 39.36 27.705 39.6 ;
      RECT MASK 1 28.085 39.36 28.145 39.6 ;
      RECT MASK 1 28.525 39.36 28.585 39.6 ;
      RECT MASK 1 28.965 39.36 29.025 39.6 ;
      RECT MASK 1 29.405 39.36 29.465 39.6 ;
      RECT MASK 1 29.845 39.36 29.905 39.6 ;
      RECT MASK 1 30.285 39.36 30.345 39.6 ;
      RECT MASK 1 30.725 39.36 30.785 39.6 ;
      RECT MASK 1 31.183 39.36 31.243 39.6 ;
      RECT MASK 1 31.623 39.36 31.683 39.6 ;
      RECT MASK 1 32.063 39.36 32.123 39.6 ;
      RECT MASK 1 32.503 39.36 32.563 39.6 ;
      RECT MASK 1 32.943 39.36 33.003 39.6 ;
      RECT MASK 1 33.383 39.36 33.443 39.6 ;
      RECT MASK 1 33.823 39.36 33.883 39.6 ;
      RECT MASK 1 34.263 39.36 34.323 39.6 ;
      RECT MASK 1 34.703 39.36 34.763 39.6 ;
      RECT MASK 1 35.143 39.36 35.203 39.6 ;
      RECT MASK 1 35.583 39.36 35.643 39.6 ;
      RECT MASK 1 36.023 39.36 36.083 39.6 ;
      RECT MASK 1 36.463 39.36 36.523 39.6 ;
      RECT MASK 1 36.903 39.36 36.963 39.6 ;
      RECT MASK 1 37.343 39.36 37.403 39.6 ;
      RECT MASK 1 37.801 39.36 37.861 39.6 ;
      RECT MASK 1 38.241 39.36 38.301 39.6 ;
      RECT MASK 1 38.681 39.36 38.741 39.6 ;
      RECT MASK 1 39.121 39.36 39.181 39.6 ;
      RECT MASK 1 39.561 39.36 39.621 39.6 ;
      RECT MASK 1 40.001 39.36 40.061 39.6 ;
      RECT MASK 1 40.441 39.36 40.501 39.6 ;
      RECT MASK 1 40.881 39.36 40.941 39.6 ;
      RECT MASK 1 41.321 39.36 41.381 39.6 ;
      RECT MASK 1 41.761 39.36 41.821 39.6 ;
      RECT MASK 1 43.081 39.36 43.141 39.6 ;
      RECT MASK 1 43.521 39.36 43.581 39.6 ;
      RECT MASK 1 43.961 39.36 44.021 39.6 ;
      RECT MASK 1 44.419 39.36 44.479 39.6 ;
      RECT MASK 1 44.859 39.36 44.919 39.6 ;
      RECT MASK 1 45.299 39.36 45.359 39.6 ;
      RECT MASK 1 45.739 39.36 45.799 39.6 ;
      RECT MASK 1 46.179 39.36 46.239 39.6 ;
      RECT MASK 1 46.619 39.36 46.679 39.6 ;
      RECT MASK 1 47.059 39.36 47.119 39.6 ;
      RECT MASK 1 47.499 39.36 47.559 39.6 ;
      RECT MASK 1 47.939 39.36 47.999 39.6 ;
      RECT MASK 1 48.379 39.36 48.439 39.6 ;
      RECT MASK 1 48.819 39.36 48.879 39.6 ;
      RECT MASK 1 49.259 39.36 49.319 39.6 ;
      RECT MASK 1 49.699 39.36 49.759 39.6 ;
      RECT MASK 1 50.139 39.36 50.199 39.6 ;
      RECT MASK 1 50.579 39.36 50.639 39.6 ;
      RECT MASK 1 51.037 39.36 51.097 39.6 ;
      RECT MASK 1 51.477 39.36 51.537 39.6 ;
      RECT MASK 1 51.917 39.36 51.977 39.6 ;
      RECT MASK 1 52.357 39.36 52.417 39.6 ;
      RECT MASK 1 52.797 39.36 52.857 39.6 ;
      RECT MASK 1 53.237 39.36 53.297 39.6 ;
      RECT MASK 1 53.677 39.36 53.737 39.6 ;
      RECT MASK 1 54.117 39.36 54.177 39.6 ;
      RECT MASK 1 54.557 39.36 54.617 39.6 ;
      RECT MASK 1 54.997 39.36 55.057 39.6 ;
      RECT MASK 1 55.437 39.36 55.497 39.6 ;
      RECT MASK 1 55.877 39.36 55.937 39.6 ;
      RECT MASK 1 56.317 39.36 56.377 39.6 ;
      RECT MASK 1 56.757 39.36 56.817 39.6 ;
      RECT MASK 1 57.197 39.36 57.257 39.6 ;
      RECT MASK 1 57.655 39.36 57.715 39.6 ;
      RECT MASK 1 58.095 39.36 58.155 39.6 ;
      RECT MASK 1 58.535 39.36 58.595 39.6 ;
      RECT MASK 1 58.975 39.36 59.035 39.6 ;
      RECT MASK 1 59.415 39.36 59.475 39.6 ;
      RECT MASK 1 59.855 39.36 59.915 39.6 ;
      RECT MASK 1 60.295 39.36 60.355 39.6 ;
      RECT MASK 1 60.735 39.36 60.795 39.6 ;
      RECT MASK 1 61.175 39.36 61.235 39.6 ;
      RECT MASK 1 61.615 39.36 61.675 39.6 ;
      RECT MASK 1 62.055 39.36 62.115 39.6 ;
      RECT MASK 1 62.495 39.36 62.555 39.6 ;
      RECT MASK 1 62.935 39.36 62.995 39.6 ;
      RECT MASK 1 63.375 39.36 63.435 39.6 ;
      RECT MASK 1 63.815 39.36 63.875 39.6 ;
      RECT MASK 1 64.273 39.36 64.333 39.6 ;
      RECT MASK 1 64.713 39.36 64.773 39.6 ;
      RECT MASK 1 65.153 39.36 65.213 39.6 ;
      RECT MASK 1 65.593 39.36 65.653 39.6 ;
      RECT MASK 1 66.033 39.36 66.093 39.6 ;
      RECT MASK 1 66.473 39.36 66.533 39.6 ;
      RECT MASK 1 66.913 39.36 66.973 39.6 ;
      RECT MASK 1 67.353 39.36 67.413 39.6 ;
      RECT MASK 1 67.793 39.36 67.853 39.6 ;
      RECT MASK 1 68.233 39.36 68.293 39.6 ;
      RECT MASK 1 68.673 39.36 68.733 39.6 ;
      RECT MASK 1 69.113 39.36 69.173 39.6 ;
      RECT MASK 1 69.553 39.36 69.613 39.6 ;
      RECT MASK 1 69.993 39.36 70.053 39.6 ;
      RECT MASK 1 70.433 39.36 70.493 39.6 ;
      RECT MASK 1 70.891 39.36 70.951 39.6 ;
      RECT MASK 1 71.331 39.36 71.391 39.6 ;
      RECT MASK 1 71.771 39.36 71.831 39.6 ;
      RECT MASK 1 72.211 39.36 72.271 39.6 ;
      RECT MASK 1 72.651 39.36 72.711 39.6 ;
      RECT MASK 1 73.091 39.36 73.151 39.6 ;
      RECT MASK 1 73.531 39.36 73.591 39.6 ;
      RECT MASK 1 73.971 39.36 74.031 39.6 ;
      RECT MASK 1 74.411 39.36 74.471 39.6 ;
      RECT MASK 1 74.851 39.36 74.911 39.6 ;
      RECT MASK 1 75.291 39.36 75.351 39.6 ;
      RECT MASK 1 75.731 39.36 75.791 39.6 ;
      RECT MASK 1 76.171 39.36 76.231 39.6 ;
      RECT MASK 1 76.611 39.36 76.671 39.6 ;
      RECT MASK 1 77.051 39.36 77.111 39.6 ;
      RECT MASK 1 77.509 39.36 77.569 39.6 ;
      RECT MASK 1 77.949 39.36 78.009 39.6 ;
      RECT MASK 1 78.389 39.36 78.449 39.6 ;
      RECT MASK 1 78.829 39.36 78.889 39.6 ;
      RECT MASK 1 79.269 39.36 79.329 39.6 ;
      RECT MASK 1 79.709 39.36 79.769 39.6 ;
      RECT MASK 1 80.149 39.36 80.209 39.6 ;
      RECT MASK 1 80.589 39.36 80.649 39.6 ;
      RECT MASK 1 81.029 39.36 81.089 39.6 ;
      RECT MASK 1 81.469 39.36 81.529 39.6 ;
      RECT MASK 1 81.909 39.36 81.969 39.6 ;
      RECT MASK 1 82.349 39.36 82.409 39.6 ;
      RECT MASK 1 83.669 39.36 83.729 39.6 ;
      RECT MASK 1 84.127 39.36 84.187 39.6 ;
      RECT MASK 1 84.567 39.36 84.627 39.6 ;
      RECT MASK 1 85.007 39.36 85.067 39.6 ;
      RECT MASK 1 85.447 39.36 85.507 39.6 ;
      RECT MASK 1 85.887 39.36 85.947 39.6 ;
      RECT MASK 1 86.327 39.36 86.387 39.6 ;
      RECT MASK 1 86.767 39.36 86.827 39.6 ;
      RECT MASK 1 87.207 39.36 87.267 39.6 ;
      RECT MASK 1 87.647 39.36 87.707 39.6 ;
      RECT MASK 1 88.087 39.36 88.147 39.6 ;
      RECT MASK 1 88.527 39.36 88.587 39.6 ;
      RECT MASK 1 88.967 39.36 89.027 39.6 ;
      RECT MASK 1 89.407 39.36 89.467 39.6 ;
      RECT MASK 1 89.847 39.36 89.907 39.6 ;
      RECT MASK 1 90.287 39.36 90.347 39.6 ;
      RECT MASK 1 90.745 39.36 90.805 39.6 ;
      RECT MASK 1 91.185 39.36 91.245 39.6 ;
      RECT MASK 1 91.625 39.36 91.685 39.6 ;
      RECT MASK 1 92.065 39.36 92.125 39.6 ;
      RECT MASK 1 92.505 39.36 92.565 39.6 ;
      RECT MASK 1 92.945 39.36 93.005 39.6 ;
      RECT MASK 1 93.385 39.36 93.445 39.6 ;
      RECT MASK 1 93.825 39.36 93.885 39.6 ;
      RECT MASK 1 94.265 39.36 94.325 39.6 ;
      RECT MASK 1 94.705 39.36 94.765 39.6 ;
      RECT MASK 1 95.145 39.36 95.205 39.6 ;
      RECT MASK 1 95.585 39.36 95.645 39.6 ;
      RECT MASK 1 96.025 39.36 96.085 39.6 ;
      RECT MASK 1 96.465 39.36 96.525 39.6 ;
      RECT MASK 1 96.905 39.36 96.965 39.6 ;
      RECT MASK 1 97.363 39.36 97.423 39.6 ;
      RECT MASK 1 97.803 39.36 97.863 39.6 ;
      RECT MASK 1 98.243 39.36 98.303 39.6 ;
      RECT MASK 1 98.683 39.36 98.743 39.6 ;
      RECT MASK 1 99.123 39.36 99.183 39.6 ;
      RECT MASK 1 99.563 39.36 99.623 39.6 ;
      RECT MASK 1 100.003 39.36 100.063 39.6 ;
      RECT MASK 1 100.443 39.36 100.503 39.6 ;
      RECT MASK 1 100.883 39.36 100.943 39.6 ;
      RECT MASK 1 101.323 39.36 101.383 39.6 ;
      RECT MASK 1 101.763 39.36 101.823 39.6 ;
      RECT MASK 1 102.203 39.36 102.263 39.6 ;
      RECT MASK 1 102.643 39.36 102.703 39.6 ;
      RECT MASK 1 103.083 39.36 103.143 39.6 ;
      RECT MASK 1 103.523 39.36 103.583 39.6 ;
      RECT MASK 1 103.981 39.36 104.041 39.6 ;
      RECT MASK 1 104.421 39.36 104.481 39.6 ;
      RECT MASK 1 104.861 39.36 104.921 39.6 ;
      RECT MASK 1 105.301 39.36 105.361 39.6 ;
      RECT MASK 1 105.741 39.36 105.801 39.6 ;
      RECT MASK 1 106.181 39.36 106.241 39.6 ;
      RECT MASK 1 106.621 39.36 106.681 39.6 ;
      RECT MASK 1 107.061 39.36 107.121 39.6 ;
      RECT MASK 1 107.501 39.36 107.561 39.6 ;
      RECT MASK 1 107.941 39.36 108.001 39.6 ;
      RECT MASK 1 108.381 39.36 108.441 39.6 ;
      RECT MASK 1 108.821 39.36 108.881 39.6 ;
      RECT MASK 1 109.261 39.36 109.321 39.6 ;
      RECT MASK 1 109.701 39.36 109.761 39.6 ;
      RECT MASK 1 110.141 39.36 110.201 39.6 ;
      RECT MASK 1 4.711 39.78 4.771 40.02 ;
      RECT MASK 1 5.151 39.78 5.211 40.02 ;
      RECT MASK 1 5.591 39.78 5.651 40.02 ;
      RECT MASK 1 6.031 39.78 6.091 40.02 ;
      RECT MASK 1 6.471 39.78 6.531 40.02 ;
      RECT MASK 1 6.911 39.78 6.971 40.02 ;
      RECT MASK 1 7.351 39.78 7.411 40.02 ;
      RECT MASK 1 7.791 39.78 7.851 40.02 ;
      RECT MASK 1 8.231 39.78 8.291 40.02 ;
      RECT MASK 1 8.671 39.78 8.731 40.02 ;
      RECT MASK 1 9.111 39.78 9.171 40.02 ;
      RECT MASK 1 9.551 39.78 9.611 40.02 ;
      RECT MASK 1 9.991 39.78 10.051 40.02 ;
      RECT MASK 1 10.431 39.78 10.491 40.02 ;
      RECT MASK 1 10.871 39.78 10.931 40.02 ;
      RECT MASK 1 11.329 39.78 11.389 40.02 ;
      RECT MASK 1 11.769 39.78 11.829 40.02 ;
      RECT MASK 1 12.209 39.78 12.269 40.02 ;
      RECT MASK 1 12.649 39.78 12.709 40.02 ;
      RECT MASK 1 13.089 39.78 13.149 40.02 ;
      RECT MASK 1 13.529 39.78 13.589 40.02 ;
      RECT MASK 1 13.969 39.78 14.029 40.02 ;
      RECT MASK 1 14.409 39.78 14.469 40.02 ;
      RECT MASK 1 14.849 39.78 14.909 40.02 ;
      RECT MASK 1 15.289 39.78 15.349 40.02 ;
      RECT MASK 1 15.729 39.78 15.789 40.02 ;
      RECT MASK 1 16.169 39.78 16.229 40.02 ;
      RECT MASK 1 16.609 39.78 16.669 40.02 ;
      RECT MASK 1 17.049 39.78 17.109 40.02 ;
      RECT MASK 1 17.489 39.78 17.549 40.02 ;
      RECT MASK 1 17.947 39.78 18.007 40.02 ;
      RECT MASK 1 18.387 39.78 18.447 40.02 ;
      RECT MASK 1 18.827 39.78 18.887 40.02 ;
      RECT MASK 1 19.267 39.78 19.327 40.02 ;
      RECT MASK 1 19.707 39.78 19.767 40.02 ;
      RECT MASK 1 20.147 39.78 20.207 40.02 ;
      RECT MASK 1 20.587 39.78 20.647 40.02 ;
      RECT MASK 1 21.027 39.78 21.087 40.02 ;
      RECT MASK 1 21.467 39.78 21.527 40.02 ;
      RECT MASK 1 21.907 39.78 21.967 40.02 ;
      RECT MASK 1 22.347 39.78 22.407 40.02 ;
      RECT MASK 1 22.787 39.78 22.847 40.02 ;
      RECT MASK 1 23.227 39.78 23.287 40.02 ;
      RECT MASK 1 23.667 39.78 23.727 40.02 ;
      RECT MASK 1 24.107 39.78 24.167 40.02 ;
      RECT MASK 1 24.565 39.78 24.625 40.02 ;
      RECT MASK 1 25.005 39.78 25.065 40.02 ;
      RECT MASK 1 25.445 39.78 25.505 40.02 ;
      RECT MASK 1 25.885 39.78 25.945 40.02 ;
      RECT MASK 1 26.325 39.78 26.385 40.02 ;
      RECT MASK 1 26.765 39.78 26.825 40.02 ;
      RECT MASK 1 27.205 39.78 27.265 40.02 ;
      RECT MASK 1 27.645 39.78 27.705 40.02 ;
      RECT MASK 1 28.085 39.78 28.145 40.02 ;
      RECT MASK 1 28.525 39.78 28.585 40.02 ;
      RECT MASK 1 28.965 39.78 29.025 40.02 ;
      RECT MASK 1 29.405 39.78 29.465 40.02 ;
      RECT MASK 1 29.845 39.78 29.905 40.02 ;
      RECT MASK 1 30.285 39.78 30.345 40.02 ;
      RECT MASK 1 30.725 39.78 30.785 40.02 ;
      RECT MASK 1 31.183 39.78 31.243 40.02 ;
      RECT MASK 1 31.623 39.78 31.683 40.02 ;
      RECT MASK 1 32.063 39.78 32.123 40.02 ;
      RECT MASK 1 32.503 39.78 32.563 40.02 ;
      RECT MASK 1 32.943 39.78 33.003 40.02 ;
      RECT MASK 1 33.383 39.78 33.443 40.02 ;
      RECT MASK 1 33.823 39.78 33.883 40.02 ;
      RECT MASK 1 34.263 39.78 34.323 40.02 ;
      RECT MASK 1 34.703 39.78 34.763 40.02 ;
      RECT MASK 1 35.143 39.78 35.203 40.02 ;
      RECT MASK 1 35.583 39.78 35.643 40.02 ;
      RECT MASK 1 36.023 39.78 36.083 40.02 ;
      RECT MASK 1 36.463 39.78 36.523 40.02 ;
      RECT MASK 1 36.903 39.78 36.963 40.02 ;
      RECT MASK 1 37.343 39.78 37.403 40.02 ;
      RECT MASK 1 37.801 39.78 37.861 40.02 ;
      RECT MASK 1 38.241 39.78 38.301 40.02 ;
      RECT MASK 1 38.681 39.78 38.741 40.02 ;
      RECT MASK 1 39.121 39.78 39.181 40.02 ;
      RECT MASK 1 39.561 39.78 39.621 40.02 ;
      RECT MASK 1 40.001 39.78 40.061 40.02 ;
      RECT MASK 1 40.441 39.78 40.501 40.02 ;
      RECT MASK 1 40.881 39.78 40.941 40.02 ;
      RECT MASK 1 41.321 39.78 41.381 40.02 ;
      RECT MASK 1 41.761 39.78 41.821 40.02 ;
      RECT MASK 1 43.081 39.78 43.141 40.02 ;
      RECT MASK 1 43.521 39.78 43.581 40.02 ;
      RECT MASK 1 43.961 39.78 44.021 40.02 ;
      RECT MASK 1 44.419 39.78 44.479 40.02 ;
      RECT MASK 1 44.859 39.78 44.919 40.02 ;
      RECT MASK 1 45.299 39.78 45.359 40.02 ;
      RECT MASK 1 45.739 39.78 45.799 40.02 ;
      RECT MASK 1 46.179 39.78 46.239 40.02 ;
      RECT MASK 1 46.619 39.78 46.679 40.02 ;
      RECT MASK 1 47.059 39.78 47.119 40.02 ;
      RECT MASK 1 47.499 39.78 47.559 40.02 ;
      RECT MASK 1 47.939 39.78 47.999 40.02 ;
      RECT MASK 1 48.379 39.78 48.439 40.02 ;
      RECT MASK 1 48.819 39.78 48.879 40.02 ;
      RECT MASK 1 49.259 39.78 49.319 40.02 ;
      RECT MASK 1 49.699 39.78 49.759 40.02 ;
      RECT MASK 1 50.139 39.78 50.199 40.02 ;
      RECT MASK 1 50.579 39.78 50.639 40.02 ;
      RECT MASK 1 51.037 39.78 51.097 40.02 ;
      RECT MASK 1 51.477 39.78 51.537 40.02 ;
      RECT MASK 1 51.917 39.78 51.977 40.02 ;
      RECT MASK 1 52.357 39.78 52.417 40.02 ;
      RECT MASK 1 52.797 39.78 52.857 40.02 ;
      RECT MASK 1 53.237 39.78 53.297 40.02 ;
      RECT MASK 1 53.677 39.78 53.737 40.02 ;
      RECT MASK 1 54.117 39.78 54.177 40.02 ;
      RECT MASK 1 54.557 39.78 54.617 40.02 ;
      RECT MASK 1 54.997 39.78 55.057 40.02 ;
      RECT MASK 1 55.437 39.78 55.497 40.02 ;
      RECT MASK 1 55.877 39.78 55.937 40.02 ;
      RECT MASK 1 56.317 39.78 56.377 40.02 ;
      RECT MASK 1 56.757 39.78 56.817 40.02 ;
      RECT MASK 1 57.197 39.78 57.257 40.02 ;
      RECT MASK 1 57.655 39.78 57.715 40.02 ;
      RECT MASK 1 58.095 39.78 58.155 40.02 ;
      RECT MASK 1 58.535 39.78 58.595 40.02 ;
      RECT MASK 1 58.975 39.78 59.035 40.02 ;
      RECT MASK 1 59.415 39.78 59.475 40.02 ;
      RECT MASK 1 59.855 39.78 59.915 40.02 ;
      RECT MASK 1 60.295 39.78 60.355 40.02 ;
      RECT MASK 1 60.735 39.78 60.795 40.02 ;
      RECT MASK 1 61.175 39.78 61.235 40.02 ;
      RECT MASK 1 61.615 39.78 61.675 40.02 ;
      RECT MASK 1 62.055 39.78 62.115 40.02 ;
      RECT MASK 1 62.495 39.78 62.555 40.02 ;
      RECT MASK 1 62.935 39.78 62.995 40.02 ;
      RECT MASK 1 63.375 39.78 63.435 40.02 ;
      RECT MASK 1 63.815 39.78 63.875 40.02 ;
      RECT MASK 1 64.273 39.78 64.333 40.02 ;
      RECT MASK 1 64.713 39.78 64.773 40.02 ;
      RECT MASK 1 65.153 39.78 65.213 40.02 ;
      RECT MASK 1 65.593 39.78 65.653 40.02 ;
      RECT MASK 1 66.033 39.78 66.093 40.02 ;
      RECT MASK 1 66.473 39.78 66.533 40.02 ;
      RECT MASK 1 66.913 39.78 66.973 40.02 ;
      RECT MASK 1 67.353 39.78 67.413 40.02 ;
      RECT MASK 1 67.793 39.78 67.853 40.02 ;
      RECT MASK 1 68.233 39.78 68.293 40.02 ;
      RECT MASK 1 68.673 39.78 68.733 40.02 ;
      RECT MASK 1 69.113 39.78 69.173 40.02 ;
      RECT MASK 1 69.553 39.78 69.613 40.02 ;
      RECT MASK 1 69.993 39.78 70.053 40.02 ;
      RECT MASK 1 70.433 39.78 70.493 40.02 ;
      RECT MASK 1 70.891 39.78 70.951 40.02 ;
      RECT MASK 1 71.331 39.78 71.391 40.02 ;
      RECT MASK 1 71.771 39.78 71.831 40.02 ;
      RECT MASK 1 72.211 39.78 72.271 40.02 ;
      RECT MASK 1 72.651 39.78 72.711 40.02 ;
      RECT MASK 1 73.091 39.78 73.151 40.02 ;
      RECT MASK 1 73.531 39.78 73.591 40.02 ;
      RECT MASK 1 73.971 39.78 74.031 40.02 ;
      RECT MASK 1 74.411 39.78 74.471 40.02 ;
      RECT MASK 1 74.851 39.78 74.911 40.02 ;
      RECT MASK 1 75.291 39.78 75.351 40.02 ;
      RECT MASK 1 75.731 39.78 75.791 40.02 ;
      RECT MASK 1 76.171 39.78 76.231 40.02 ;
      RECT MASK 1 76.611 39.78 76.671 40.02 ;
      RECT MASK 1 77.051 39.78 77.111 40.02 ;
      RECT MASK 1 77.509 39.78 77.569 40.02 ;
      RECT MASK 1 77.949 39.78 78.009 40.02 ;
      RECT MASK 1 78.389 39.78 78.449 40.02 ;
      RECT MASK 1 78.829 39.78 78.889 40.02 ;
      RECT MASK 1 79.269 39.78 79.329 40.02 ;
      RECT MASK 1 79.709 39.78 79.769 40.02 ;
      RECT MASK 1 80.149 39.78 80.209 40.02 ;
      RECT MASK 1 80.589 39.78 80.649 40.02 ;
      RECT MASK 1 81.029 39.78 81.089 40.02 ;
      RECT MASK 1 81.469 39.78 81.529 40.02 ;
      RECT MASK 1 81.909 39.78 81.969 40.02 ;
      RECT MASK 1 82.349 39.78 82.409 40.02 ;
      RECT MASK 1 83.669 39.78 83.729 40.02 ;
      RECT MASK 1 84.127 39.78 84.187 40.02 ;
      RECT MASK 1 84.567 39.78 84.627 40.02 ;
      RECT MASK 1 85.007 39.78 85.067 40.02 ;
      RECT MASK 1 85.447 39.78 85.507 40.02 ;
      RECT MASK 1 85.887 39.78 85.947 40.02 ;
      RECT MASK 1 86.327 39.78 86.387 40.02 ;
      RECT MASK 1 86.767 39.78 86.827 40.02 ;
      RECT MASK 1 87.207 39.78 87.267 40.02 ;
      RECT MASK 1 87.647 39.78 87.707 40.02 ;
      RECT MASK 1 88.087 39.78 88.147 40.02 ;
      RECT MASK 1 88.527 39.78 88.587 40.02 ;
      RECT MASK 1 88.967 39.78 89.027 40.02 ;
      RECT MASK 1 89.407 39.78 89.467 40.02 ;
      RECT MASK 1 89.847 39.78 89.907 40.02 ;
      RECT MASK 1 90.287 39.78 90.347 40.02 ;
      RECT MASK 1 90.745 39.78 90.805 40.02 ;
      RECT MASK 1 91.185 39.78 91.245 40.02 ;
      RECT MASK 1 91.625 39.78 91.685 40.02 ;
      RECT MASK 1 92.065 39.78 92.125 40.02 ;
      RECT MASK 1 92.505 39.78 92.565 40.02 ;
      RECT MASK 1 92.945 39.78 93.005 40.02 ;
      RECT MASK 1 93.385 39.78 93.445 40.02 ;
      RECT MASK 1 93.825 39.78 93.885 40.02 ;
      RECT MASK 1 94.265 39.78 94.325 40.02 ;
      RECT MASK 1 94.705 39.78 94.765 40.02 ;
      RECT MASK 1 95.145 39.78 95.205 40.02 ;
      RECT MASK 1 95.585 39.78 95.645 40.02 ;
      RECT MASK 1 96.025 39.78 96.085 40.02 ;
      RECT MASK 1 96.465 39.78 96.525 40.02 ;
      RECT MASK 1 96.905 39.78 96.965 40.02 ;
      RECT MASK 1 97.363 39.78 97.423 40.02 ;
      RECT MASK 1 97.803 39.78 97.863 40.02 ;
      RECT MASK 1 98.243 39.78 98.303 40.02 ;
      RECT MASK 1 98.683 39.78 98.743 40.02 ;
      RECT MASK 1 99.123 39.78 99.183 40.02 ;
      RECT MASK 1 99.563 39.78 99.623 40.02 ;
      RECT MASK 1 100.003 39.78 100.063 40.02 ;
      RECT MASK 1 100.443 39.78 100.503 40.02 ;
      RECT MASK 1 100.883 39.78 100.943 40.02 ;
      RECT MASK 1 101.323 39.78 101.383 40.02 ;
      RECT MASK 1 101.763 39.78 101.823 40.02 ;
      RECT MASK 1 102.203 39.78 102.263 40.02 ;
      RECT MASK 1 102.643 39.78 102.703 40.02 ;
      RECT MASK 1 103.083 39.78 103.143 40.02 ;
      RECT MASK 1 103.523 39.78 103.583 40.02 ;
      RECT MASK 1 103.981 39.78 104.041 40.02 ;
      RECT MASK 1 104.421 39.78 104.481 40.02 ;
      RECT MASK 1 104.861 39.78 104.921 40.02 ;
      RECT MASK 1 105.301 39.78 105.361 40.02 ;
      RECT MASK 1 105.741 39.78 105.801 40.02 ;
      RECT MASK 1 106.181 39.78 106.241 40.02 ;
      RECT MASK 1 106.621 39.78 106.681 40.02 ;
      RECT MASK 1 107.061 39.78 107.121 40.02 ;
      RECT MASK 1 107.501 39.78 107.561 40.02 ;
      RECT MASK 1 107.941 39.78 108.001 40.02 ;
      RECT MASK 1 108.381 39.78 108.441 40.02 ;
      RECT MASK 1 108.821 39.78 108.881 40.02 ;
      RECT MASK 1 109.261 39.78 109.321 40.02 ;
      RECT MASK 1 109.701 39.78 109.761 40.02 ;
      RECT MASK 1 110.141 39.78 110.201 40.02 ;
      RECT MASK 1 4.681 40.219 4.801 51.431 ;
      RECT MASK 1 5.121 40.219 5.241 51.431 ;
      RECT MASK 1 5.561 40.219 5.681 51.431 ;
      RECT MASK 1 6.001 40.219 6.121 51.431 ;
      RECT MASK 1 6.441 40.219 6.561 51.431 ;
      RECT MASK 1 6.881 40.219 7.001 51.431 ;
      RECT MASK 1 7.321 40.219 7.441 51.431 ;
      RECT MASK 1 7.761 40.219 7.881 51.431 ;
      RECT MASK 1 8.201 40.219 8.321 51.431 ;
      RECT MASK 1 8.641 40.219 8.761 51.431 ;
      RECT MASK 1 9.081 40.219 9.201 51.431 ;
      RECT MASK 1 9.521 40.219 9.641 51.431 ;
      RECT MASK 1 9.961 40.219 10.081 51.431 ;
      RECT MASK 1 10.401 40.219 10.521 51.431 ;
      RECT MASK 1 10.841 40.219 10.961 51.431 ;
      RECT MASK 1 11.299 40.219 11.419 51.431 ;
      RECT MASK 1 11.739 40.219 11.859 51.431 ;
      RECT MASK 1 12.179 40.219 12.299 51.431 ;
      RECT MASK 1 12.619 40.219 12.739 51.431 ;
      RECT MASK 1 13.059 40.219 13.179 51.431 ;
      RECT MASK 1 13.499 40.219 13.619 51.431 ;
      RECT MASK 1 13.939 40.219 14.059 51.431 ;
      RECT MASK 1 14.379 40.219 14.499 51.431 ;
      RECT MASK 1 14.819 40.219 14.939 51.431 ;
      RECT MASK 1 15.259 40.219 15.379 51.431 ;
      RECT MASK 1 15.699 40.219 15.819 51.431 ;
      RECT MASK 1 16.139 40.219 16.259 51.431 ;
      RECT MASK 1 16.579 40.219 16.699 51.431 ;
      RECT MASK 1 17.019 40.219 17.139 51.431 ;
      RECT MASK 1 17.459 40.219 17.579 51.431 ;
      RECT MASK 1 17.917 40.219 18.037 51.431 ;
      RECT MASK 1 18.357 40.219 18.477 51.431 ;
      RECT MASK 1 18.797 40.219 18.917 51.431 ;
      RECT MASK 1 19.237 40.219 19.357 51.431 ;
      RECT MASK 1 19.677 40.219 19.797 51.431 ;
      RECT MASK 1 20.117 40.219 20.237 51.431 ;
      RECT MASK 1 20.557 40.219 20.677 51.431 ;
      RECT MASK 1 20.997 40.219 21.117 51.431 ;
      RECT MASK 1 21.437 40.219 21.557 51.431 ;
      RECT MASK 1 21.877 40.219 21.997 51.431 ;
      RECT MASK 1 22.317 40.219 22.437 51.431 ;
      RECT MASK 1 22.757 40.219 22.877 51.431 ;
      RECT MASK 1 23.197 40.219 23.317 51.431 ;
      RECT MASK 1 23.637 40.219 23.757 51.431 ;
      RECT MASK 1 24.077 40.219 24.197 51.431 ;
      RECT MASK 1 24.535 40.219 24.655 51.431 ;
      RECT MASK 1 24.975 40.219 25.095 51.431 ;
      RECT MASK 1 25.415 40.219 25.535 51.431 ;
      RECT MASK 1 25.855 40.219 25.975 51.431 ;
      RECT MASK 1 26.295 40.219 26.415 51.431 ;
      RECT MASK 1 26.735 40.219 26.855 51.431 ;
      RECT MASK 1 27.175 40.219 27.295 51.431 ;
      RECT MASK 1 27.615 40.219 27.735 51.431 ;
      RECT MASK 1 28.055 40.219 28.175 51.431 ;
      RECT MASK 1 28.495 40.219 28.615 51.431 ;
      RECT MASK 1 28.935 40.219 29.055 51.431 ;
      RECT MASK 1 29.375 40.219 29.495 51.431 ;
      RECT MASK 1 29.815 40.219 29.935 51.431 ;
      RECT MASK 1 30.255 40.219 30.375 51.431 ;
      RECT MASK 1 30.695 40.219 30.815 51.431 ;
      RECT MASK 1 31.153 40.219 31.273 51.431 ;
      RECT MASK 1 31.593 40.219 31.713 51.431 ;
      RECT MASK 1 32.033 40.219 32.153 51.431 ;
      RECT MASK 1 32.473 40.219 32.593 51.431 ;
      RECT MASK 1 32.913 40.219 33.033 51.431 ;
      RECT MASK 1 33.353 40.219 33.473 51.431 ;
      RECT MASK 1 33.793 40.219 33.913 51.431 ;
      RECT MASK 1 34.233 40.219 34.353 51.431 ;
      RECT MASK 1 34.673 40.219 34.793 51.431 ;
      RECT MASK 1 35.113 40.219 35.233 51.431 ;
      RECT MASK 1 35.553 40.219 35.673 51.431 ;
      RECT MASK 1 35.993 40.219 36.113 51.431 ;
      RECT MASK 1 36.433 40.219 36.553 51.431 ;
      RECT MASK 1 36.873 40.219 36.993 51.431 ;
      RECT MASK 1 37.313 40.219 37.433 51.431 ;
      RECT MASK 1 37.771 40.219 37.891 51.431 ;
      RECT MASK 1 38.211 40.219 38.331 51.431 ;
      RECT MASK 1 38.651 40.219 38.771 51.431 ;
      RECT MASK 1 39.091 40.219 39.211 51.431 ;
      RECT MASK 1 39.531 40.219 39.651 51.431 ;
      RECT MASK 1 39.971 40.219 40.091 51.431 ;
      RECT MASK 1 40.411 40.219 40.531 51.431 ;
      RECT MASK 1 40.851 40.219 40.971 51.431 ;
      RECT MASK 1 41.291 40.219 41.411 51.431 ;
      RECT MASK 1 41.731 40.219 41.851 51.431 ;
      RECT MASK 1 42.171 40.219 42.291 51.431 ;
      RECT MASK 1 42.611 40.219 42.731 51.431 ;
      RECT MASK 1 43.051 40.219 43.171 51.431 ;
      RECT MASK 1 43.491 40.219 43.611 51.431 ;
      RECT MASK 1 43.931 40.219 44.051 51.431 ;
      RECT MASK 1 44.389 40.219 44.509 51.431 ;
      RECT MASK 1 44.829 40.219 44.949 51.431 ;
      RECT MASK 1 45.269 40.219 45.389 51.431 ;
      RECT MASK 1 45.709 40.219 45.829 51.431 ;
      RECT MASK 1 46.149 40.219 46.269 51.431 ;
      RECT MASK 1 46.589 40.219 46.709 51.431 ;
      RECT MASK 1 47.029 40.219 47.149 51.431 ;
      RECT MASK 1 47.469 40.219 47.589 51.431 ;
      RECT MASK 1 47.909 40.219 48.029 51.431 ;
      RECT MASK 1 48.349 40.219 48.469 51.431 ;
      RECT MASK 1 48.789 40.219 48.909 51.431 ;
      RECT MASK 1 49.229 40.219 49.349 51.431 ;
      RECT MASK 1 49.669 40.219 49.789 51.431 ;
      RECT MASK 1 50.109 40.219 50.229 51.431 ;
      RECT MASK 1 50.549 40.219 50.669 51.431 ;
      RECT MASK 1 51.007 40.219 51.127 51.431 ;
      RECT MASK 1 51.447 40.219 51.567 51.431 ;
      RECT MASK 1 51.887 40.219 52.007 51.431 ;
      RECT MASK 1 52.327 40.219 52.447 51.431 ;
      RECT MASK 1 52.767 40.219 52.887 51.431 ;
      RECT MASK 1 53.207 40.219 53.327 51.431 ;
      RECT MASK 1 53.647 40.219 53.767 51.431 ;
      RECT MASK 1 54.087 40.219 54.207 51.431 ;
      RECT MASK 1 54.527 40.219 54.647 51.431 ;
      RECT MASK 1 54.967 40.219 55.087 51.431 ;
      RECT MASK 1 55.407 40.219 55.527 51.431 ;
      RECT MASK 1 55.847 40.219 55.967 51.431 ;
      RECT MASK 1 56.287 40.219 56.407 51.431 ;
      RECT MASK 1 56.727 40.219 56.847 51.431 ;
      RECT MASK 1 57.167 40.219 57.287 51.431 ;
      RECT MASK 1 57.625 40.219 57.745 51.431 ;
      RECT MASK 1 58.065 40.219 58.185 51.431 ;
      RECT MASK 1 58.505 40.219 58.625 51.431 ;
      RECT MASK 1 58.945 40.219 59.065 51.431 ;
      RECT MASK 1 59.385 40.219 59.505 51.431 ;
      RECT MASK 1 59.825 40.219 59.945 51.431 ;
      RECT MASK 1 60.265 40.219 60.385 51.431 ;
      RECT MASK 1 60.705 40.219 60.825 51.431 ;
      RECT MASK 1 61.145 40.219 61.265 51.431 ;
      RECT MASK 1 61.585 40.219 61.705 51.431 ;
      RECT MASK 1 62.025 40.219 62.145 51.431 ;
      RECT MASK 1 62.465 40.219 62.585 51.431 ;
      RECT MASK 1 62.905 40.219 63.025 51.431 ;
      RECT MASK 1 63.345 40.219 63.465 51.431 ;
      RECT MASK 1 63.785 40.219 63.905 51.431 ;
      RECT MASK 1 64.243 40.219 64.363 51.431 ;
      RECT MASK 1 64.683 40.219 64.803 51.431 ;
      RECT MASK 1 65.123 40.219 65.243 51.431 ;
      RECT MASK 1 65.563 40.219 65.683 51.431 ;
      RECT MASK 1 66.003 40.219 66.123 51.431 ;
      RECT MASK 1 66.443 40.219 66.563 51.431 ;
      RECT MASK 1 66.883 40.219 67.003 51.431 ;
      RECT MASK 1 67.323 40.219 67.443 51.431 ;
      RECT MASK 1 67.763 40.219 67.883 51.431 ;
      RECT MASK 1 68.203 40.219 68.323 51.431 ;
      RECT MASK 1 68.643 40.219 68.763 51.431 ;
      RECT MASK 1 69.083 40.219 69.203 51.431 ;
      RECT MASK 1 69.523 40.219 69.643 51.431 ;
      RECT MASK 1 69.963 40.219 70.083 51.431 ;
      RECT MASK 1 70.403 40.219 70.523 51.431 ;
      RECT MASK 1 70.861 40.219 70.981 51.431 ;
      RECT MASK 1 71.301 40.219 71.421 51.431 ;
      RECT MASK 1 71.741 40.219 71.861 51.431 ;
      RECT MASK 1 72.181 40.219 72.301 51.431 ;
      RECT MASK 1 72.621 40.219 72.741 51.431 ;
      RECT MASK 1 73.061 40.219 73.181 51.431 ;
      RECT MASK 1 73.501 40.219 73.621 51.431 ;
      RECT MASK 1 73.941 40.219 74.061 51.431 ;
      RECT MASK 1 74.381 40.219 74.501 51.431 ;
      RECT MASK 1 74.821 40.219 74.941 51.431 ;
      RECT MASK 1 75.261 40.219 75.381 51.431 ;
      RECT MASK 1 75.701 40.219 75.821 51.431 ;
      RECT MASK 1 76.141 40.219 76.261 51.431 ;
      RECT MASK 1 76.581 40.219 76.701 51.431 ;
      RECT MASK 1 77.021 40.219 77.141 51.431 ;
      RECT MASK 1 77.479 40.219 77.599 51.431 ;
      RECT MASK 1 77.919 40.219 78.039 51.431 ;
      RECT MASK 1 78.359 40.219 78.479 51.431 ;
      RECT MASK 1 78.799 40.219 78.919 51.431 ;
      RECT MASK 1 79.239 40.219 79.359 51.431 ;
      RECT MASK 1 79.679 40.219 79.799 51.431 ;
      RECT MASK 1 80.119 40.219 80.239 51.431 ;
      RECT MASK 1 80.559 40.219 80.679 51.431 ;
      RECT MASK 1 80.999 40.219 81.119 51.431 ;
      RECT MASK 1 81.439 40.219 81.559 51.431 ;
      RECT MASK 1 81.879 40.219 81.999 51.431 ;
      RECT MASK 1 82.319 40.219 82.439 51.431 ;
      RECT MASK 1 82.759 40.219 82.879 51.431 ;
      RECT MASK 1 83.199 40.219 83.319 51.431 ;
      RECT MASK 1 83.639 40.219 83.759 51.431 ;
      RECT MASK 1 84.097 40.219 84.217 51.431 ;
      RECT MASK 1 84.537 40.219 84.657 51.431 ;
      RECT MASK 1 84.977 40.219 85.097 51.431 ;
      RECT MASK 1 85.417 40.219 85.537 51.431 ;
      RECT MASK 1 85.857 40.219 85.977 51.431 ;
      RECT MASK 1 86.297 40.219 86.417 51.431 ;
      RECT MASK 1 86.737 40.219 86.857 51.431 ;
      RECT MASK 1 87.177 40.219 87.297 51.431 ;
      RECT MASK 1 87.617 40.219 87.737 51.431 ;
      RECT MASK 1 88.057 40.219 88.177 51.431 ;
      RECT MASK 1 88.497 40.219 88.617 51.431 ;
      RECT MASK 1 88.937 40.219 89.057 51.431 ;
      RECT MASK 1 89.377 40.219 89.497 51.431 ;
      RECT MASK 1 89.817 40.219 89.937 51.431 ;
      RECT MASK 1 90.257 40.219 90.377 51.431 ;
      RECT MASK 1 90.715 40.219 90.835 51.431 ;
      RECT MASK 1 91.155 40.219 91.275 51.431 ;
      RECT MASK 1 91.595 40.219 91.715 51.431 ;
      RECT MASK 1 92.035 40.219 92.155 51.431 ;
      RECT MASK 1 92.475 40.219 92.595 51.431 ;
      RECT MASK 1 92.915 40.219 93.035 51.431 ;
      RECT MASK 1 93.355 40.219 93.475 51.431 ;
      RECT MASK 1 93.795 40.219 93.915 51.431 ;
      RECT MASK 1 94.235 40.219 94.355 51.431 ;
      RECT MASK 1 94.675 40.219 94.795 51.431 ;
      RECT MASK 1 95.115 40.219 95.235 51.431 ;
      RECT MASK 1 95.555 40.219 95.675 51.431 ;
      RECT MASK 1 95.995 40.219 96.115 51.431 ;
      RECT MASK 1 96.435 40.219 96.555 51.431 ;
      RECT MASK 1 96.875 40.219 96.995 51.431 ;
      RECT MASK 1 97.333 40.219 97.453 51.431 ;
      RECT MASK 1 97.773 40.219 97.893 51.431 ;
      RECT MASK 1 98.213 40.219 98.333 51.431 ;
      RECT MASK 1 98.653 40.219 98.773 51.431 ;
      RECT MASK 1 99.093 40.219 99.213 51.431 ;
      RECT MASK 1 99.533 40.219 99.653 51.431 ;
      RECT MASK 1 99.973 40.219 100.093 51.431 ;
      RECT MASK 1 100.413 40.219 100.533 51.431 ;
      RECT MASK 1 100.853 40.219 100.973 51.431 ;
      RECT MASK 1 101.293 40.219 101.413 51.431 ;
      RECT MASK 1 101.733 40.219 101.853 51.431 ;
      RECT MASK 1 102.173 40.219 102.293 51.431 ;
      RECT MASK 1 102.613 40.219 102.733 51.431 ;
      RECT MASK 1 103.053 40.219 103.173 51.431 ;
      RECT MASK 1 103.493 40.219 103.613 51.431 ;
      RECT MASK 1 103.951 40.219 104.071 51.431 ;
      RECT MASK 1 104.391 40.219 104.511 51.431 ;
      RECT MASK 1 104.831 40.219 104.951 51.431 ;
      RECT MASK 1 105.271 40.219 105.391 51.431 ;
      RECT MASK 1 105.711 40.219 105.831 51.431 ;
      RECT MASK 1 106.151 40.219 106.271 51.431 ;
      RECT MASK 1 106.591 40.219 106.711 51.431 ;
      RECT MASK 1 107.031 40.219 107.151 51.431 ;
      RECT MASK 1 107.471 40.219 107.591 51.431 ;
      RECT MASK 1 107.911 40.219 108.031 51.431 ;
      RECT MASK 1 108.351 40.219 108.471 51.431 ;
      RECT MASK 1 108.791 40.219 108.911 51.431 ;
      RECT MASK 1 109.231 40.219 109.351 51.431 ;
      RECT MASK 1 109.671 40.219 109.791 51.431 ;
      RECT MASK 1 110.111 40.219 110.231 51.431 ;
      RECT MASK 1 112.8065 40.879 112.9265 41.939 ;
      RECT MASK 1 113.2465 40.879 113.3665 41.939 ;
      RECT MASK 1 113.6865 40.879 113.8065 41.939 ;
      RECT MASK 1 114.1265 40.879 114.2465 41.939 ;
      RECT MASK 1 114.5665 40.879 114.6865 41.939 ;
      RECT MASK 1 115.0065 40.879 115.1265 41.939 ;
      RECT MASK 1 115.4465 40.879 115.5665 41.939 ;
      RECT MASK 1 115.8865 40.879 116.0065 41.939 ;
      RECT MASK 1 116.3265 40.879 116.4465 41.939 ;
      RECT MASK 1 117.6465 40.879 117.7665 41.939 ;
      RECT MASK 1 118.0865 40.879 118.2065 41.939 ;
      RECT MASK 1 118.5265 40.879 118.6465 41.939 ;
      RECT MASK 1 118.9665 40.879 119.0865 41.939 ;
      RECT MASK 1 119.4065 40.879 119.5265 41.939 ;
      RECT MASK 1 119.8465 40.879 119.9665 41.939 ;
      RECT MASK 1 120.2865 40.879 120.4065 41.939 ;
      RECT MASK 1 120.7265 40.879 120.8465 41.939 ;
      RECT MASK 1 121.1665 40.879 121.2865 41.939 ;
      RECT MASK 1 121.6065 40.879 121.7265 41.939 ;
      RECT MASK 1 122.0465 40.879 122.1665 41.939 ;
      RECT MASK 1 122.4865 40.879 122.6065 41.939 ;
      RECT MASK 1 122.9265 40.879 123.0465 41.939 ;
      RECT MASK 1 123.3665 40.879 123.4865 41.939 ;
      RECT MASK 1 123.8065 40.879 123.9265 41.939 ;
      RECT MASK 1 112.8065 42.199 112.9265 43.289 ;
      RECT MASK 1 113.2465 42.199 113.3665 43.289 ;
      RECT MASK 1 113.6865 42.199 113.8065 43.289 ;
      RECT MASK 1 114.1265 42.199 114.2465 43.289 ;
      RECT MASK 1 114.5665 42.199 114.6865 43.289 ;
      RECT MASK 1 115.0065 42.199 115.1265 43.289 ;
      RECT MASK 1 115.4465 42.199 115.5665 43.289 ;
      RECT MASK 1 115.8865 42.199 116.0065 43.289 ;
      RECT MASK 1 116.3265 42.199 116.4465 43.289 ;
      RECT MASK 1 117.6465 42.199 117.7665 43.289 ;
      RECT MASK 1 118.0865 42.199 118.2065 43.289 ;
      RECT MASK 1 118.5265 42.199 118.6465 43.289 ;
      RECT MASK 1 118.9665 42.199 119.0865 43.289 ;
      RECT MASK 1 119.4065 42.199 119.5265 43.289 ;
      RECT MASK 1 119.8465 42.199 119.9665 43.289 ;
      RECT MASK 1 120.2865 42.199 120.4065 43.289 ;
      RECT MASK 1 120.7265 42.199 120.8465 43.289 ;
      RECT MASK 1 121.1665 42.199 121.2865 43.289 ;
      RECT MASK 1 121.6065 42.199 121.7265 43.289 ;
      RECT MASK 1 122.0465 42.199 122.1665 43.289 ;
      RECT MASK 1 122.4865 42.199 122.6065 43.289 ;
      RECT MASK 1 122.9265 42.199 123.0465 43.289 ;
      RECT MASK 1 123.3665 42.199 123.4865 43.289 ;
      RECT MASK 1 123.8065 42.199 123.9265 43.289 ;
      RECT MASK 1 112.8065 43.549 112.9265 44.639 ;
      RECT MASK 1 113.2465 43.549 113.3665 44.639 ;
      RECT MASK 1 113.6865 43.549 113.8065 44.639 ;
      RECT MASK 1 114.1265 43.549 114.2465 44.639 ;
      RECT MASK 1 114.5665 43.549 114.6865 44.639 ;
      RECT MASK 1 115.0065 43.549 115.1265 44.639 ;
      RECT MASK 1 115.4465 43.549 115.5665 44.639 ;
      RECT MASK 1 115.8865 43.549 116.0065 44.639 ;
      RECT MASK 1 116.3265 43.549 116.4465 44.639 ;
      RECT MASK 1 117.6465 43.549 117.7665 44.639 ;
      RECT MASK 1 118.0865 43.549 118.2065 44.639 ;
      RECT MASK 1 118.5265 43.549 118.6465 44.639 ;
      RECT MASK 1 118.9665 43.549 119.0865 44.639 ;
      RECT MASK 1 119.4065 43.549 119.5265 44.639 ;
      RECT MASK 1 119.8465 43.549 119.9665 44.639 ;
      RECT MASK 1 120.2865 43.549 120.4065 44.639 ;
      RECT MASK 1 120.7265 43.549 120.8465 44.639 ;
      RECT MASK 1 121.1665 43.549 121.2865 44.639 ;
      RECT MASK 1 121.6065 43.549 121.7265 44.639 ;
      RECT MASK 1 122.0465 43.549 122.1665 44.639 ;
      RECT MASK 1 122.4865 43.549 122.6065 44.639 ;
      RECT MASK 1 122.9265 43.549 123.0465 44.639 ;
      RECT MASK 1 123.3665 43.549 123.4865 44.639 ;
      RECT MASK 1 123.8065 43.549 123.9265 44.639 ;
      RECT MASK 1 112.8065 44.899 112.9265 46.709 ;
      RECT MASK 1 113.2465 44.899 113.3665 46.709 ;
      RECT MASK 1 113.6865 44.899 113.8065 46.709 ;
      RECT MASK 1 114.1265 44.899 114.2465 46.709 ;
      RECT MASK 1 114.5665 44.899 114.6865 46.709 ;
      RECT MASK 1 115.0065 44.899 115.1265 46.709 ;
      RECT MASK 1 115.4465 44.899 115.5665 46.709 ;
      RECT MASK 1 115.8865 44.899 116.0065 46.709 ;
      RECT MASK 1 116.3265 44.899 116.4465 46.709 ;
      RECT MASK 1 117.6465 44.899 117.7665 46.709 ;
      RECT MASK 1 118.0865 44.899 118.2065 46.709 ;
      RECT MASK 1 118.5265 44.899 118.6465 46.709 ;
      RECT MASK 1 118.9665 44.899 119.0865 46.709 ;
      RECT MASK 1 119.4065 44.899 119.5265 46.709 ;
      RECT MASK 1 119.8465 44.899 119.9665 46.709 ;
      RECT MASK 1 120.2865 44.899 120.4065 46.709 ;
      RECT MASK 1 120.7265 44.899 120.8465 46.709 ;
      RECT MASK 1 121.1665 44.899 121.2865 46.709 ;
      RECT MASK 1 121.6065 44.899 121.7265 46.709 ;
      RECT MASK 1 122.0465 44.899 122.1665 46.709 ;
      RECT MASK 1 122.4865 44.899 122.6065 46.709 ;
      RECT MASK 1 122.9265 44.899 123.0465 46.709 ;
      RECT MASK 1 123.3665 44.899 123.4865 46.709 ;
      RECT MASK 1 123.8065 44.899 123.9265 46.709 ;
      RECT MASK 1 112.8065 46.969 112.9265 48.119 ;
      RECT MASK 1 113.2465 46.969 113.3665 48.119 ;
      RECT MASK 1 113.6865 46.969 113.8065 48.119 ;
      RECT MASK 1 114.1265 46.969 114.2465 48.119 ;
      RECT MASK 1 114.5665 46.969 114.6865 48.119 ;
      RECT MASK 1 115.0065 46.969 115.1265 48.119 ;
      RECT MASK 1 115.4465 46.969 115.5665 48.119 ;
      RECT MASK 1 115.8865 46.969 116.0065 48.119 ;
      RECT MASK 1 116.3265 46.969 116.4465 48.119 ;
      RECT MASK 1 117.6465 46.969 117.7665 48.059 ;
      RECT MASK 1 118.0865 46.969 118.2065 48.059 ;
      RECT MASK 1 118.5265 46.969 118.6465 48.059 ;
      RECT MASK 1 118.9665 46.969 119.0865 48.059 ;
      RECT MASK 1 119.4065 46.969 119.5265 48.059 ;
      RECT MASK 1 119.8465 46.969 119.9665 48.059 ;
      RECT MASK 1 120.2865 46.969 120.4065 48.059 ;
      RECT MASK 1 120.7265 46.969 120.8465 48.059 ;
      RECT MASK 1 121.1665 46.969 121.2865 48.059 ;
      RECT MASK 1 121.6065 46.969 121.7265 48.059 ;
      RECT MASK 1 122.0465 46.969 122.1665 48.059 ;
      RECT MASK 1 122.4865 46.969 122.6065 48.059 ;
      RECT MASK 1 122.9265 46.969 123.0465 48.059 ;
      RECT MASK 1 123.3665 46.969 123.4865 48.059 ;
      RECT MASK 1 123.8065 46.969 123.9265 48.059 ;
      RECT MASK 1 112.8065 48.379 112.9265 49.409 ;
      RECT MASK 1 113.2465 48.379 113.3665 49.409 ;
      RECT MASK 1 113.6865 48.379 113.8065 49.409 ;
      RECT MASK 1 114.1265 48.379 114.2465 49.409 ;
      RECT MASK 1 114.5665 48.379 114.6865 49.409 ;
      RECT MASK 1 115.0065 48.379 115.1265 49.409 ;
      RECT MASK 1 115.4465 48.379 115.5665 49.409 ;
      RECT MASK 1 115.8865 48.379 116.0065 49.409 ;
      RECT MASK 1 116.3265 48.379 116.4465 49.409 ;
      RECT MASK 1 112.8065 49.669 112.9265 50.759 ;
      RECT MASK 1 113.2465 49.669 113.3665 50.759 ;
      RECT MASK 1 113.6865 49.669 113.8065 50.759 ;
      RECT MASK 1 114.1265 49.669 114.2465 50.759 ;
      RECT MASK 1 114.5665 49.669 114.6865 50.759 ;
      RECT MASK 1 115.0065 49.669 115.1265 50.759 ;
      RECT MASK 1 115.4465 49.669 115.5665 50.759 ;
      RECT MASK 1 115.8865 49.669 116.0065 50.759 ;
      RECT MASK 1 116.3265 49.669 116.4465 50.759 ;
      RECT MASK 1 4.711 51.6 4.771 51.84 ;
      RECT MASK 1 5.151 51.6 5.211 51.84 ;
      RECT MASK 1 5.591 51.6 5.651 51.84 ;
      RECT MASK 1 6.031 51.6 6.091 51.84 ;
      RECT MASK 1 6.471 51.6 6.531 51.84 ;
      RECT MASK 1 6.911 51.6 6.971 51.84 ;
      RECT MASK 1 7.351 51.6 7.411 51.84 ;
      RECT MASK 1 7.791 51.6 7.851 51.84 ;
      RECT MASK 1 8.231 51.6 8.291 51.84 ;
      RECT MASK 1 8.671 51.6 8.731 51.84 ;
      RECT MASK 1 9.111 51.6 9.171 51.84 ;
      RECT MASK 1 9.551 51.6 9.611 51.84 ;
      RECT MASK 1 9.991 51.6 10.051 51.84 ;
      RECT MASK 1 10.431 51.6 10.491 51.84 ;
      RECT MASK 1 10.871 51.6 10.931 51.84 ;
      RECT MASK 1 11.329 51.6 11.389 51.84 ;
      RECT MASK 1 11.769 51.6 11.829 51.84 ;
      RECT MASK 1 12.209 51.6 12.269 51.84 ;
      RECT MASK 1 12.649 51.6 12.709 51.84 ;
      RECT MASK 1 13.089 51.6 13.149 51.84 ;
      RECT MASK 1 13.529 51.6 13.589 51.84 ;
      RECT MASK 1 13.969 51.6 14.029 51.84 ;
      RECT MASK 1 14.409 51.6 14.469 51.84 ;
      RECT MASK 1 14.849 51.6 14.909 51.84 ;
      RECT MASK 1 15.289 51.6 15.349 51.84 ;
      RECT MASK 1 15.729 51.6 15.789 51.84 ;
      RECT MASK 1 16.169 51.6 16.229 51.84 ;
      RECT MASK 1 16.609 51.6 16.669 51.84 ;
      RECT MASK 1 17.049 51.6 17.109 51.84 ;
      RECT MASK 1 17.489 51.6 17.549 51.84 ;
      RECT MASK 1 17.947 51.6 18.007 51.84 ;
      RECT MASK 1 18.387 51.6 18.447 51.84 ;
      RECT MASK 1 18.827 51.6 18.887 51.84 ;
      RECT MASK 1 19.267 51.6 19.327 51.84 ;
      RECT MASK 1 19.707 51.6 19.767 51.84 ;
      RECT MASK 1 20.147 51.6 20.207 51.84 ;
      RECT MASK 1 20.587 51.6 20.647 51.84 ;
      RECT MASK 1 21.027 51.6 21.087 51.84 ;
      RECT MASK 1 21.467 51.6 21.527 51.84 ;
      RECT MASK 1 21.907 51.6 21.967 51.84 ;
      RECT MASK 1 22.347 51.6 22.407 51.84 ;
      RECT MASK 1 22.787 51.6 22.847 51.84 ;
      RECT MASK 1 23.227 51.6 23.287 51.84 ;
      RECT MASK 1 23.667 51.6 23.727 51.84 ;
      RECT MASK 1 24.107 51.6 24.167 51.84 ;
      RECT MASK 1 24.565 51.6 24.625 51.84 ;
      RECT MASK 1 25.005 51.6 25.065 51.84 ;
      RECT MASK 1 25.445 51.6 25.505 51.84 ;
      RECT MASK 1 25.885 51.6 25.945 51.84 ;
      RECT MASK 1 26.325 51.6 26.385 51.84 ;
      RECT MASK 1 26.765 51.6 26.825 51.84 ;
      RECT MASK 1 27.205 51.6 27.265 51.84 ;
      RECT MASK 1 27.645 51.6 27.705 51.84 ;
      RECT MASK 1 28.085 51.6 28.145 51.84 ;
      RECT MASK 1 28.525 51.6 28.585 51.84 ;
      RECT MASK 1 28.965 51.6 29.025 51.84 ;
      RECT MASK 1 29.405 51.6 29.465 51.84 ;
      RECT MASK 1 29.845 51.6 29.905 51.84 ;
      RECT MASK 1 30.285 51.6 30.345 51.84 ;
      RECT MASK 1 30.725 51.6 30.785 51.84 ;
      RECT MASK 1 31.183 51.6 31.243 51.84 ;
      RECT MASK 1 31.623 51.6 31.683 51.84 ;
      RECT MASK 1 32.063 51.6 32.123 51.84 ;
      RECT MASK 1 32.503 51.6 32.563 51.84 ;
      RECT MASK 1 32.943 51.6 33.003 51.84 ;
      RECT MASK 1 33.383 51.6 33.443 51.84 ;
      RECT MASK 1 33.823 51.6 33.883 51.84 ;
      RECT MASK 1 34.263 51.6 34.323 51.84 ;
      RECT MASK 1 34.703 51.6 34.763 51.84 ;
      RECT MASK 1 35.143 51.6 35.203 51.84 ;
      RECT MASK 1 35.583 51.6 35.643 51.84 ;
      RECT MASK 1 36.023 51.6 36.083 51.84 ;
      RECT MASK 1 36.463 51.6 36.523 51.84 ;
      RECT MASK 1 36.903 51.6 36.963 51.84 ;
      RECT MASK 1 37.343 51.6 37.403 51.84 ;
      RECT MASK 1 37.801 51.6 37.861 51.84 ;
      RECT MASK 1 38.241 51.6 38.301 51.84 ;
      RECT MASK 1 38.681 51.6 38.741 51.84 ;
      RECT MASK 1 39.121 51.6 39.181 51.84 ;
      RECT MASK 1 39.561 51.6 39.621 51.84 ;
      RECT MASK 1 40.001 51.6 40.061 51.84 ;
      RECT MASK 1 40.441 51.6 40.501 51.84 ;
      RECT MASK 1 40.881 51.6 40.941 51.84 ;
      RECT MASK 1 41.321 51.6 41.381 51.84 ;
      RECT MASK 1 41.761 51.6 41.821 51.84 ;
      RECT MASK 1 43.081 51.6 43.141 51.84 ;
      RECT MASK 1 43.521 51.6 43.581 51.84 ;
      RECT MASK 1 43.961 51.6 44.021 51.84 ;
      RECT MASK 1 44.419 51.6 44.479 51.84 ;
      RECT MASK 1 44.859 51.6 44.919 51.84 ;
      RECT MASK 1 45.299 51.6 45.359 51.84 ;
      RECT MASK 1 45.739 51.6 45.799 51.84 ;
      RECT MASK 1 46.179 51.6 46.239 51.84 ;
      RECT MASK 1 46.619 51.6 46.679 51.84 ;
      RECT MASK 1 47.059 51.6 47.119 51.84 ;
      RECT MASK 1 47.499 51.6 47.559 51.84 ;
      RECT MASK 1 47.939 51.6 47.999 51.84 ;
      RECT MASK 1 48.379 51.6 48.439 51.84 ;
      RECT MASK 1 48.819 51.6 48.879 51.84 ;
      RECT MASK 1 49.259 51.6 49.319 51.84 ;
      RECT MASK 1 49.699 51.6 49.759 51.84 ;
      RECT MASK 1 50.139 51.6 50.199 51.84 ;
      RECT MASK 1 50.579 51.6 50.639 51.84 ;
      RECT MASK 1 51.037 51.6 51.097 51.84 ;
      RECT MASK 1 51.477 51.6 51.537 51.84 ;
      RECT MASK 1 51.917 51.6 51.977 51.84 ;
      RECT MASK 1 52.357 51.6 52.417 51.84 ;
      RECT MASK 1 52.797 51.6 52.857 51.84 ;
      RECT MASK 1 53.237 51.6 53.297 51.84 ;
      RECT MASK 1 53.677 51.6 53.737 51.84 ;
      RECT MASK 1 54.117 51.6 54.177 51.84 ;
      RECT MASK 1 54.557 51.6 54.617 51.84 ;
      RECT MASK 1 54.997 51.6 55.057 51.84 ;
      RECT MASK 1 55.437 51.6 55.497 51.84 ;
      RECT MASK 1 55.877 51.6 55.937 51.84 ;
      RECT MASK 1 56.317 51.6 56.377 51.84 ;
      RECT MASK 1 56.757 51.6 56.817 51.84 ;
      RECT MASK 1 57.197 51.6 57.257 51.84 ;
      RECT MASK 1 57.655 51.6 57.715 51.84 ;
      RECT MASK 1 58.095 51.6 58.155 51.84 ;
      RECT MASK 1 58.535 51.6 58.595 51.84 ;
      RECT MASK 1 58.975 51.6 59.035 51.84 ;
      RECT MASK 1 59.415 51.6 59.475 51.84 ;
      RECT MASK 1 59.855 51.6 59.915 51.84 ;
      RECT MASK 1 60.295 51.6 60.355 51.84 ;
      RECT MASK 1 60.735 51.6 60.795 51.84 ;
      RECT MASK 1 61.175 51.6 61.235 51.84 ;
      RECT MASK 1 61.615 51.6 61.675 51.84 ;
      RECT MASK 1 62.055 51.6 62.115 51.84 ;
      RECT MASK 1 62.495 51.6 62.555 51.84 ;
      RECT MASK 1 62.935 51.6 62.995 51.84 ;
      RECT MASK 1 63.375 51.6 63.435 51.84 ;
      RECT MASK 1 63.815 51.6 63.875 51.84 ;
      RECT MASK 1 64.273 51.6 64.333 51.84 ;
      RECT MASK 1 64.713 51.6 64.773 51.84 ;
      RECT MASK 1 65.153 51.6 65.213 51.84 ;
      RECT MASK 1 65.593 51.6 65.653 51.84 ;
      RECT MASK 1 66.033 51.6 66.093 51.84 ;
      RECT MASK 1 66.473 51.6 66.533 51.84 ;
      RECT MASK 1 66.913 51.6 66.973 51.84 ;
      RECT MASK 1 67.353 51.6 67.413 51.84 ;
      RECT MASK 1 67.793 51.6 67.853 51.84 ;
      RECT MASK 1 68.233 51.6 68.293 51.84 ;
      RECT MASK 1 68.673 51.6 68.733 51.84 ;
      RECT MASK 1 69.113 51.6 69.173 51.84 ;
      RECT MASK 1 69.553 51.6 69.613 51.84 ;
      RECT MASK 1 69.993 51.6 70.053 51.84 ;
      RECT MASK 1 70.433 51.6 70.493 51.84 ;
      RECT MASK 1 70.891 51.6 70.951 51.84 ;
      RECT MASK 1 71.331 51.6 71.391 51.84 ;
      RECT MASK 1 71.771 51.6 71.831 51.84 ;
      RECT MASK 1 72.211 51.6 72.271 51.84 ;
      RECT MASK 1 72.651 51.6 72.711 51.84 ;
      RECT MASK 1 73.091 51.6 73.151 51.84 ;
      RECT MASK 1 73.531 51.6 73.591 51.84 ;
      RECT MASK 1 73.971 51.6 74.031 51.84 ;
      RECT MASK 1 74.411 51.6 74.471 51.84 ;
      RECT MASK 1 74.851 51.6 74.911 51.84 ;
      RECT MASK 1 75.291 51.6 75.351 51.84 ;
      RECT MASK 1 75.731 51.6 75.791 51.84 ;
      RECT MASK 1 76.171 51.6 76.231 51.84 ;
      RECT MASK 1 76.611 51.6 76.671 51.84 ;
      RECT MASK 1 77.051 51.6 77.111 51.84 ;
      RECT MASK 1 77.509 51.6 77.569 51.84 ;
      RECT MASK 1 77.949 51.6 78.009 51.84 ;
      RECT MASK 1 78.389 51.6 78.449 51.84 ;
      RECT MASK 1 78.829 51.6 78.889 51.84 ;
      RECT MASK 1 79.269 51.6 79.329 51.84 ;
      RECT MASK 1 79.709 51.6 79.769 51.84 ;
      RECT MASK 1 80.149 51.6 80.209 51.84 ;
      RECT MASK 1 80.589 51.6 80.649 51.84 ;
      RECT MASK 1 81.029 51.6 81.089 51.84 ;
      RECT MASK 1 81.469 51.6 81.529 51.84 ;
      RECT MASK 1 81.909 51.6 81.969 51.84 ;
      RECT MASK 1 82.349 51.6 82.409 51.84 ;
      RECT MASK 1 83.669 51.6 83.729 51.84 ;
      RECT MASK 1 84.127 51.6 84.187 51.84 ;
      RECT MASK 1 84.567 51.6 84.627 51.84 ;
      RECT MASK 1 85.007 51.6 85.067 51.84 ;
      RECT MASK 1 85.447 51.6 85.507 51.84 ;
      RECT MASK 1 85.887 51.6 85.947 51.84 ;
      RECT MASK 1 86.327 51.6 86.387 51.84 ;
      RECT MASK 1 86.767 51.6 86.827 51.84 ;
      RECT MASK 1 87.207 51.6 87.267 51.84 ;
      RECT MASK 1 87.647 51.6 87.707 51.84 ;
      RECT MASK 1 88.087 51.6 88.147 51.84 ;
      RECT MASK 1 88.527 51.6 88.587 51.84 ;
      RECT MASK 1 88.967 51.6 89.027 51.84 ;
      RECT MASK 1 89.407 51.6 89.467 51.84 ;
      RECT MASK 1 89.847 51.6 89.907 51.84 ;
      RECT MASK 1 90.287 51.6 90.347 51.84 ;
      RECT MASK 1 90.745 51.6 90.805 51.84 ;
      RECT MASK 1 91.185 51.6 91.245 51.84 ;
      RECT MASK 1 91.625 51.6 91.685 51.84 ;
      RECT MASK 1 92.065 51.6 92.125 51.84 ;
      RECT MASK 1 92.505 51.6 92.565 51.84 ;
      RECT MASK 1 92.945 51.6 93.005 51.84 ;
      RECT MASK 1 93.385 51.6 93.445 51.84 ;
      RECT MASK 1 93.825 51.6 93.885 51.84 ;
      RECT MASK 1 94.265 51.6 94.325 51.84 ;
      RECT MASK 1 94.705 51.6 94.765 51.84 ;
      RECT MASK 1 95.145 51.6 95.205 51.84 ;
      RECT MASK 1 95.585 51.6 95.645 51.84 ;
      RECT MASK 1 96.025 51.6 96.085 51.84 ;
      RECT MASK 1 96.465 51.6 96.525 51.84 ;
      RECT MASK 1 96.905 51.6 96.965 51.84 ;
      RECT MASK 1 97.363 51.6 97.423 51.84 ;
      RECT MASK 1 97.803 51.6 97.863 51.84 ;
      RECT MASK 1 98.243 51.6 98.303 51.84 ;
      RECT MASK 1 98.683 51.6 98.743 51.84 ;
      RECT MASK 1 99.123 51.6 99.183 51.84 ;
      RECT MASK 1 99.563 51.6 99.623 51.84 ;
      RECT MASK 1 100.003 51.6 100.063 51.84 ;
      RECT MASK 1 100.443 51.6 100.503 51.84 ;
      RECT MASK 1 100.883 51.6 100.943 51.84 ;
      RECT MASK 1 101.323 51.6 101.383 51.84 ;
      RECT MASK 1 101.763 51.6 101.823 51.84 ;
      RECT MASK 1 102.203 51.6 102.263 51.84 ;
      RECT MASK 1 102.643 51.6 102.703 51.84 ;
      RECT MASK 1 103.083 51.6 103.143 51.84 ;
      RECT MASK 1 103.523 51.6 103.583 51.84 ;
      RECT MASK 1 103.981 51.6 104.041 51.84 ;
      RECT MASK 1 104.421 51.6 104.481 51.84 ;
      RECT MASK 1 104.861 51.6 104.921 51.84 ;
      RECT MASK 1 105.301 51.6 105.361 51.84 ;
      RECT MASK 1 105.741 51.6 105.801 51.84 ;
      RECT MASK 1 106.181 51.6 106.241 51.84 ;
      RECT MASK 1 106.621 51.6 106.681 51.84 ;
      RECT MASK 1 107.061 51.6 107.121 51.84 ;
      RECT MASK 1 107.501 51.6 107.561 51.84 ;
      RECT MASK 1 107.941 51.6 108.001 51.84 ;
      RECT MASK 1 108.381 51.6 108.441 51.84 ;
      RECT MASK 1 108.821 51.6 108.881 51.84 ;
      RECT MASK 1 109.261 51.6 109.321 51.84 ;
      RECT MASK 1 109.701 51.6 109.761 51.84 ;
      RECT MASK 1 110.141 51.6 110.201 51.84 ;
      RECT MASK 1 4.711 52.02 4.771 52.26 ;
      RECT MASK 1 5.151 52.02 5.211 52.26 ;
      RECT MASK 1 5.591 52.02 5.651 52.26 ;
      RECT MASK 1 6.031 52.02 6.091 52.26 ;
      RECT MASK 1 6.471 52.02 6.531 52.26 ;
      RECT MASK 1 6.911 52.02 6.971 52.26 ;
      RECT MASK 1 7.351 52.02 7.411 52.26 ;
      RECT MASK 1 7.791 52.02 7.851 52.26 ;
      RECT MASK 1 8.231 52.02 8.291 52.26 ;
      RECT MASK 1 8.671 52.02 8.731 52.26 ;
      RECT MASK 1 9.111 52.02 9.171 52.26 ;
      RECT MASK 1 9.551 52.02 9.611 52.26 ;
      RECT MASK 1 9.991 52.02 10.051 52.26 ;
      RECT MASK 1 10.431 52.02 10.491 52.26 ;
      RECT MASK 1 10.871 52.02 10.931 52.26 ;
      RECT MASK 1 11.329 52.02 11.389 52.26 ;
      RECT MASK 1 11.769 52.02 11.829 52.26 ;
      RECT MASK 1 12.209 52.02 12.269 52.26 ;
      RECT MASK 1 12.649 52.02 12.709 52.26 ;
      RECT MASK 1 13.089 52.02 13.149 52.26 ;
      RECT MASK 1 13.529 52.02 13.589 52.26 ;
      RECT MASK 1 13.969 52.02 14.029 52.26 ;
      RECT MASK 1 14.409 52.02 14.469 52.26 ;
      RECT MASK 1 14.849 52.02 14.909 52.26 ;
      RECT MASK 1 15.289 52.02 15.349 52.26 ;
      RECT MASK 1 15.729 52.02 15.789 52.26 ;
      RECT MASK 1 16.169 52.02 16.229 52.26 ;
      RECT MASK 1 16.609 52.02 16.669 52.26 ;
      RECT MASK 1 17.049 52.02 17.109 52.26 ;
      RECT MASK 1 17.489 52.02 17.549 52.26 ;
      RECT MASK 1 17.947 52.02 18.007 52.26 ;
      RECT MASK 1 18.387 52.02 18.447 52.26 ;
      RECT MASK 1 18.827 52.02 18.887 52.26 ;
      RECT MASK 1 19.267 52.02 19.327 52.26 ;
      RECT MASK 1 19.707 52.02 19.767 52.26 ;
      RECT MASK 1 20.147 52.02 20.207 52.26 ;
      RECT MASK 1 20.587 52.02 20.647 52.26 ;
      RECT MASK 1 21.027 52.02 21.087 52.26 ;
      RECT MASK 1 21.467 52.02 21.527 52.26 ;
      RECT MASK 1 21.907 52.02 21.967 52.26 ;
      RECT MASK 1 22.347 52.02 22.407 52.26 ;
      RECT MASK 1 22.787 52.02 22.847 52.26 ;
      RECT MASK 1 23.227 52.02 23.287 52.26 ;
      RECT MASK 1 23.667 52.02 23.727 52.26 ;
      RECT MASK 1 24.107 52.02 24.167 52.26 ;
      RECT MASK 1 24.565 52.02 24.625 52.26 ;
      RECT MASK 1 25.005 52.02 25.065 52.26 ;
      RECT MASK 1 25.445 52.02 25.505 52.26 ;
      RECT MASK 1 25.885 52.02 25.945 52.26 ;
      RECT MASK 1 26.325 52.02 26.385 52.26 ;
      RECT MASK 1 26.765 52.02 26.825 52.26 ;
      RECT MASK 1 27.205 52.02 27.265 52.26 ;
      RECT MASK 1 27.645 52.02 27.705 52.26 ;
      RECT MASK 1 28.085 52.02 28.145 52.26 ;
      RECT MASK 1 28.525 52.02 28.585 52.26 ;
      RECT MASK 1 28.965 52.02 29.025 52.26 ;
      RECT MASK 1 29.405 52.02 29.465 52.26 ;
      RECT MASK 1 29.845 52.02 29.905 52.26 ;
      RECT MASK 1 30.285 52.02 30.345 52.26 ;
      RECT MASK 1 30.725 52.02 30.785 52.26 ;
      RECT MASK 1 31.183 52.02 31.243 52.26 ;
      RECT MASK 1 31.623 52.02 31.683 52.26 ;
      RECT MASK 1 32.063 52.02 32.123 52.26 ;
      RECT MASK 1 32.503 52.02 32.563 52.26 ;
      RECT MASK 1 32.943 52.02 33.003 52.26 ;
      RECT MASK 1 33.383 52.02 33.443 52.26 ;
      RECT MASK 1 33.823 52.02 33.883 52.26 ;
      RECT MASK 1 34.263 52.02 34.323 52.26 ;
      RECT MASK 1 34.703 52.02 34.763 52.26 ;
      RECT MASK 1 35.143 52.02 35.203 52.26 ;
      RECT MASK 1 35.583 52.02 35.643 52.26 ;
      RECT MASK 1 36.023 52.02 36.083 52.26 ;
      RECT MASK 1 36.463 52.02 36.523 52.26 ;
      RECT MASK 1 36.903 52.02 36.963 52.26 ;
      RECT MASK 1 37.343 52.02 37.403 52.26 ;
      RECT MASK 1 37.801 52.02 37.861 52.26 ;
      RECT MASK 1 38.241 52.02 38.301 52.26 ;
      RECT MASK 1 38.681 52.02 38.741 52.26 ;
      RECT MASK 1 39.121 52.02 39.181 52.26 ;
      RECT MASK 1 39.561 52.02 39.621 52.26 ;
      RECT MASK 1 40.001 52.02 40.061 52.26 ;
      RECT MASK 1 40.441 52.02 40.501 52.26 ;
      RECT MASK 1 40.881 52.02 40.941 52.26 ;
      RECT MASK 1 41.321 52.02 41.381 52.26 ;
      RECT MASK 1 41.761 52.02 41.821 52.26 ;
      RECT MASK 1 43.081 52.02 43.141 52.26 ;
      RECT MASK 1 43.521 52.02 43.581 52.26 ;
      RECT MASK 1 43.961 52.02 44.021 52.26 ;
      RECT MASK 1 44.419 52.02 44.479 52.26 ;
      RECT MASK 1 44.859 52.02 44.919 52.26 ;
      RECT MASK 1 45.299 52.02 45.359 52.26 ;
      RECT MASK 1 45.739 52.02 45.799 52.26 ;
      RECT MASK 1 46.179 52.02 46.239 52.26 ;
      RECT MASK 1 46.619 52.02 46.679 52.26 ;
      RECT MASK 1 47.059 52.02 47.119 52.26 ;
      RECT MASK 1 47.499 52.02 47.559 52.26 ;
      RECT MASK 1 47.939 52.02 47.999 52.26 ;
      RECT MASK 1 48.379 52.02 48.439 52.26 ;
      RECT MASK 1 48.819 52.02 48.879 52.26 ;
      RECT MASK 1 49.259 52.02 49.319 52.26 ;
      RECT MASK 1 49.699 52.02 49.759 52.26 ;
      RECT MASK 1 50.139 52.02 50.199 52.26 ;
      RECT MASK 1 50.579 52.02 50.639 52.26 ;
      RECT MASK 1 51.037 52.02 51.097 52.26 ;
      RECT MASK 1 51.477 52.02 51.537 52.26 ;
      RECT MASK 1 51.917 52.02 51.977 52.26 ;
      RECT MASK 1 52.357 52.02 52.417 52.26 ;
      RECT MASK 1 52.797 52.02 52.857 52.26 ;
      RECT MASK 1 53.237 52.02 53.297 52.26 ;
      RECT MASK 1 53.677 52.02 53.737 52.26 ;
      RECT MASK 1 54.117 52.02 54.177 52.26 ;
      RECT MASK 1 54.557 52.02 54.617 52.26 ;
      RECT MASK 1 54.997 52.02 55.057 52.26 ;
      RECT MASK 1 55.437 52.02 55.497 52.26 ;
      RECT MASK 1 55.877 52.02 55.937 52.26 ;
      RECT MASK 1 56.317 52.02 56.377 52.26 ;
      RECT MASK 1 56.757 52.02 56.817 52.26 ;
      RECT MASK 1 57.197 52.02 57.257 52.26 ;
      RECT MASK 1 57.655 52.02 57.715 52.26 ;
      RECT MASK 1 58.095 52.02 58.155 52.26 ;
      RECT MASK 1 58.535 52.02 58.595 52.26 ;
      RECT MASK 1 58.975 52.02 59.035 52.26 ;
      RECT MASK 1 59.415 52.02 59.475 52.26 ;
      RECT MASK 1 59.855 52.02 59.915 52.26 ;
      RECT MASK 1 60.295 52.02 60.355 52.26 ;
      RECT MASK 1 60.735 52.02 60.795 52.26 ;
      RECT MASK 1 61.175 52.02 61.235 52.26 ;
      RECT MASK 1 61.615 52.02 61.675 52.26 ;
      RECT MASK 1 62.055 52.02 62.115 52.26 ;
      RECT MASK 1 62.495 52.02 62.555 52.26 ;
      RECT MASK 1 62.935 52.02 62.995 52.26 ;
      RECT MASK 1 63.375 52.02 63.435 52.26 ;
      RECT MASK 1 63.815 52.02 63.875 52.26 ;
      RECT MASK 1 64.273 52.02 64.333 52.26 ;
      RECT MASK 1 64.713 52.02 64.773 52.26 ;
      RECT MASK 1 65.153 52.02 65.213 52.26 ;
      RECT MASK 1 65.593 52.02 65.653 52.26 ;
      RECT MASK 1 66.033 52.02 66.093 52.26 ;
      RECT MASK 1 66.473 52.02 66.533 52.26 ;
      RECT MASK 1 66.913 52.02 66.973 52.26 ;
      RECT MASK 1 67.353 52.02 67.413 52.26 ;
      RECT MASK 1 67.793 52.02 67.853 52.26 ;
      RECT MASK 1 68.233 52.02 68.293 52.26 ;
      RECT MASK 1 68.673 52.02 68.733 52.26 ;
      RECT MASK 1 69.113 52.02 69.173 52.26 ;
      RECT MASK 1 69.553 52.02 69.613 52.26 ;
      RECT MASK 1 69.993 52.02 70.053 52.26 ;
      RECT MASK 1 70.433 52.02 70.493 52.26 ;
      RECT MASK 1 70.891 52.02 70.951 52.26 ;
      RECT MASK 1 71.331 52.02 71.391 52.26 ;
      RECT MASK 1 71.771 52.02 71.831 52.26 ;
      RECT MASK 1 72.211 52.02 72.271 52.26 ;
      RECT MASK 1 72.651 52.02 72.711 52.26 ;
      RECT MASK 1 73.091 52.02 73.151 52.26 ;
      RECT MASK 1 73.531 52.02 73.591 52.26 ;
      RECT MASK 1 73.971 52.02 74.031 52.26 ;
      RECT MASK 1 74.411 52.02 74.471 52.26 ;
      RECT MASK 1 74.851 52.02 74.911 52.26 ;
      RECT MASK 1 75.291 52.02 75.351 52.26 ;
      RECT MASK 1 75.731 52.02 75.791 52.26 ;
      RECT MASK 1 76.171 52.02 76.231 52.26 ;
      RECT MASK 1 76.611 52.02 76.671 52.26 ;
      RECT MASK 1 77.051 52.02 77.111 52.26 ;
      RECT MASK 1 77.509 52.02 77.569 52.26 ;
      RECT MASK 1 77.949 52.02 78.009 52.26 ;
      RECT MASK 1 78.389 52.02 78.449 52.26 ;
      RECT MASK 1 78.829 52.02 78.889 52.26 ;
      RECT MASK 1 79.269 52.02 79.329 52.26 ;
      RECT MASK 1 79.709 52.02 79.769 52.26 ;
      RECT MASK 1 80.149 52.02 80.209 52.26 ;
      RECT MASK 1 80.589 52.02 80.649 52.26 ;
      RECT MASK 1 81.029 52.02 81.089 52.26 ;
      RECT MASK 1 81.469 52.02 81.529 52.26 ;
      RECT MASK 1 81.909 52.02 81.969 52.26 ;
      RECT MASK 1 82.349 52.02 82.409 52.26 ;
      RECT MASK 1 83.669 52.02 83.729 52.26 ;
      RECT MASK 1 84.127 52.02 84.187 52.26 ;
      RECT MASK 1 84.567 52.02 84.627 52.26 ;
      RECT MASK 1 85.007 52.02 85.067 52.26 ;
      RECT MASK 1 85.447 52.02 85.507 52.26 ;
      RECT MASK 1 85.887 52.02 85.947 52.26 ;
      RECT MASK 1 86.327 52.02 86.387 52.26 ;
      RECT MASK 1 86.767 52.02 86.827 52.26 ;
      RECT MASK 1 87.207 52.02 87.267 52.26 ;
      RECT MASK 1 87.647 52.02 87.707 52.26 ;
      RECT MASK 1 88.087 52.02 88.147 52.26 ;
      RECT MASK 1 88.527 52.02 88.587 52.26 ;
      RECT MASK 1 88.967 52.02 89.027 52.26 ;
      RECT MASK 1 89.407 52.02 89.467 52.26 ;
      RECT MASK 1 89.847 52.02 89.907 52.26 ;
      RECT MASK 1 90.287 52.02 90.347 52.26 ;
      RECT MASK 1 90.745 52.02 90.805 52.26 ;
      RECT MASK 1 91.185 52.02 91.245 52.26 ;
      RECT MASK 1 91.625 52.02 91.685 52.26 ;
      RECT MASK 1 92.065 52.02 92.125 52.26 ;
      RECT MASK 1 92.505 52.02 92.565 52.26 ;
      RECT MASK 1 92.945 52.02 93.005 52.26 ;
      RECT MASK 1 93.385 52.02 93.445 52.26 ;
      RECT MASK 1 93.825 52.02 93.885 52.26 ;
      RECT MASK 1 94.265 52.02 94.325 52.26 ;
      RECT MASK 1 94.705 52.02 94.765 52.26 ;
      RECT MASK 1 95.145 52.02 95.205 52.26 ;
      RECT MASK 1 95.585 52.02 95.645 52.26 ;
      RECT MASK 1 96.025 52.02 96.085 52.26 ;
      RECT MASK 1 96.465 52.02 96.525 52.26 ;
      RECT MASK 1 96.905 52.02 96.965 52.26 ;
      RECT MASK 1 97.363 52.02 97.423 52.26 ;
      RECT MASK 1 97.803 52.02 97.863 52.26 ;
      RECT MASK 1 98.243 52.02 98.303 52.26 ;
      RECT MASK 1 98.683 52.02 98.743 52.26 ;
      RECT MASK 1 99.123 52.02 99.183 52.26 ;
      RECT MASK 1 99.563 52.02 99.623 52.26 ;
      RECT MASK 1 100.003 52.02 100.063 52.26 ;
      RECT MASK 1 100.443 52.02 100.503 52.26 ;
      RECT MASK 1 100.883 52.02 100.943 52.26 ;
      RECT MASK 1 101.323 52.02 101.383 52.26 ;
      RECT MASK 1 101.763 52.02 101.823 52.26 ;
      RECT MASK 1 102.203 52.02 102.263 52.26 ;
      RECT MASK 1 102.643 52.02 102.703 52.26 ;
      RECT MASK 1 103.083 52.02 103.143 52.26 ;
      RECT MASK 1 103.523 52.02 103.583 52.26 ;
      RECT MASK 1 103.981 52.02 104.041 52.26 ;
      RECT MASK 1 104.421 52.02 104.481 52.26 ;
      RECT MASK 1 104.861 52.02 104.921 52.26 ;
      RECT MASK 1 105.301 52.02 105.361 52.26 ;
      RECT MASK 1 105.741 52.02 105.801 52.26 ;
      RECT MASK 1 106.181 52.02 106.241 52.26 ;
      RECT MASK 1 106.621 52.02 106.681 52.26 ;
      RECT MASK 1 107.061 52.02 107.121 52.26 ;
      RECT MASK 1 107.501 52.02 107.561 52.26 ;
      RECT MASK 1 107.941 52.02 108.001 52.26 ;
      RECT MASK 1 108.381 52.02 108.441 52.26 ;
      RECT MASK 1 108.821 52.02 108.881 52.26 ;
      RECT MASK 1 109.261 52.02 109.321 52.26 ;
      RECT MASK 1 109.701 52.02 109.761 52.26 ;
      RECT MASK 1 110.141 52.02 110.201 52.26 ;
      RECT MASK 1 4.681 52.459 4.801 63.671 ;
      RECT MASK 1 5.121 52.459 5.241 63.671 ;
      RECT MASK 1 5.561 52.459 5.681 63.671 ;
      RECT MASK 1 6.001 52.459 6.121 63.671 ;
      RECT MASK 1 6.441 52.459 6.561 63.671 ;
      RECT MASK 1 6.881 52.459 7.001 63.671 ;
      RECT MASK 1 7.321 52.459 7.441 63.671 ;
      RECT MASK 1 7.761 52.459 7.881 63.671 ;
      RECT MASK 1 8.201 52.459 8.321 63.671 ;
      RECT MASK 1 8.641 52.459 8.761 63.671 ;
      RECT MASK 1 9.081 52.459 9.201 63.671 ;
      RECT MASK 1 9.521 52.459 9.641 63.671 ;
      RECT MASK 1 9.961 52.459 10.081 63.671 ;
      RECT MASK 1 10.401 52.459 10.521 63.671 ;
      RECT MASK 1 10.841 52.459 10.961 63.671 ;
      RECT MASK 1 11.299 52.459 11.419 63.671 ;
      RECT MASK 1 11.739 52.459 11.859 63.671 ;
      RECT MASK 1 12.179 52.459 12.299 63.671 ;
      RECT MASK 1 12.619 52.459 12.739 63.671 ;
      RECT MASK 1 13.059 52.459 13.179 63.671 ;
      RECT MASK 1 13.499 52.459 13.619 63.671 ;
      RECT MASK 1 13.939 52.459 14.059 63.671 ;
      RECT MASK 1 14.379 52.459 14.499 63.671 ;
      RECT MASK 1 14.819 52.459 14.939 63.671 ;
      RECT MASK 1 15.259 52.459 15.379 63.671 ;
      RECT MASK 1 15.699 52.459 15.819 63.671 ;
      RECT MASK 1 16.139 52.459 16.259 63.671 ;
      RECT MASK 1 16.579 52.459 16.699 63.671 ;
      RECT MASK 1 17.019 52.459 17.139 63.671 ;
      RECT MASK 1 17.459 52.459 17.579 63.671 ;
      RECT MASK 1 17.917 52.459 18.037 63.671 ;
      RECT MASK 1 18.357 52.459 18.477 63.671 ;
      RECT MASK 1 18.797 52.459 18.917 63.671 ;
      RECT MASK 1 19.237 52.459 19.357 63.671 ;
      RECT MASK 1 19.677 52.459 19.797 63.671 ;
      RECT MASK 1 20.117 52.459 20.237 63.671 ;
      RECT MASK 1 20.557 52.459 20.677 63.671 ;
      RECT MASK 1 20.997 52.459 21.117 63.671 ;
      RECT MASK 1 21.437 52.459 21.557 63.671 ;
      RECT MASK 1 21.877 52.459 21.997 63.671 ;
      RECT MASK 1 22.317 52.459 22.437 63.671 ;
      RECT MASK 1 22.757 52.459 22.877 63.671 ;
      RECT MASK 1 23.197 52.459 23.317 63.671 ;
      RECT MASK 1 23.637 52.459 23.757 63.671 ;
      RECT MASK 1 24.077 52.459 24.197 63.671 ;
      RECT MASK 1 24.535 52.459 24.655 63.671 ;
      RECT MASK 1 24.975 52.459 25.095 63.671 ;
      RECT MASK 1 25.415 52.459 25.535 63.671 ;
      RECT MASK 1 25.855 52.459 25.975 63.671 ;
      RECT MASK 1 26.295 52.459 26.415 63.671 ;
      RECT MASK 1 26.735 52.459 26.855 63.671 ;
      RECT MASK 1 27.175 52.459 27.295 63.671 ;
      RECT MASK 1 27.615 52.459 27.735 63.671 ;
      RECT MASK 1 28.055 52.459 28.175 63.671 ;
      RECT MASK 1 28.495 52.459 28.615 63.671 ;
      RECT MASK 1 28.935 52.459 29.055 63.671 ;
      RECT MASK 1 29.375 52.459 29.495 63.671 ;
      RECT MASK 1 29.815 52.459 29.935 63.671 ;
      RECT MASK 1 30.255 52.459 30.375 63.671 ;
      RECT MASK 1 30.695 52.459 30.815 63.671 ;
      RECT MASK 1 31.153 52.459 31.273 63.671 ;
      RECT MASK 1 31.593 52.459 31.713 63.671 ;
      RECT MASK 1 32.033 52.459 32.153 63.671 ;
      RECT MASK 1 32.473 52.459 32.593 63.671 ;
      RECT MASK 1 32.913 52.459 33.033 63.671 ;
      RECT MASK 1 33.353 52.459 33.473 63.671 ;
      RECT MASK 1 33.793 52.459 33.913 63.671 ;
      RECT MASK 1 34.233 52.459 34.353 63.671 ;
      RECT MASK 1 34.673 52.459 34.793 63.671 ;
      RECT MASK 1 35.113 52.459 35.233 63.671 ;
      RECT MASK 1 35.553 52.459 35.673 63.671 ;
      RECT MASK 1 35.993 52.459 36.113 63.671 ;
      RECT MASK 1 36.433 52.459 36.553 63.671 ;
      RECT MASK 1 36.873 52.459 36.993 63.671 ;
      RECT MASK 1 37.313 52.459 37.433 63.671 ;
      RECT MASK 1 37.771 52.459 37.891 63.671 ;
      RECT MASK 1 38.211 52.459 38.331 63.671 ;
      RECT MASK 1 38.651 52.459 38.771 63.671 ;
      RECT MASK 1 39.091 52.459 39.211 63.671 ;
      RECT MASK 1 39.531 52.459 39.651 63.671 ;
      RECT MASK 1 39.971 52.459 40.091 63.671 ;
      RECT MASK 1 40.411 52.459 40.531 63.671 ;
      RECT MASK 1 40.851 52.459 40.971 63.671 ;
      RECT MASK 1 41.291 52.459 41.411 63.671 ;
      RECT MASK 1 41.731 52.459 41.851 63.671 ;
      RECT MASK 1 42.171 52.459 42.291 63.671 ;
      RECT MASK 1 42.611 52.459 42.731 63.671 ;
      RECT MASK 1 43.051 52.459 43.171 63.671 ;
      RECT MASK 1 43.491 52.459 43.611 63.671 ;
      RECT MASK 1 43.931 52.459 44.051 63.671 ;
      RECT MASK 1 44.389 52.459 44.509 63.671 ;
      RECT MASK 1 44.829 52.459 44.949 63.671 ;
      RECT MASK 1 45.269 52.459 45.389 63.671 ;
      RECT MASK 1 45.709 52.459 45.829 63.671 ;
      RECT MASK 1 46.149 52.459 46.269 63.671 ;
      RECT MASK 1 46.589 52.459 46.709 63.671 ;
      RECT MASK 1 47.029 52.459 47.149 63.671 ;
      RECT MASK 1 47.469 52.459 47.589 63.671 ;
      RECT MASK 1 47.909 52.459 48.029 63.671 ;
      RECT MASK 1 48.349 52.459 48.469 63.671 ;
      RECT MASK 1 48.789 52.459 48.909 63.671 ;
      RECT MASK 1 49.229 52.459 49.349 63.671 ;
      RECT MASK 1 49.669 52.459 49.789 63.671 ;
      RECT MASK 1 50.109 52.459 50.229 63.671 ;
      RECT MASK 1 50.549 52.459 50.669 63.671 ;
      RECT MASK 1 51.007 52.459 51.127 63.671 ;
      RECT MASK 1 51.447 52.459 51.567 63.671 ;
      RECT MASK 1 51.887 52.459 52.007 63.671 ;
      RECT MASK 1 52.327 52.459 52.447 63.671 ;
      RECT MASK 1 52.767 52.459 52.887 63.671 ;
      RECT MASK 1 53.207 52.459 53.327 63.671 ;
      RECT MASK 1 53.647 52.459 53.767 63.671 ;
      RECT MASK 1 54.087 52.459 54.207 63.671 ;
      RECT MASK 1 54.527 52.459 54.647 63.671 ;
      RECT MASK 1 54.967 52.459 55.087 63.671 ;
      RECT MASK 1 55.407 52.459 55.527 63.671 ;
      RECT MASK 1 55.847 52.459 55.967 63.671 ;
      RECT MASK 1 56.287 52.459 56.407 63.671 ;
      RECT MASK 1 56.727 52.459 56.847 63.671 ;
      RECT MASK 1 57.167 52.459 57.287 63.671 ;
      RECT MASK 1 57.625 52.459 57.745 63.671 ;
      RECT MASK 1 58.065 52.459 58.185 63.671 ;
      RECT MASK 1 58.505 52.459 58.625 63.671 ;
      RECT MASK 1 58.945 52.459 59.065 63.671 ;
      RECT MASK 1 59.385 52.459 59.505 63.671 ;
      RECT MASK 1 59.825 52.459 59.945 63.671 ;
      RECT MASK 1 60.265 52.459 60.385 63.671 ;
      RECT MASK 1 60.705 52.459 60.825 63.671 ;
      RECT MASK 1 61.145 52.459 61.265 63.671 ;
      RECT MASK 1 61.585 52.459 61.705 63.671 ;
      RECT MASK 1 62.025 52.459 62.145 63.671 ;
      RECT MASK 1 62.465 52.459 62.585 63.671 ;
      RECT MASK 1 62.905 52.459 63.025 63.671 ;
      RECT MASK 1 63.345 52.459 63.465 63.671 ;
      RECT MASK 1 63.785 52.459 63.905 63.671 ;
      RECT MASK 1 64.243 52.459 64.363 63.671 ;
      RECT MASK 1 64.683 52.459 64.803 63.671 ;
      RECT MASK 1 65.123 52.459 65.243 63.671 ;
      RECT MASK 1 65.563 52.459 65.683 63.671 ;
      RECT MASK 1 66.003 52.459 66.123 63.671 ;
      RECT MASK 1 66.443 52.459 66.563 63.671 ;
      RECT MASK 1 66.883 52.459 67.003 63.671 ;
      RECT MASK 1 67.323 52.459 67.443 63.671 ;
      RECT MASK 1 67.763 52.459 67.883 63.671 ;
      RECT MASK 1 68.203 52.459 68.323 63.671 ;
      RECT MASK 1 68.643 52.459 68.763 63.671 ;
      RECT MASK 1 69.083 52.459 69.203 63.671 ;
      RECT MASK 1 69.523 52.459 69.643 63.671 ;
      RECT MASK 1 69.963 52.459 70.083 63.671 ;
      RECT MASK 1 70.403 52.459 70.523 63.671 ;
      RECT MASK 1 70.861 52.459 70.981 63.671 ;
      RECT MASK 1 71.301 52.459 71.421 63.671 ;
      RECT MASK 1 71.741 52.459 71.861 63.671 ;
      RECT MASK 1 72.181 52.459 72.301 63.671 ;
      RECT MASK 1 72.621 52.459 72.741 63.671 ;
      RECT MASK 1 73.061 52.459 73.181 63.671 ;
      RECT MASK 1 73.501 52.459 73.621 63.671 ;
      RECT MASK 1 73.941 52.459 74.061 63.671 ;
      RECT MASK 1 74.381 52.459 74.501 63.671 ;
      RECT MASK 1 74.821 52.459 74.941 63.671 ;
      RECT MASK 1 75.261 52.459 75.381 63.671 ;
      RECT MASK 1 75.701 52.459 75.821 63.671 ;
      RECT MASK 1 76.141 52.459 76.261 63.671 ;
      RECT MASK 1 76.581 52.459 76.701 63.671 ;
      RECT MASK 1 77.021 52.459 77.141 63.671 ;
      RECT MASK 1 77.479 52.459 77.599 63.671 ;
      RECT MASK 1 77.919 52.459 78.039 63.671 ;
      RECT MASK 1 78.359 52.459 78.479 63.671 ;
      RECT MASK 1 78.799 52.459 78.919 63.671 ;
      RECT MASK 1 79.239 52.459 79.359 63.671 ;
      RECT MASK 1 79.679 52.459 79.799 63.671 ;
      RECT MASK 1 80.119 52.459 80.239 63.671 ;
      RECT MASK 1 80.559 52.459 80.679 63.671 ;
      RECT MASK 1 80.999 52.459 81.119 63.671 ;
      RECT MASK 1 81.439 52.459 81.559 63.671 ;
      RECT MASK 1 81.879 52.459 81.999 63.671 ;
      RECT MASK 1 82.319 52.459 82.439 63.671 ;
      RECT MASK 1 82.759 52.459 82.879 63.671 ;
      RECT MASK 1 83.199 52.459 83.319 63.671 ;
      RECT MASK 1 83.639 52.459 83.759 63.671 ;
      RECT MASK 1 84.097 52.459 84.217 63.671 ;
      RECT MASK 1 84.537 52.459 84.657 63.671 ;
      RECT MASK 1 84.977 52.459 85.097 63.671 ;
      RECT MASK 1 85.417 52.459 85.537 63.671 ;
      RECT MASK 1 85.857 52.459 85.977 63.671 ;
      RECT MASK 1 86.297 52.459 86.417 63.671 ;
      RECT MASK 1 86.737 52.459 86.857 63.671 ;
      RECT MASK 1 87.177 52.459 87.297 63.671 ;
      RECT MASK 1 87.617 52.459 87.737 63.671 ;
      RECT MASK 1 88.057 52.459 88.177 63.671 ;
      RECT MASK 1 88.497 52.459 88.617 63.671 ;
      RECT MASK 1 88.937 52.459 89.057 63.671 ;
      RECT MASK 1 89.377 52.459 89.497 63.671 ;
      RECT MASK 1 89.817 52.459 89.937 63.671 ;
      RECT MASK 1 90.257 52.459 90.377 63.671 ;
      RECT MASK 1 90.715 52.459 90.835 63.671 ;
      RECT MASK 1 91.155 52.459 91.275 63.671 ;
      RECT MASK 1 91.595 52.459 91.715 63.671 ;
      RECT MASK 1 92.035 52.459 92.155 63.671 ;
      RECT MASK 1 92.475 52.459 92.595 63.671 ;
      RECT MASK 1 92.915 52.459 93.035 63.671 ;
      RECT MASK 1 93.355 52.459 93.475 63.671 ;
      RECT MASK 1 93.795 52.459 93.915 63.671 ;
      RECT MASK 1 94.235 52.459 94.355 63.671 ;
      RECT MASK 1 94.675 52.459 94.795 63.671 ;
      RECT MASK 1 95.115 52.459 95.235 63.671 ;
      RECT MASK 1 95.555 52.459 95.675 63.671 ;
      RECT MASK 1 95.995 52.459 96.115 63.671 ;
      RECT MASK 1 96.435 52.459 96.555 63.671 ;
      RECT MASK 1 96.875 52.459 96.995 63.671 ;
      RECT MASK 1 97.333 52.459 97.453 63.671 ;
      RECT MASK 1 97.773 52.459 97.893 63.671 ;
      RECT MASK 1 98.213 52.459 98.333 63.671 ;
      RECT MASK 1 98.653 52.459 98.773 63.671 ;
      RECT MASK 1 99.093 52.459 99.213 63.671 ;
      RECT MASK 1 99.533 52.459 99.653 63.671 ;
      RECT MASK 1 99.973 52.459 100.093 63.671 ;
      RECT MASK 1 100.413 52.459 100.533 63.671 ;
      RECT MASK 1 100.853 52.459 100.973 63.671 ;
      RECT MASK 1 101.293 52.459 101.413 63.671 ;
      RECT MASK 1 101.733 52.459 101.853 63.671 ;
      RECT MASK 1 102.173 52.459 102.293 63.671 ;
      RECT MASK 1 102.613 52.459 102.733 63.671 ;
      RECT MASK 1 103.053 52.459 103.173 63.671 ;
      RECT MASK 1 103.493 52.459 103.613 63.671 ;
      RECT MASK 1 103.951 52.459 104.071 63.671 ;
      RECT MASK 1 104.391 52.459 104.511 63.671 ;
      RECT MASK 1 104.831 52.459 104.951 63.671 ;
      RECT MASK 1 105.271 52.459 105.391 63.671 ;
      RECT MASK 1 105.711 52.459 105.831 63.671 ;
      RECT MASK 1 106.151 52.459 106.271 63.671 ;
      RECT MASK 1 106.591 52.459 106.711 63.671 ;
      RECT MASK 1 107.031 52.459 107.151 63.671 ;
      RECT MASK 1 107.471 52.459 107.591 63.671 ;
      RECT MASK 1 107.911 52.459 108.031 63.671 ;
      RECT MASK 1 108.351 52.459 108.471 63.671 ;
      RECT MASK 1 108.791 52.459 108.911 63.671 ;
      RECT MASK 1 109.231 52.459 109.351 63.671 ;
      RECT MASK 1 109.671 52.459 109.791 63.671 ;
      RECT MASK 1 110.111 52.459 110.231 63.671 ;
      RECT MASK 1 112.8065 53.149 112.9265 54.179 ;
      RECT MASK 1 113.2465 53.149 113.3665 54.179 ;
      RECT MASK 1 113.6865 53.149 113.8065 54.179 ;
      RECT MASK 1 114.1265 53.149 114.2465 54.179 ;
      RECT MASK 1 114.5665 53.149 114.6865 54.179 ;
      RECT MASK 1 115.0065 53.149 115.1265 54.179 ;
      RECT MASK 1 115.4465 53.149 115.5665 54.179 ;
      RECT MASK 1 115.8865 53.149 116.0065 54.179 ;
      RECT MASK 1 116.3265 53.149 116.4465 54.179 ;
      RECT MASK 1 117.6465 53.149 117.7665 54.179 ;
      RECT MASK 1 118.0865 53.149 118.2065 54.179 ;
      RECT MASK 1 118.5265 53.149 118.6465 54.179 ;
      RECT MASK 1 118.9665 53.149 119.0865 54.179 ;
      RECT MASK 1 119.4065 53.149 119.5265 54.179 ;
      RECT MASK 1 119.8465 53.149 119.9665 54.179 ;
      RECT MASK 1 120.2865 53.149 120.4065 54.179 ;
      RECT MASK 1 120.7265 53.149 120.8465 54.179 ;
      RECT MASK 1 121.1665 53.149 121.2865 54.179 ;
      RECT MASK 1 121.6065 53.149 121.7265 54.179 ;
      RECT MASK 1 122.0465 53.149 122.1665 54.179 ;
      RECT MASK 1 122.4865 53.149 122.6065 54.179 ;
      RECT MASK 1 122.9265 53.149 123.0465 54.179 ;
      RECT MASK 1 112.8065 54.499 112.9265 55.529 ;
      RECT MASK 1 113.2465 54.499 113.3665 55.529 ;
      RECT MASK 1 113.6865 54.499 113.8065 55.529 ;
      RECT MASK 1 114.1265 54.499 114.2465 55.529 ;
      RECT MASK 1 114.5665 54.499 114.6865 55.529 ;
      RECT MASK 1 115.0065 54.499 115.1265 55.529 ;
      RECT MASK 1 115.4465 54.499 115.5665 55.529 ;
      RECT MASK 1 115.8865 54.499 116.0065 55.529 ;
      RECT MASK 1 116.3265 54.499 116.4465 55.529 ;
      RECT MASK 1 112.8065 55.789 112.9265 56.879 ;
      RECT MASK 1 113.2465 55.789 113.3665 56.879 ;
      RECT MASK 1 113.6865 55.789 113.8065 56.879 ;
      RECT MASK 1 114.1265 55.789 114.2465 56.879 ;
      RECT MASK 1 114.5665 55.789 114.6865 56.879 ;
      RECT MASK 1 115.0065 55.789 115.1265 56.879 ;
      RECT MASK 1 115.4465 55.789 115.5665 56.879 ;
      RECT MASK 1 115.8865 55.789 116.0065 56.879 ;
      RECT MASK 1 116.3265 55.789 116.4465 56.879 ;
      RECT MASK 1 117.6465 55.849 117.7665 56.879 ;
      RECT MASK 1 118.0865 55.849 118.2065 56.879 ;
      RECT MASK 1 118.5265 55.849 118.6465 56.879 ;
      RECT MASK 1 118.9665 55.849 119.0865 56.879 ;
      RECT MASK 1 119.4065 55.849 119.5265 56.879 ;
      RECT MASK 1 119.8465 55.849 119.9665 56.879 ;
      RECT MASK 1 120.2865 55.849 120.4065 56.879 ;
      RECT MASK 1 120.7265 55.849 120.8465 56.879 ;
      RECT MASK 1 121.1665 55.849 121.2865 56.879 ;
      RECT MASK 1 121.6065 55.849 121.7265 56.879 ;
      RECT MASK 1 122.0465 55.849 122.1665 56.879 ;
      RECT MASK 1 122.4865 55.849 122.6065 56.879 ;
      RECT MASK 1 122.9265 55.849 123.0465 56.879 ;
      RECT MASK 1 123.3665 55.849 123.4865 56.879 ;
      RECT MASK 1 123.8065 55.849 123.9265 56.879 ;
      RECT MASK 1 112.8065 57.139 112.9265 58.949 ;
      RECT MASK 1 113.2465 57.139 113.3665 58.949 ;
      RECT MASK 1 113.6865 57.139 113.8065 58.949 ;
      RECT MASK 1 114.1265 57.139 114.2465 58.949 ;
      RECT MASK 1 114.5665 57.139 114.6865 58.949 ;
      RECT MASK 1 115.0065 57.139 115.1265 58.949 ;
      RECT MASK 1 115.4465 57.139 115.5665 58.949 ;
      RECT MASK 1 115.8865 57.139 116.0065 58.949 ;
      RECT MASK 1 116.3265 57.139 116.4465 58.949 ;
      RECT MASK 1 117.6465 57.199 117.7665 58.949 ;
      RECT MASK 1 118.0865 57.199 118.2065 58.949 ;
      RECT MASK 1 118.5265 57.199 118.6465 58.949 ;
      RECT MASK 1 118.9665 57.199 119.0865 58.949 ;
      RECT MASK 1 119.4065 57.199 119.5265 58.949 ;
      RECT MASK 1 119.8465 57.199 119.9665 58.949 ;
      RECT MASK 1 120.2865 57.199 120.4065 58.949 ;
      RECT MASK 1 120.7265 57.199 120.8465 58.949 ;
      RECT MASK 1 121.1665 57.199 121.2865 58.949 ;
      RECT MASK 1 121.6065 57.199 121.7265 58.949 ;
      RECT MASK 1 122.0465 57.199 122.1665 58.949 ;
      RECT MASK 1 122.4865 57.199 122.6065 58.949 ;
      RECT MASK 1 122.9265 57.199 123.0465 58.949 ;
      RECT MASK 1 123.3665 57.199 123.4865 58.949 ;
      RECT MASK 1 123.8065 57.199 123.9265 58.949 ;
      RECT MASK 1 112.8065 59.209 112.9265 60.359 ;
      RECT MASK 1 113.2465 59.209 113.3665 60.359 ;
      RECT MASK 1 113.6865 59.209 113.8065 60.359 ;
      RECT MASK 1 114.1265 59.209 114.2465 60.359 ;
      RECT MASK 1 114.5665 59.209 114.6865 60.359 ;
      RECT MASK 1 115.0065 59.209 115.1265 60.359 ;
      RECT MASK 1 115.4465 59.209 115.5665 60.359 ;
      RECT MASK 1 115.8865 59.209 116.0065 60.359 ;
      RECT MASK 1 116.3265 59.209 116.4465 60.359 ;
      RECT MASK 1 117.6465 59.209 117.7665 60.359 ;
      RECT MASK 1 118.0865 59.209 118.2065 60.359 ;
      RECT MASK 1 118.5265 59.209 118.6465 60.359 ;
      RECT MASK 1 118.9665 59.209 119.0865 60.359 ;
      RECT MASK 1 119.4065 59.209 119.5265 60.359 ;
      RECT MASK 1 119.8465 59.209 119.9665 60.359 ;
      RECT MASK 1 120.2865 59.209 120.4065 60.359 ;
      RECT MASK 1 120.7265 59.209 120.8465 60.359 ;
      RECT MASK 1 121.1665 59.209 121.2865 60.359 ;
      RECT MASK 1 121.6065 59.209 121.7265 60.359 ;
      RECT MASK 1 122.0465 59.209 122.1665 60.359 ;
      RECT MASK 1 122.4865 59.209 122.6065 60.359 ;
      RECT MASK 1 122.9265 59.209 123.0465 60.359 ;
      RECT MASK 1 123.3665 59.209 123.4865 60.359 ;
      RECT MASK 1 123.8065 59.209 123.9265 60.359 ;
      RECT MASK 1 112.8065 60.619 112.9265 61.649 ;
      RECT MASK 1 113.2465 60.619 113.3665 61.649 ;
      RECT MASK 1 113.6865 60.619 113.8065 61.649 ;
      RECT MASK 1 114.1265 60.619 114.2465 61.649 ;
      RECT MASK 1 114.5665 60.619 114.6865 61.649 ;
      RECT MASK 1 115.0065 60.619 115.1265 61.649 ;
      RECT MASK 1 115.4465 60.619 115.5665 61.649 ;
      RECT MASK 1 115.8865 60.619 116.0065 61.649 ;
      RECT MASK 1 116.3265 60.619 116.4465 61.649 ;
      RECT MASK 1 117.6465 60.619 117.7665 61.649 ;
      RECT MASK 1 118.0865 60.619 118.2065 61.649 ;
      RECT MASK 1 118.5265 60.619 118.6465 61.649 ;
      RECT MASK 1 118.9665 60.619 119.0865 61.649 ;
      RECT MASK 1 119.4065 60.619 119.5265 61.649 ;
      RECT MASK 1 119.8465 60.619 119.9665 61.649 ;
      RECT MASK 1 120.2865 60.619 120.4065 61.649 ;
      RECT MASK 1 120.7265 60.619 120.8465 61.649 ;
      RECT MASK 1 121.1665 60.619 121.2865 61.649 ;
      RECT MASK 1 121.6065 60.619 121.7265 61.649 ;
      RECT MASK 1 122.0465 60.619 122.1665 61.649 ;
      RECT MASK 1 122.4865 60.619 122.6065 61.649 ;
      RECT MASK 1 122.9265 60.619 123.0465 61.649 ;
      RECT MASK 1 123.3665 60.619 123.4865 61.649 ;
      RECT MASK 1 123.8065 60.619 123.9265 61.649 ;
      RECT MASK 1 112.8065 61.909 112.9265 62.999 ;
      RECT MASK 1 113.2465 61.909 113.3665 62.999 ;
      RECT MASK 1 113.6865 61.909 113.8065 62.999 ;
      RECT MASK 1 114.1265 61.909 114.2465 62.999 ;
      RECT MASK 1 114.5665 61.909 114.6865 62.999 ;
      RECT MASK 1 115.0065 61.909 115.1265 62.999 ;
      RECT MASK 1 115.4465 61.909 115.5665 62.999 ;
      RECT MASK 1 115.8865 61.909 116.0065 62.999 ;
      RECT MASK 1 116.3265 61.909 116.4465 62.999 ;
      RECT MASK 1 117.6465 61.909 117.7665 62.999 ;
      RECT MASK 1 118.0865 61.909 118.2065 62.999 ;
      RECT MASK 1 118.5265 61.909 118.6465 62.999 ;
      RECT MASK 1 118.9665 61.909 119.0865 62.999 ;
      RECT MASK 1 119.4065 61.909 119.5265 62.999 ;
      RECT MASK 1 119.8465 61.909 119.9665 62.999 ;
      RECT MASK 1 120.2865 61.909 120.4065 62.999 ;
      RECT MASK 1 120.7265 61.909 120.8465 62.999 ;
      RECT MASK 1 121.1665 61.909 121.2865 62.999 ;
      RECT MASK 1 121.6065 61.909 121.7265 62.999 ;
      RECT MASK 1 122.0465 61.909 122.1665 62.999 ;
      RECT MASK 1 122.4865 61.909 122.6065 62.999 ;
      RECT MASK 1 122.9265 61.909 123.0465 62.999 ;
      RECT MASK 1 123.3665 61.909 123.4865 62.999 ;
      RECT MASK 1 123.8065 61.909 123.9265 62.999 ;
      RECT MASK 1 112.8065 63.259 112.9265 65.069 ;
      RECT MASK 1 113.2465 63.259 113.3665 65.069 ;
      RECT MASK 1 113.6865 63.259 113.8065 65.069 ;
      RECT MASK 1 114.1265 63.259 114.2465 65.069 ;
      RECT MASK 1 114.5665 63.259 114.6865 65.069 ;
      RECT MASK 1 115.0065 63.259 115.1265 65.069 ;
      RECT MASK 1 115.4465 63.259 115.5665 65.069 ;
      RECT MASK 1 115.8865 63.259 116.0065 65.069 ;
      RECT MASK 1 116.3265 63.259 116.4465 65.069 ;
      RECT MASK 1 117.6465 63.259 117.7665 65.069 ;
      RECT MASK 1 118.0865 63.259 118.2065 65.069 ;
      RECT MASK 1 118.5265 63.259 118.6465 65.069 ;
      RECT MASK 1 118.9665 63.259 119.0865 65.069 ;
      RECT MASK 1 119.4065 63.259 119.5265 65.069 ;
      RECT MASK 1 119.8465 63.259 119.9665 65.069 ;
      RECT MASK 1 120.2865 63.259 120.4065 65.069 ;
      RECT MASK 1 120.7265 63.259 120.8465 65.069 ;
      RECT MASK 1 121.1665 63.259 121.2865 65.069 ;
      RECT MASK 1 121.6065 63.259 121.7265 65.069 ;
      RECT MASK 1 122.0465 63.259 122.1665 65.069 ;
      RECT MASK 1 122.4865 63.259 122.6065 65.069 ;
      RECT MASK 1 122.9265 63.259 123.0465 65.069 ;
      RECT MASK 1 123.3665 63.259 123.4865 65.069 ;
      RECT MASK 1 123.8065 63.259 123.9265 65.069 ;
      RECT MASK 1 4.711 63.84 4.771 64.08 ;
      RECT MASK 1 5.151 63.84 5.211 64.08 ;
      RECT MASK 1 5.591 63.84 5.651 64.08 ;
      RECT MASK 1 6.031 63.84 6.091 64.08 ;
      RECT MASK 1 6.471 63.84 6.531 64.08 ;
      RECT MASK 1 6.911 63.84 6.971 64.08 ;
      RECT MASK 1 7.351 63.84 7.411 64.08 ;
      RECT MASK 1 7.791 63.84 7.851 64.08 ;
      RECT MASK 1 8.231 63.84 8.291 64.08 ;
      RECT MASK 1 8.671 63.84 8.731 64.08 ;
      RECT MASK 1 9.111 63.84 9.171 64.08 ;
      RECT MASK 1 9.551 63.84 9.611 64.08 ;
      RECT MASK 1 9.991 63.84 10.051 64.08 ;
      RECT MASK 1 10.431 63.84 10.491 64.08 ;
      RECT MASK 1 10.871 63.84 10.931 64.08 ;
      RECT MASK 1 11.329 63.84 11.389 64.08 ;
      RECT MASK 1 11.769 63.84 11.829 64.08 ;
      RECT MASK 1 12.209 63.84 12.269 64.08 ;
      RECT MASK 1 12.649 63.84 12.709 64.08 ;
      RECT MASK 1 13.089 63.84 13.149 64.08 ;
      RECT MASK 1 13.529 63.84 13.589 64.08 ;
      RECT MASK 1 13.969 63.84 14.029 64.08 ;
      RECT MASK 1 14.409 63.84 14.469 64.08 ;
      RECT MASK 1 14.849 63.84 14.909 64.08 ;
      RECT MASK 1 15.289 63.84 15.349 64.08 ;
      RECT MASK 1 15.729 63.84 15.789 64.08 ;
      RECT MASK 1 16.169 63.84 16.229 64.08 ;
      RECT MASK 1 16.609 63.84 16.669 64.08 ;
      RECT MASK 1 17.049 63.84 17.109 64.08 ;
      RECT MASK 1 17.489 63.84 17.549 64.08 ;
      RECT MASK 1 17.947 63.84 18.007 64.08 ;
      RECT MASK 1 18.387 63.84 18.447 64.08 ;
      RECT MASK 1 18.827 63.84 18.887 64.08 ;
      RECT MASK 1 19.267 63.84 19.327 64.08 ;
      RECT MASK 1 19.707 63.84 19.767 64.08 ;
      RECT MASK 1 20.147 63.84 20.207 64.08 ;
      RECT MASK 1 20.587 63.84 20.647 64.08 ;
      RECT MASK 1 21.027 63.84 21.087 64.08 ;
      RECT MASK 1 21.467 63.84 21.527 64.08 ;
      RECT MASK 1 21.907 63.84 21.967 64.08 ;
      RECT MASK 1 22.347 63.84 22.407 64.08 ;
      RECT MASK 1 22.787 63.84 22.847 64.08 ;
      RECT MASK 1 23.227 63.84 23.287 64.08 ;
      RECT MASK 1 23.667 63.84 23.727 64.08 ;
      RECT MASK 1 24.107 63.84 24.167 64.08 ;
      RECT MASK 1 24.565 63.84 24.625 64.08 ;
      RECT MASK 1 25.005 63.84 25.065 64.08 ;
      RECT MASK 1 25.445 63.84 25.505 64.08 ;
      RECT MASK 1 25.885 63.84 25.945 64.08 ;
      RECT MASK 1 26.325 63.84 26.385 64.08 ;
      RECT MASK 1 26.765 63.84 26.825 64.08 ;
      RECT MASK 1 27.205 63.84 27.265 64.08 ;
      RECT MASK 1 27.645 63.84 27.705 64.08 ;
      RECT MASK 1 28.085 63.84 28.145 64.08 ;
      RECT MASK 1 28.525 63.84 28.585 64.08 ;
      RECT MASK 1 28.965 63.84 29.025 64.08 ;
      RECT MASK 1 29.405 63.84 29.465 64.08 ;
      RECT MASK 1 29.845 63.84 29.905 64.08 ;
      RECT MASK 1 30.285 63.84 30.345 64.08 ;
      RECT MASK 1 30.725 63.84 30.785 64.08 ;
      RECT MASK 1 31.183 63.84 31.243 64.08 ;
      RECT MASK 1 31.623 63.84 31.683 64.08 ;
      RECT MASK 1 32.063 63.84 32.123 64.08 ;
      RECT MASK 1 32.503 63.84 32.563 64.08 ;
      RECT MASK 1 32.943 63.84 33.003 64.08 ;
      RECT MASK 1 33.383 63.84 33.443 64.08 ;
      RECT MASK 1 33.823 63.84 33.883 64.08 ;
      RECT MASK 1 34.263 63.84 34.323 64.08 ;
      RECT MASK 1 34.703 63.84 34.763 64.08 ;
      RECT MASK 1 35.143 63.84 35.203 64.08 ;
      RECT MASK 1 35.583 63.84 35.643 64.08 ;
      RECT MASK 1 36.023 63.84 36.083 64.08 ;
      RECT MASK 1 36.463 63.84 36.523 64.08 ;
      RECT MASK 1 36.903 63.84 36.963 64.08 ;
      RECT MASK 1 37.343 63.84 37.403 64.08 ;
      RECT MASK 1 37.801 63.84 37.861 64.08 ;
      RECT MASK 1 38.241 63.84 38.301 64.08 ;
      RECT MASK 1 38.681 63.84 38.741 64.08 ;
      RECT MASK 1 39.121 63.84 39.181 64.08 ;
      RECT MASK 1 39.561 63.84 39.621 64.08 ;
      RECT MASK 1 40.001 63.84 40.061 64.08 ;
      RECT MASK 1 40.441 63.84 40.501 64.08 ;
      RECT MASK 1 40.881 63.84 40.941 64.08 ;
      RECT MASK 1 41.321 63.84 41.381 64.08 ;
      RECT MASK 1 41.761 63.84 41.821 64.08 ;
      RECT MASK 1 43.081 63.84 43.141 64.08 ;
      RECT MASK 1 43.521 63.84 43.581 64.08 ;
      RECT MASK 1 43.961 63.84 44.021 64.08 ;
      RECT MASK 1 44.419 63.84 44.479 64.08 ;
      RECT MASK 1 44.859 63.84 44.919 64.08 ;
      RECT MASK 1 45.299 63.84 45.359 64.08 ;
      RECT MASK 1 45.739 63.84 45.799 64.08 ;
      RECT MASK 1 46.179 63.84 46.239 64.08 ;
      RECT MASK 1 46.619 63.84 46.679 64.08 ;
      RECT MASK 1 47.059 63.84 47.119 64.08 ;
      RECT MASK 1 47.499 63.84 47.559 64.08 ;
      RECT MASK 1 47.939 63.84 47.999 64.08 ;
      RECT MASK 1 48.379 63.84 48.439 64.08 ;
      RECT MASK 1 48.819 63.84 48.879 64.08 ;
      RECT MASK 1 49.259 63.84 49.319 64.08 ;
      RECT MASK 1 49.699 63.84 49.759 64.08 ;
      RECT MASK 1 50.139 63.84 50.199 64.08 ;
      RECT MASK 1 50.579 63.84 50.639 64.08 ;
      RECT MASK 1 51.037 63.84 51.097 64.08 ;
      RECT MASK 1 51.477 63.84 51.537 64.08 ;
      RECT MASK 1 51.917 63.84 51.977 64.08 ;
      RECT MASK 1 52.357 63.84 52.417 64.08 ;
      RECT MASK 1 52.797 63.84 52.857 64.08 ;
      RECT MASK 1 53.237 63.84 53.297 64.08 ;
      RECT MASK 1 53.677 63.84 53.737 64.08 ;
      RECT MASK 1 54.117 63.84 54.177 64.08 ;
      RECT MASK 1 54.557 63.84 54.617 64.08 ;
      RECT MASK 1 54.997 63.84 55.057 64.08 ;
      RECT MASK 1 55.437 63.84 55.497 64.08 ;
      RECT MASK 1 55.877 63.84 55.937 64.08 ;
      RECT MASK 1 56.317 63.84 56.377 64.08 ;
      RECT MASK 1 56.757 63.84 56.817 64.08 ;
      RECT MASK 1 57.197 63.84 57.257 64.08 ;
      RECT MASK 1 57.655 63.84 57.715 64.08 ;
      RECT MASK 1 58.095 63.84 58.155 64.08 ;
      RECT MASK 1 58.535 63.84 58.595 64.08 ;
      RECT MASK 1 58.975 63.84 59.035 64.08 ;
      RECT MASK 1 59.415 63.84 59.475 64.08 ;
      RECT MASK 1 59.855 63.84 59.915 64.08 ;
      RECT MASK 1 60.295 63.84 60.355 64.08 ;
      RECT MASK 1 60.735 63.84 60.795 64.08 ;
      RECT MASK 1 61.175 63.84 61.235 64.08 ;
      RECT MASK 1 61.615 63.84 61.675 64.08 ;
      RECT MASK 1 62.055 63.84 62.115 64.08 ;
      RECT MASK 1 62.495 63.84 62.555 64.08 ;
      RECT MASK 1 62.935 63.84 62.995 64.08 ;
      RECT MASK 1 63.375 63.84 63.435 64.08 ;
      RECT MASK 1 63.815 63.84 63.875 64.08 ;
      RECT MASK 1 64.273 63.84 64.333 64.08 ;
      RECT MASK 1 64.713 63.84 64.773 64.08 ;
      RECT MASK 1 65.153 63.84 65.213 64.08 ;
      RECT MASK 1 65.593 63.84 65.653 64.08 ;
      RECT MASK 1 66.033 63.84 66.093 64.08 ;
      RECT MASK 1 66.473 63.84 66.533 64.08 ;
      RECT MASK 1 66.913 63.84 66.973 64.08 ;
      RECT MASK 1 67.353 63.84 67.413 64.08 ;
      RECT MASK 1 67.793 63.84 67.853 64.08 ;
      RECT MASK 1 68.233 63.84 68.293 64.08 ;
      RECT MASK 1 68.673 63.84 68.733 64.08 ;
      RECT MASK 1 69.113 63.84 69.173 64.08 ;
      RECT MASK 1 69.553 63.84 69.613 64.08 ;
      RECT MASK 1 69.993 63.84 70.053 64.08 ;
      RECT MASK 1 70.433 63.84 70.493 64.08 ;
      RECT MASK 1 70.891 63.84 70.951 64.08 ;
      RECT MASK 1 71.331 63.84 71.391 64.08 ;
      RECT MASK 1 71.771 63.84 71.831 64.08 ;
      RECT MASK 1 72.211 63.84 72.271 64.08 ;
      RECT MASK 1 72.651 63.84 72.711 64.08 ;
      RECT MASK 1 73.091 63.84 73.151 64.08 ;
      RECT MASK 1 73.531 63.84 73.591 64.08 ;
      RECT MASK 1 73.971 63.84 74.031 64.08 ;
      RECT MASK 1 74.411 63.84 74.471 64.08 ;
      RECT MASK 1 74.851 63.84 74.911 64.08 ;
      RECT MASK 1 75.291 63.84 75.351 64.08 ;
      RECT MASK 1 75.731 63.84 75.791 64.08 ;
      RECT MASK 1 76.171 63.84 76.231 64.08 ;
      RECT MASK 1 76.611 63.84 76.671 64.08 ;
      RECT MASK 1 77.051 63.84 77.111 64.08 ;
      RECT MASK 1 77.509 63.84 77.569 64.08 ;
      RECT MASK 1 77.949 63.84 78.009 64.08 ;
      RECT MASK 1 78.389 63.84 78.449 64.08 ;
      RECT MASK 1 78.829 63.84 78.889 64.08 ;
      RECT MASK 1 79.269 63.84 79.329 64.08 ;
      RECT MASK 1 79.709 63.84 79.769 64.08 ;
      RECT MASK 1 80.149 63.84 80.209 64.08 ;
      RECT MASK 1 80.589 63.84 80.649 64.08 ;
      RECT MASK 1 81.029 63.84 81.089 64.08 ;
      RECT MASK 1 81.469 63.84 81.529 64.08 ;
      RECT MASK 1 81.909 63.84 81.969 64.08 ;
      RECT MASK 1 82.349 63.84 82.409 64.08 ;
      RECT MASK 1 83.669 63.84 83.729 64.08 ;
      RECT MASK 1 84.127 63.84 84.187 64.08 ;
      RECT MASK 1 84.567 63.84 84.627 64.08 ;
      RECT MASK 1 85.007 63.84 85.067 64.08 ;
      RECT MASK 1 85.447 63.84 85.507 64.08 ;
      RECT MASK 1 85.887 63.84 85.947 64.08 ;
      RECT MASK 1 86.327 63.84 86.387 64.08 ;
      RECT MASK 1 86.767 63.84 86.827 64.08 ;
      RECT MASK 1 87.207 63.84 87.267 64.08 ;
      RECT MASK 1 87.647 63.84 87.707 64.08 ;
      RECT MASK 1 88.087 63.84 88.147 64.08 ;
      RECT MASK 1 88.527 63.84 88.587 64.08 ;
      RECT MASK 1 88.967 63.84 89.027 64.08 ;
      RECT MASK 1 89.407 63.84 89.467 64.08 ;
      RECT MASK 1 89.847 63.84 89.907 64.08 ;
      RECT MASK 1 90.287 63.84 90.347 64.08 ;
      RECT MASK 1 90.745 63.84 90.805 64.08 ;
      RECT MASK 1 91.185 63.84 91.245 64.08 ;
      RECT MASK 1 91.625 63.84 91.685 64.08 ;
      RECT MASK 1 92.065 63.84 92.125 64.08 ;
      RECT MASK 1 92.505 63.84 92.565 64.08 ;
      RECT MASK 1 92.945 63.84 93.005 64.08 ;
      RECT MASK 1 93.385 63.84 93.445 64.08 ;
      RECT MASK 1 93.825 63.84 93.885 64.08 ;
      RECT MASK 1 94.265 63.84 94.325 64.08 ;
      RECT MASK 1 94.705 63.84 94.765 64.08 ;
      RECT MASK 1 95.145 63.84 95.205 64.08 ;
      RECT MASK 1 95.585 63.84 95.645 64.08 ;
      RECT MASK 1 96.025 63.84 96.085 64.08 ;
      RECT MASK 1 96.465 63.84 96.525 64.08 ;
      RECT MASK 1 96.905 63.84 96.965 64.08 ;
      RECT MASK 1 97.363 63.84 97.423 64.08 ;
      RECT MASK 1 97.803 63.84 97.863 64.08 ;
      RECT MASK 1 98.243 63.84 98.303 64.08 ;
      RECT MASK 1 98.683 63.84 98.743 64.08 ;
      RECT MASK 1 99.123 63.84 99.183 64.08 ;
      RECT MASK 1 99.563 63.84 99.623 64.08 ;
      RECT MASK 1 100.003 63.84 100.063 64.08 ;
      RECT MASK 1 100.443 63.84 100.503 64.08 ;
      RECT MASK 1 100.883 63.84 100.943 64.08 ;
      RECT MASK 1 101.323 63.84 101.383 64.08 ;
      RECT MASK 1 101.763 63.84 101.823 64.08 ;
      RECT MASK 1 102.203 63.84 102.263 64.08 ;
      RECT MASK 1 102.643 63.84 102.703 64.08 ;
      RECT MASK 1 103.083 63.84 103.143 64.08 ;
      RECT MASK 1 103.523 63.84 103.583 64.08 ;
      RECT MASK 1 103.981 63.84 104.041 64.08 ;
      RECT MASK 1 104.421 63.84 104.481 64.08 ;
      RECT MASK 1 104.861 63.84 104.921 64.08 ;
      RECT MASK 1 105.301 63.84 105.361 64.08 ;
      RECT MASK 1 105.741 63.84 105.801 64.08 ;
      RECT MASK 1 106.181 63.84 106.241 64.08 ;
      RECT MASK 1 106.621 63.84 106.681 64.08 ;
      RECT MASK 1 107.061 63.84 107.121 64.08 ;
      RECT MASK 1 107.501 63.84 107.561 64.08 ;
      RECT MASK 1 107.941 63.84 108.001 64.08 ;
      RECT MASK 1 108.381 63.84 108.441 64.08 ;
      RECT MASK 1 108.821 63.84 108.881 64.08 ;
      RECT MASK 1 109.261 63.84 109.321 64.08 ;
      RECT MASK 1 109.701 63.84 109.761 64.08 ;
      RECT MASK 1 110.141 63.84 110.201 64.08 ;
      RECT MASK 1 4.711 64.26 4.771 64.5 ;
      RECT MASK 1 5.151 64.26 5.211 64.5 ;
      RECT MASK 1 5.591 64.26 5.651 64.5 ;
      RECT MASK 1 6.031 64.26 6.091 64.5 ;
      RECT MASK 1 6.471 64.26 6.531 64.5 ;
      RECT MASK 1 6.911 64.26 6.971 64.5 ;
      RECT MASK 1 7.351 64.26 7.411 64.5 ;
      RECT MASK 1 7.791 64.26 7.851 64.5 ;
      RECT MASK 1 8.231 64.26 8.291 64.5 ;
      RECT MASK 1 8.671 64.26 8.731 64.5 ;
      RECT MASK 1 9.111 64.26 9.171 64.5 ;
      RECT MASK 1 9.551 64.26 9.611 64.5 ;
      RECT MASK 1 9.991 64.26 10.051 64.5 ;
      RECT MASK 1 10.431 64.26 10.491 64.5 ;
      RECT MASK 1 10.871 64.26 10.931 64.5 ;
      RECT MASK 1 11.329 64.26 11.389 64.5 ;
      RECT MASK 1 11.769 64.26 11.829 64.5 ;
      RECT MASK 1 12.209 64.26 12.269 64.5 ;
      RECT MASK 1 12.649 64.26 12.709 64.5 ;
      RECT MASK 1 13.089 64.26 13.149 64.5 ;
      RECT MASK 1 13.529 64.26 13.589 64.5 ;
      RECT MASK 1 13.969 64.26 14.029 64.5 ;
      RECT MASK 1 14.409 64.26 14.469 64.5 ;
      RECT MASK 1 14.849 64.26 14.909 64.5 ;
      RECT MASK 1 15.289 64.26 15.349 64.5 ;
      RECT MASK 1 15.729 64.26 15.789 64.5 ;
      RECT MASK 1 16.169 64.26 16.229 64.5 ;
      RECT MASK 1 16.609 64.26 16.669 64.5 ;
      RECT MASK 1 17.049 64.26 17.109 64.5 ;
      RECT MASK 1 17.489 64.26 17.549 64.5 ;
      RECT MASK 1 17.947 64.26 18.007 64.5 ;
      RECT MASK 1 18.387 64.26 18.447 64.5 ;
      RECT MASK 1 18.827 64.26 18.887 64.5 ;
      RECT MASK 1 19.267 64.26 19.327 64.5 ;
      RECT MASK 1 19.707 64.26 19.767 64.5 ;
      RECT MASK 1 20.147 64.26 20.207 64.5 ;
      RECT MASK 1 20.587 64.26 20.647 64.5 ;
      RECT MASK 1 21.027 64.26 21.087 64.5 ;
      RECT MASK 1 21.467 64.26 21.527 64.5 ;
      RECT MASK 1 21.907 64.26 21.967 64.5 ;
      RECT MASK 1 22.347 64.26 22.407 64.5 ;
      RECT MASK 1 22.787 64.26 22.847 64.5 ;
      RECT MASK 1 23.227 64.26 23.287 64.5 ;
      RECT MASK 1 23.667 64.26 23.727 64.5 ;
      RECT MASK 1 24.107 64.26 24.167 64.5 ;
      RECT MASK 1 24.565 64.26 24.625 64.5 ;
      RECT MASK 1 25.005 64.26 25.065 64.5 ;
      RECT MASK 1 25.445 64.26 25.505 64.5 ;
      RECT MASK 1 25.885 64.26 25.945 64.5 ;
      RECT MASK 1 26.325 64.26 26.385 64.5 ;
      RECT MASK 1 26.765 64.26 26.825 64.5 ;
      RECT MASK 1 27.205 64.26 27.265 64.5 ;
      RECT MASK 1 27.645 64.26 27.705 64.5 ;
      RECT MASK 1 28.085 64.26 28.145 64.5 ;
      RECT MASK 1 28.525 64.26 28.585 64.5 ;
      RECT MASK 1 28.965 64.26 29.025 64.5 ;
      RECT MASK 1 29.405 64.26 29.465 64.5 ;
      RECT MASK 1 29.845 64.26 29.905 64.5 ;
      RECT MASK 1 30.285 64.26 30.345 64.5 ;
      RECT MASK 1 30.725 64.26 30.785 64.5 ;
      RECT MASK 1 31.183 64.26 31.243 64.5 ;
      RECT MASK 1 31.623 64.26 31.683 64.5 ;
      RECT MASK 1 32.063 64.26 32.123 64.5 ;
      RECT MASK 1 32.503 64.26 32.563 64.5 ;
      RECT MASK 1 32.943 64.26 33.003 64.5 ;
      RECT MASK 1 33.383 64.26 33.443 64.5 ;
      RECT MASK 1 33.823 64.26 33.883 64.5 ;
      RECT MASK 1 34.263 64.26 34.323 64.5 ;
      RECT MASK 1 34.703 64.26 34.763 64.5 ;
      RECT MASK 1 35.143 64.26 35.203 64.5 ;
      RECT MASK 1 35.583 64.26 35.643 64.5 ;
      RECT MASK 1 36.023 64.26 36.083 64.5 ;
      RECT MASK 1 36.463 64.26 36.523 64.5 ;
      RECT MASK 1 36.903 64.26 36.963 64.5 ;
      RECT MASK 1 37.343 64.26 37.403 64.5 ;
      RECT MASK 1 37.801 64.26 37.861 64.5 ;
      RECT MASK 1 38.241 64.26 38.301 64.5 ;
      RECT MASK 1 38.681 64.26 38.741 64.5 ;
      RECT MASK 1 39.121 64.26 39.181 64.5 ;
      RECT MASK 1 39.561 64.26 39.621 64.5 ;
      RECT MASK 1 40.001 64.26 40.061 64.5 ;
      RECT MASK 1 40.441 64.26 40.501 64.5 ;
      RECT MASK 1 40.881 64.26 40.941 64.5 ;
      RECT MASK 1 41.321 64.26 41.381 64.5 ;
      RECT MASK 1 41.761 64.26 41.821 64.5 ;
      RECT MASK 1 43.081 64.26 43.141 64.5 ;
      RECT MASK 1 43.521 64.26 43.581 64.5 ;
      RECT MASK 1 43.961 64.26 44.021 64.5 ;
      RECT MASK 1 44.419 64.26 44.479 64.5 ;
      RECT MASK 1 44.859 64.26 44.919 64.5 ;
      RECT MASK 1 45.299 64.26 45.359 64.5 ;
      RECT MASK 1 45.739 64.26 45.799 64.5 ;
      RECT MASK 1 46.179 64.26 46.239 64.5 ;
      RECT MASK 1 46.619 64.26 46.679 64.5 ;
      RECT MASK 1 47.059 64.26 47.119 64.5 ;
      RECT MASK 1 47.499 64.26 47.559 64.5 ;
      RECT MASK 1 47.939 64.26 47.999 64.5 ;
      RECT MASK 1 48.379 64.26 48.439 64.5 ;
      RECT MASK 1 48.819 64.26 48.879 64.5 ;
      RECT MASK 1 49.259 64.26 49.319 64.5 ;
      RECT MASK 1 49.699 64.26 49.759 64.5 ;
      RECT MASK 1 50.139 64.26 50.199 64.5 ;
      RECT MASK 1 50.579 64.26 50.639 64.5 ;
      RECT MASK 1 51.037 64.26 51.097 64.5 ;
      RECT MASK 1 51.477 64.26 51.537 64.5 ;
      RECT MASK 1 51.917 64.26 51.977 64.5 ;
      RECT MASK 1 52.357 64.26 52.417 64.5 ;
      RECT MASK 1 52.797 64.26 52.857 64.5 ;
      RECT MASK 1 53.237 64.26 53.297 64.5 ;
      RECT MASK 1 53.677 64.26 53.737 64.5 ;
      RECT MASK 1 54.117 64.26 54.177 64.5 ;
      RECT MASK 1 54.557 64.26 54.617 64.5 ;
      RECT MASK 1 54.997 64.26 55.057 64.5 ;
      RECT MASK 1 55.437 64.26 55.497 64.5 ;
      RECT MASK 1 55.877 64.26 55.937 64.5 ;
      RECT MASK 1 56.317 64.26 56.377 64.5 ;
      RECT MASK 1 56.757 64.26 56.817 64.5 ;
      RECT MASK 1 57.197 64.26 57.257 64.5 ;
      RECT MASK 1 57.655 64.26 57.715 64.5 ;
      RECT MASK 1 58.095 64.26 58.155 64.5 ;
      RECT MASK 1 58.535 64.26 58.595 64.5 ;
      RECT MASK 1 58.975 64.26 59.035 64.5 ;
      RECT MASK 1 59.415 64.26 59.475 64.5 ;
      RECT MASK 1 59.855 64.26 59.915 64.5 ;
      RECT MASK 1 60.295 64.26 60.355 64.5 ;
      RECT MASK 1 60.735 64.26 60.795 64.5 ;
      RECT MASK 1 61.175 64.26 61.235 64.5 ;
      RECT MASK 1 61.615 64.26 61.675 64.5 ;
      RECT MASK 1 62.055 64.26 62.115 64.5 ;
      RECT MASK 1 62.495 64.26 62.555 64.5 ;
      RECT MASK 1 62.935 64.26 62.995 64.5 ;
      RECT MASK 1 63.375 64.26 63.435 64.5 ;
      RECT MASK 1 63.815 64.26 63.875 64.5 ;
      RECT MASK 1 64.273 64.26 64.333 64.5 ;
      RECT MASK 1 64.713 64.26 64.773 64.5 ;
      RECT MASK 1 65.153 64.26 65.213 64.5 ;
      RECT MASK 1 65.593 64.26 65.653 64.5 ;
      RECT MASK 1 66.033 64.26 66.093 64.5 ;
      RECT MASK 1 66.473 64.26 66.533 64.5 ;
      RECT MASK 1 66.913 64.26 66.973 64.5 ;
      RECT MASK 1 67.353 64.26 67.413 64.5 ;
      RECT MASK 1 67.793 64.26 67.853 64.5 ;
      RECT MASK 1 68.233 64.26 68.293 64.5 ;
      RECT MASK 1 68.673 64.26 68.733 64.5 ;
      RECT MASK 1 69.113 64.26 69.173 64.5 ;
      RECT MASK 1 69.553 64.26 69.613 64.5 ;
      RECT MASK 1 69.993 64.26 70.053 64.5 ;
      RECT MASK 1 70.433 64.26 70.493 64.5 ;
      RECT MASK 1 70.891 64.26 70.951 64.5 ;
      RECT MASK 1 71.331 64.26 71.391 64.5 ;
      RECT MASK 1 71.771 64.26 71.831 64.5 ;
      RECT MASK 1 72.211 64.26 72.271 64.5 ;
      RECT MASK 1 72.651 64.26 72.711 64.5 ;
      RECT MASK 1 73.091 64.26 73.151 64.5 ;
      RECT MASK 1 73.531 64.26 73.591 64.5 ;
      RECT MASK 1 73.971 64.26 74.031 64.5 ;
      RECT MASK 1 74.411 64.26 74.471 64.5 ;
      RECT MASK 1 74.851 64.26 74.911 64.5 ;
      RECT MASK 1 75.291 64.26 75.351 64.5 ;
      RECT MASK 1 75.731 64.26 75.791 64.5 ;
      RECT MASK 1 76.171 64.26 76.231 64.5 ;
      RECT MASK 1 76.611 64.26 76.671 64.5 ;
      RECT MASK 1 77.051 64.26 77.111 64.5 ;
      RECT MASK 1 77.509 64.26 77.569 64.5 ;
      RECT MASK 1 77.949 64.26 78.009 64.5 ;
      RECT MASK 1 78.389 64.26 78.449 64.5 ;
      RECT MASK 1 78.829 64.26 78.889 64.5 ;
      RECT MASK 1 79.269 64.26 79.329 64.5 ;
      RECT MASK 1 79.709 64.26 79.769 64.5 ;
      RECT MASK 1 80.149 64.26 80.209 64.5 ;
      RECT MASK 1 80.589 64.26 80.649 64.5 ;
      RECT MASK 1 81.029 64.26 81.089 64.5 ;
      RECT MASK 1 81.469 64.26 81.529 64.5 ;
      RECT MASK 1 81.909 64.26 81.969 64.5 ;
      RECT MASK 1 82.349 64.26 82.409 64.5 ;
      RECT MASK 1 83.669 64.26 83.729 64.5 ;
      RECT MASK 1 84.127 64.26 84.187 64.5 ;
      RECT MASK 1 84.567 64.26 84.627 64.5 ;
      RECT MASK 1 85.007 64.26 85.067 64.5 ;
      RECT MASK 1 85.447 64.26 85.507 64.5 ;
      RECT MASK 1 85.887 64.26 85.947 64.5 ;
      RECT MASK 1 86.327 64.26 86.387 64.5 ;
      RECT MASK 1 86.767 64.26 86.827 64.5 ;
      RECT MASK 1 87.207 64.26 87.267 64.5 ;
      RECT MASK 1 87.647 64.26 87.707 64.5 ;
      RECT MASK 1 88.087 64.26 88.147 64.5 ;
      RECT MASK 1 88.527 64.26 88.587 64.5 ;
      RECT MASK 1 88.967 64.26 89.027 64.5 ;
      RECT MASK 1 89.407 64.26 89.467 64.5 ;
      RECT MASK 1 89.847 64.26 89.907 64.5 ;
      RECT MASK 1 90.287 64.26 90.347 64.5 ;
      RECT MASK 1 90.745 64.26 90.805 64.5 ;
      RECT MASK 1 91.185 64.26 91.245 64.5 ;
      RECT MASK 1 91.625 64.26 91.685 64.5 ;
      RECT MASK 1 92.065 64.26 92.125 64.5 ;
      RECT MASK 1 92.505 64.26 92.565 64.5 ;
      RECT MASK 1 92.945 64.26 93.005 64.5 ;
      RECT MASK 1 93.385 64.26 93.445 64.5 ;
      RECT MASK 1 93.825 64.26 93.885 64.5 ;
      RECT MASK 1 94.265 64.26 94.325 64.5 ;
      RECT MASK 1 94.705 64.26 94.765 64.5 ;
      RECT MASK 1 95.145 64.26 95.205 64.5 ;
      RECT MASK 1 95.585 64.26 95.645 64.5 ;
      RECT MASK 1 96.025 64.26 96.085 64.5 ;
      RECT MASK 1 96.465 64.26 96.525 64.5 ;
      RECT MASK 1 96.905 64.26 96.965 64.5 ;
      RECT MASK 1 97.363 64.26 97.423 64.5 ;
      RECT MASK 1 97.803 64.26 97.863 64.5 ;
      RECT MASK 1 98.243 64.26 98.303 64.5 ;
      RECT MASK 1 98.683 64.26 98.743 64.5 ;
      RECT MASK 1 99.123 64.26 99.183 64.5 ;
      RECT MASK 1 99.563 64.26 99.623 64.5 ;
      RECT MASK 1 100.003 64.26 100.063 64.5 ;
      RECT MASK 1 100.443 64.26 100.503 64.5 ;
      RECT MASK 1 100.883 64.26 100.943 64.5 ;
      RECT MASK 1 101.323 64.26 101.383 64.5 ;
      RECT MASK 1 101.763 64.26 101.823 64.5 ;
      RECT MASK 1 102.203 64.26 102.263 64.5 ;
      RECT MASK 1 102.643 64.26 102.703 64.5 ;
      RECT MASK 1 103.083 64.26 103.143 64.5 ;
      RECT MASK 1 103.523 64.26 103.583 64.5 ;
      RECT MASK 1 103.981 64.26 104.041 64.5 ;
      RECT MASK 1 104.421 64.26 104.481 64.5 ;
      RECT MASK 1 104.861 64.26 104.921 64.5 ;
      RECT MASK 1 105.301 64.26 105.361 64.5 ;
      RECT MASK 1 105.741 64.26 105.801 64.5 ;
      RECT MASK 1 106.181 64.26 106.241 64.5 ;
      RECT MASK 1 106.621 64.26 106.681 64.5 ;
      RECT MASK 1 107.061 64.26 107.121 64.5 ;
      RECT MASK 1 107.501 64.26 107.561 64.5 ;
      RECT MASK 1 107.941 64.26 108.001 64.5 ;
      RECT MASK 1 108.381 64.26 108.441 64.5 ;
      RECT MASK 1 108.821 64.26 108.881 64.5 ;
      RECT MASK 1 109.261 64.26 109.321 64.5 ;
      RECT MASK 1 109.701 64.26 109.761 64.5 ;
      RECT MASK 1 110.141 64.26 110.201 64.5 ;
      RECT MASK 1 4.681 64.699 4.801 75.911 ;
      RECT MASK 1 5.121 64.699 5.241 75.911 ;
      RECT MASK 1 5.561 64.699 5.681 75.911 ;
      RECT MASK 1 6.001 64.699 6.121 75.911 ;
      RECT MASK 1 6.441 64.699 6.561 75.911 ;
      RECT MASK 1 6.881 64.699 7.001 75.911 ;
      RECT MASK 1 7.321 64.699 7.441 75.911 ;
      RECT MASK 1 7.761 64.699 7.881 75.911 ;
      RECT MASK 1 8.201 64.699 8.321 75.911 ;
      RECT MASK 1 8.641 64.699 8.761 75.911 ;
      RECT MASK 1 9.081 64.699 9.201 75.911 ;
      RECT MASK 1 9.521 64.699 9.641 75.911 ;
      RECT MASK 1 9.961 64.699 10.081 75.911 ;
      RECT MASK 1 10.401 64.699 10.521 75.911 ;
      RECT MASK 1 10.841 64.699 10.961 75.911 ;
      RECT MASK 1 11.299 64.699 11.419 75.911 ;
      RECT MASK 1 11.739 64.699 11.859 75.911 ;
      RECT MASK 1 12.179 64.699 12.299 75.911 ;
      RECT MASK 1 12.619 64.699 12.739 75.911 ;
      RECT MASK 1 13.059 64.699 13.179 75.911 ;
      RECT MASK 1 13.499 64.699 13.619 75.911 ;
      RECT MASK 1 13.939 64.699 14.059 75.911 ;
      RECT MASK 1 14.379 64.699 14.499 75.911 ;
      RECT MASK 1 14.819 64.699 14.939 75.911 ;
      RECT MASK 1 15.259 64.699 15.379 75.911 ;
      RECT MASK 1 15.699 64.699 15.819 75.911 ;
      RECT MASK 1 16.139 64.699 16.259 75.911 ;
      RECT MASK 1 16.579 64.699 16.699 75.911 ;
      RECT MASK 1 17.019 64.699 17.139 75.911 ;
      RECT MASK 1 17.459 64.699 17.579 75.911 ;
      RECT MASK 1 17.917 64.699 18.037 75.911 ;
      RECT MASK 1 18.357 64.699 18.477 75.911 ;
      RECT MASK 1 18.797 64.699 18.917 75.911 ;
      RECT MASK 1 19.237 64.699 19.357 75.911 ;
      RECT MASK 1 19.677 64.699 19.797 75.911 ;
      RECT MASK 1 20.117 64.699 20.237 75.911 ;
      RECT MASK 1 20.557 64.699 20.677 75.911 ;
      RECT MASK 1 20.997 64.699 21.117 75.911 ;
      RECT MASK 1 21.437 64.699 21.557 75.911 ;
      RECT MASK 1 21.877 64.699 21.997 75.911 ;
      RECT MASK 1 22.317 64.699 22.437 75.911 ;
      RECT MASK 1 22.757 64.699 22.877 75.911 ;
      RECT MASK 1 23.197 64.699 23.317 75.911 ;
      RECT MASK 1 23.637 64.699 23.757 75.911 ;
      RECT MASK 1 24.077 64.699 24.197 75.911 ;
      RECT MASK 1 24.535 64.699 24.655 75.911 ;
      RECT MASK 1 24.975 64.699 25.095 75.911 ;
      RECT MASK 1 25.415 64.699 25.535 75.911 ;
      RECT MASK 1 25.855 64.699 25.975 75.911 ;
      RECT MASK 1 26.295 64.699 26.415 75.911 ;
      RECT MASK 1 26.735 64.699 26.855 75.911 ;
      RECT MASK 1 27.175 64.699 27.295 75.911 ;
      RECT MASK 1 27.615 64.699 27.735 75.911 ;
      RECT MASK 1 28.055 64.699 28.175 75.911 ;
      RECT MASK 1 28.495 64.699 28.615 75.911 ;
      RECT MASK 1 28.935 64.699 29.055 75.911 ;
      RECT MASK 1 29.375 64.699 29.495 75.911 ;
      RECT MASK 1 29.815 64.699 29.935 75.911 ;
      RECT MASK 1 30.255 64.699 30.375 75.911 ;
      RECT MASK 1 30.695 64.699 30.815 75.911 ;
      RECT MASK 1 31.153 64.699 31.273 75.911 ;
      RECT MASK 1 31.593 64.699 31.713 75.911 ;
      RECT MASK 1 32.033 64.699 32.153 75.911 ;
      RECT MASK 1 32.473 64.699 32.593 75.911 ;
      RECT MASK 1 32.913 64.699 33.033 75.911 ;
      RECT MASK 1 33.353 64.699 33.473 75.911 ;
      RECT MASK 1 33.793 64.699 33.913 75.911 ;
      RECT MASK 1 34.233 64.699 34.353 75.911 ;
      RECT MASK 1 34.673 64.699 34.793 75.911 ;
      RECT MASK 1 35.113 64.699 35.233 75.911 ;
      RECT MASK 1 35.553 64.699 35.673 75.911 ;
      RECT MASK 1 35.993 64.699 36.113 75.911 ;
      RECT MASK 1 36.433 64.699 36.553 75.911 ;
      RECT MASK 1 36.873 64.699 36.993 75.911 ;
      RECT MASK 1 37.313 64.699 37.433 75.911 ;
      RECT MASK 1 37.771 64.699 37.891 75.911 ;
      RECT MASK 1 38.211 64.699 38.331 75.911 ;
      RECT MASK 1 38.651 64.699 38.771 75.911 ;
      RECT MASK 1 39.091 64.699 39.211 75.911 ;
      RECT MASK 1 39.531 64.699 39.651 75.911 ;
      RECT MASK 1 39.971 64.699 40.091 75.911 ;
      RECT MASK 1 40.411 64.699 40.531 75.911 ;
      RECT MASK 1 40.851 64.699 40.971 75.911 ;
      RECT MASK 1 41.291 64.699 41.411 75.911 ;
      RECT MASK 1 41.731 64.699 41.851 75.911 ;
      RECT MASK 1 42.171 64.699 42.291 75.911 ;
      RECT MASK 1 42.611 64.699 42.731 75.911 ;
      RECT MASK 1 43.051 64.699 43.171 75.911 ;
      RECT MASK 1 43.491 64.699 43.611 75.911 ;
      RECT MASK 1 43.931 64.699 44.051 75.911 ;
      RECT MASK 1 44.389 64.699 44.509 75.911 ;
      RECT MASK 1 44.829 64.699 44.949 75.911 ;
      RECT MASK 1 45.269 64.699 45.389 75.911 ;
      RECT MASK 1 45.709 64.699 45.829 75.911 ;
      RECT MASK 1 46.149 64.699 46.269 75.911 ;
      RECT MASK 1 46.589 64.699 46.709 75.911 ;
      RECT MASK 1 47.029 64.699 47.149 75.911 ;
      RECT MASK 1 47.469 64.699 47.589 75.911 ;
      RECT MASK 1 47.909 64.699 48.029 75.911 ;
      RECT MASK 1 48.349 64.699 48.469 75.911 ;
      RECT MASK 1 48.789 64.699 48.909 75.911 ;
      RECT MASK 1 49.229 64.699 49.349 75.911 ;
      RECT MASK 1 49.669 64.699 49.789 75.911 ;
      RECT MASK 1 50.109 64.699 50.229 75.911 ;
      RECT MASK 1 50.549 64.699 50.669 75.911 ;
      RECT MASK 1 51.007 64.699 51.127 75.911 ;
      RECT MASK 1 51.447 64.699 51.567 75.911 ;
      RECT MASK 1 51.887 64.699 52.007 75.911 ;
      RECT MASK 1 52.327 64.699 52.447 75.911 ;
      RECT MASK 1 52.767 64.699 52.887 75.911 ;
      RECT MASK 1 53.207 64.699 53.327 75.911 ;
      RECT MASK 1 53.647 64.699 53.767 75.911 ;
      RECT MASK 1 54.087 64.699 54.207 75.911 ;
      RECT MASK 1 54.527 64.699 54.647 75.911 ;
      RECT MASK 1 54.967 64.699 55.087 75.911 ;
      RECT MASK 1 55.407 64.699 55.527 75.911 ;
      RECT MASK 1 55.847 64.699 55.967 75.911 ;
      RECT MASK 1 56.287 64.699 56.407 75.911 ;
      RECT MASK 1 56.727 64.699 56.847 75.911 ;
      RECT MASK 1 57.167 64.699 57.287 75.911 ;
      RECT MASK 1 57.625 64.699 57.745 75.911 ;
      RECT MASK 1 58.065 64.699 58.185 75.911 ;
      RECT MASK 1 58.505 64.699 58.625 75.911 ;
      RECT MASK 1 58.945 64.699 59.065 75.911 ;
      RECT MASK 1 59.385 64.699 59.505 75.911 ;
      RECT MASK 1 59.825 64.699 59.945 75.911 ;
      RECT MASK 1 60.265 64.699 60.385 75.911 ;
      RECT MASK 1 60.705 64.699 60.825 75.911 ;
      RECT MASK 1 61.145 64.699 61.265 75.911 ;
      RECT MASK 1 61.585 64.699 61.705 75.911 ;
      RECT MASK 1 62.025 64.699 62.145 75.911 ;
      RECT MASK 1 62.465 64.699 62.585 75.911 ;
      RECT MASK 1 62.905 64.699 63.025 75.911 ;
      RECT MASK 1 63.345 64.699 63.465 75.911 ;
      RECT MASK 1 63.785 64.699 63.905 75.911 ;
      RECT MASK 1 64.243 64.699 64.363 75.911 ;
      RECT MASK 1 64.683 64.699 64.803 75.911 ;
      RECT MASK 1 65.123 64.699 65.243 75.911 ;
      RECT MASK 1 65.563 64.699 65.683 75.911 ;
      RECT MASK 1 66.003 64.699 66.123 75.911 ;
      RECT MASK 1 66.443 64.699 66.563 75.911 ;
      RECT MASK 1 66.883 64.699 67.003 75.911 ;
      RECT MASK 1 67.323 64.699 67.443 75.911 ;
      RECT MASK 1 67.763 64.699 67.883 75.911 ;
      RECT MASK 1 68.203 64.699 68.323 75.911 ;
      RECT MASK 1 68.643 64.699 68.763 75.911 ;
      RECT MASK 1 69.083 64.699 69.203 75.911 ;
      RECT MASK 1 69.523 64.699 69.643 75.911 ;
      RECT MASK 1 69.963 64.699 70.083 75.911 ;
      RECT MASK 1 70.403 64.699 70.523 75.911 ;
      RECT MASK 1 70.861 64.699 70.981 75.911 ;
      RECT MASK 1 71.301 64.699 71.421 75.911 ;
      RECT MASK 1 71.741 64.699 71.861 75.911 ;
      RECT MASK 1 72.181 64.699 72.301 75.911 ;
      RECT MASK 1 72.621 64.699 72.741 75.911 ;
      RECT MASK 1 73.061 64.699 73.181 75.911 ;
      RECT MASK 1 73.501 64.699 73.621 75.911 ;
      RECT MASK 1 73.941 64.699 74.061 75.911 ;
      RECT MASK 1 74.381 64.699 74.501 75.911 ;
      RECT MASK 1 74.821 64.699 74.941 75.911 ;
      RECT MASK 1 75.261 64.699 75.381 75.911 ;
      RECT MASK 1 75.701 64.699 75.821 75.911 ;
      RECT MASK 1 76.141 64.699 76.261 75.911 ;
      RECT MASK 1 76.581 64.699 76.701 75.911 ;
      RECT MASK 1 77.021 64.699 77.141 75.911 ;
      RECT MASK 1 77.479 64.699 77.599 75.911 ;
      RECT MASK 1 77.919 64.699 78.039 75.911 ;
      RECT MASK 1 78.359 64.699 78.479 75.911 ;
      RECT MASK 1 78.799 64.699 78.919 75.911 ;
      RECT MASK 1 79.239 64.699 79.359 75.911 ;
      RECT MASK 1 79.679 64.699 79.799 75.911 ;
      RECT MASK 1 80.119 64.699 80.239 75.911 ;
      RECT MASK 1 80.559 64.699 80.679 75.911 ;
      RECT MASK 1 80.999 64.699 81.119 75.911 ;
      RECT MASK 1 81.439 64.699 81.559 75.911 ;
      RECT MASK 1 81.879 64.699 81.999 75.911 ;
      RECT MASK 1 82.319 64.699 82.439 75.911 ;
      RECT MASK 1 82.759 64.699 82.879 75.911 ;
      RECT MASK 1 83.199 64.699 83.319 75.911 ;
      RECT MASK 1 83.639 64.699 83.759 75.911 ;
      RECT MASK 1 84.097 64.699 84.217 75.911 ;
      RECT MASK 1 84.537 64.699 84.657 75.911 ;
      RECT MASK 1 84.977 64.699 85.097 75.911 ;
      RECT MASK 1 85.417 64.699 85.537 75.911 ;
      RECT MASK 1 85.857 64.699 85.977 75.911 ;
      RECT MASK 1 86.297 64.699 86.417 75.911 ;
      RECT MASK 1 86.737 64.699 86.857 75.911 ;
      RECT MASK 1 87.177 64.699 87.297 75.911 ;
      RECT MASK 1 87.617 64.699 87.737 75.911 ;
      RECT MASK 1 88.057 64.699 88.177 75.911 ;
      RECT MASK 1 88.497 64.699 88.617 75.911 ;
      RECT MASK 1 88.937 64.699 89.057 75.911 ;
      RECT MASK 1 89.377 64.699 89.497 75.911 ;
      RECT MASK 1 89.817 64.699 89.937 75.911 ;
      RECT MASK 1 90.257 64.699 90.377 75.911 ;
      RECT MASK 1 90.715 64.699 90.835 75.911 ;
      RECT MASK 1 91.155 64.699 91.275 75.911 ;
      RECT MASK 1 91.595 64.699 91.715 75.911 ;
      RECT MASK 1 92.035 64.699 92.155 75.911 ;
      RECT MASK 1 92.475 64.699 92.595 75.911 ;
      RECT MASK 1 92.915 64.699 93.035 75.911 ;
      RECT MASK 1 93.355 64.699 93.475 75.911 ;
      RECT MASK 1 93.795 64.699 93.915 75.911 ;
      RECT MASK 1 94.235 64.699 94.355 75.911 ;
      RECT MASK 1 94.675 64.699 94.795 75.911 ;
      RECT MASK 1 95.115 64.699 95.235 75.911 ;
      RECT MASK 1 95.555 64.699 95.675 75.911 ;
      RECT MASK 1 95.995 64.699 96.115 75.911 ;
      RECT MASK 1 96.435 64.699 96.555 75.911 ;
      RECT MASK 1 96.875 64.699 96.995 75.911 ;
      RECT MASK 1 97.333 64.699 97.453 75.911 ;
      RECT MASK 1 97.773 64.699 97.893 75.911 ;
      RECT MASK 1 98.213 64.699 98.333 75.911 ;
      RECT MASK 1 98.653 64.699 98.773 75.911 ;
      RECT MASK 1 99.093 64.699 99.213 75.911 ;
      RECT MASK 1 99.533 64.699 99.653 75.911 ;
      RECT MASK 1 99.973 64.699 100.093 75.911 ;
      RECT MASK 1 100.413 64.699 100.533 75.911 ;
      RECT MASK 1 100.853 64.699 100.973 75.911 ;
      RECT MASK 1 101.293 64.699 101.413 75.911 ;
      RECT MASK 1 101.733 64.699 101.853 75.911 ;
      RECT MASK 1 102.173 64.699 102.293 75.911 ;
      RECT MASK 1 102.613 64.699 102.733 75.911 ;
      RECT MASK 1 103.053 64.699 103.173 75.911 ;
      RECT MASK 1 103.493 64.699 103.613 75.911 ;
      RECT MASK 1 103.951 64.699 104.071 75.911 ;
      RECT MASK 1 104.391 64.699 104.511 75.911 ;
      RECT MASK 1 104.831 64.699 104.951 75.911 ;
      RECT MASK 1 105.271 64.699 105.391 75.911 ;
      RECT MASK 1 105.711 64.699 105.831 75.911 ;
      RECT MASK 1 106.151 64.699 106.271 75.911 ;
      RECT MASK 1 106.591 64.699 106.711 75.911 ;
      RECT MASK 1 107.031 64.699 107.151 75.911 ;
      RECT MASK 1 107.471 64.699 107.591 75.911 ;
      RECT MASK 1 107.911 64.699 108.031 75.911 ;
      RECT MASK 1 108.351 64.699 108.471 75.911 ;
      RECT MASK 1 108.791 64.699 108.911 75.911 ;
      RECT MASK 1 109.231 64.699 109.351 75.911 ;
      RECT MASK 1 109.671 64.699 109.791 75.911 ;
      RECT MASK 1 110.111 64.699 110.231 75.911 ;
      RECT MASK 1 112.8065 65.329 112.9265 66.419 ;
      RECT MASK 1 113.2465 65.329 113.3665 66.419 ;
      RECT MASK 1 113.6865 65.329 113.8065 66.419 ;
      RECT MASK 1 114.1265 65.329 114.2465 66.419 ;
      RECT MASK 1 114.5665 65.329 114.6865 66.419 ;
      RECT MASK 1 115.0065 65.329 115.1265 66.419 ;
      RECT MASK 1 115.4465 65.329 115.5665 66.419 ;
      RECT MASK 1 115.8865 65.329 116.0065 66.419 ;
      RECT MASK 1 116.3265 65.329 116.4465 66.419 ;
      RECT MASK 1 117.6465 65.329 117.7665 66.419 ;
      RECT MASK 1 118.0865 65.329 118.2065 66.419 ;
      RECT MASK 1 118.5265 65.329 118.6465 66.419 ;
      RECT MASK 1 118.9665 65.329 119.0865 66.419 ;
      RECT MASK 1 119.4065 65.329 119.5265 66.419 ;
      RECT MASK 1 119.8465 65.329 119.9665 66.419 ;
      RECT MASK 1 120.2865 65.329 120.4065 66.419 ;
      RECT MASK 1 120.7265 65.329 120.8465 66.419 ;
      RECT MASK 1 121.1665 65.329 121.2865 66.419 ;
      RECT MASK 1 121.6065 65.329 121.7265 66.419 ;
      RECT MASK 1 122.0465 65.329 122.1665 66.419 ;
      RECT MASK 1 122.4865 65.329 122.6065 66.419 ;
      RECT MASK 1 122.9265 65.329 123.0465 66.419 ;
      RECT MASK 1 123.3665 65.329 123.4865 66.419 ;
      RECT MASK 1 123.8065 65.329 123.9265 66.419 ;
      RECT MASK 1 112.8065 66.679 112.9265 67.769 ;
      RECT MASK 1 113.2465 66.679 113.3665 67.769 ;
      RECT MASK 1 113.6865 66.679 113.8065 67.769 ;
      RECT MASK 1 114.1265 66.679 114.2465 67.769 ;
      RECT MASK 1 114.5665 66.679 114.6865 67.769 ;
      RECT MASK 1 115.0065 66.679 115.1265 67.769 ;
      RECT MASK 1 115.4465 66.679 115.5665 67.769 ;
      RECT MASK 1 115.8865 66.679 116.0065 67.769 ;
      RECT MASK 1 116.3265 66.679 116.4465 67.769 ;
      RECT MASK 1 117.6465 66.679 117.7665 67.769 ;
      RECT MASK 1 118.0865 66.679 118.2065 67.769 ;
      RECT MASK 1 118.5265 66.679 118.6465 67.769 ;
      RECT MASK 1 118.9665 66.679 119.0865 67.769 ;
      RECT MASK 1 119.4065 66.679 119.5265 67.769 ;
      RECT MASK 1 119.8465 66.679 119.9665 67.769 ;
      RECT MASK 1 120.2865 66.679 120.4065 67.769 ;
      RECT MASK 1 120.7265 66.679 120.8465 67.769 ;
      RECT MASK 1 121.1665 66.679 121.2865 67.769 ;
      RECT MASK 1 121.6065 66.679 121.7265 67.769 ;
      RECT MASK 1 122.0465 66.679 122.1665 67.769 ;
      RECT MASK 1 122.4865 66.679 122.6065 67.769 ;
      RECT MASK 1 122.9265 66.679 123.0465 67.769 ;
      RECT MASK 1 123.3665 66.679 123.4865 67.769 ;
      RECT MASK 1 123.8065 66.679 123.9265 67.769 ;
      RECT MASK 1 112.8065 68.029 112.9265 69.119 ;
      RECT MASK 1 113.2465 68.029 113.3665 69.119 ;
      RECT MASK 1 113.6865 68.029 113.8065 69.119 ;
      RECT MASK 1 114.1265 68.029 114.2465 69.119 ;
      RECT MASK 1 114.5665 68.029 114.6865 69.119 ;
      RECT MASK 1 115.0065 68.029 115.1265 69.119 ;
      RECT MASK 1 115.4465 68.029 115.5665 69.119 ;
      RECT MASK 1 115.8865 68.029 116.0065 69.119 ;
      RECT MASK 1 116.3265 68.029 116.4465 69.119 ;
      RECT MASK 1 117.6465 68.029 117.7665 69.119 ;
      RECT MASK 1 118.0865 68.029 118.2065 69.119 ;
      RECT MASK 1 118.5265 68.029 118.6465 69.119 ;
      RECT MASK 1 118.9665 68.029 119.0865 69.119 ;
      RECT MASK 1 119.4065 68.029 119.5265 69.119 ;
      RECT MASK 1 119.8465 68.029 119.9665 69.119 ;
      RECT MASK 1 120.2865 68.029 120.4065 69.119 ;
      RECT MASK 1 120.7265 68.029 120.8465 69.119 ;
      RECT MASK 1 121.1665 68.029 121.2865 69.119 ;
      RECT MASK 1 121.6065 68.029 121.7265 69.119 ;
      RECT MASK 1 122.0465 68.029 122.1665 69.119 ;
      RECT MASK 1 122.4865 68.029 122.6065 69.119 ;
      RECT MASK 1 122.9265 68.029 123.0465 69.119 ;
      RECT MASK 1 123.3665 68.029 123.4865 69.119 ;
      RECT MASK 1 123.8065 68.029 123.9265 69.119 ;
      RECT MASK 1 112.8065 69.379 112.9265 71.189 ;
      RECT MASK 1 114.5665 69.379 114.6865 71.189 ;
      RECT MASK 1 115.0065 69.379 115.1265 71.189 ;
      RECT MASK 1 115.4465 69.379 115.5665 71.189 ;
      RECT MASK 1 115.8865 69.379 116.0065 71.189 ;
      RECT MASK 1 116.3265 69.379 116.4465 71.189 ;
      RECT MASK 1 117.6465 69.379 117.7665 71.189 ;
      RECT MASK 1 118.0865 69.379 118.2065 71.189 ;
      RECT MASK 1 118.5265 69.379 118.6465 71.189 ;
      RECT MASK 1 118.9665 69.379 119.0865 71.189 ;
      RECT MASK 1 119.4065 69.379 119.5265 71.189 ;
      RECT MASK 1 119.8465 69.379 119.9665 71.189 ;
      RECT MASK 1 120.2865 69.379 120.4065 71.189 ;
      RECT MASK 1 120.7265 69.379 120.8465 71.189 ;
      RECT MASK 1 121.1665 69.379 121.2865 71.189 ;
      RECT MASK 1 121.6065 69.379 121.7265 71.189 ;
      RECT MASK 1 122.0465 69.379 122.1665 71.189 ;
      RECT MASK 1 122.4865 69.379 122.6065 71.189 ;
      RECT MASK 1 122.9265 69.379 123.0465 71.189 ;
      RECT MASK 1 123.3665 69.379 123.4865 71.189 ;
      RECT MASK 1 123.8065 69.379 123.9265 71.189 ;
      RECT MASK 1 113.2465 70.8925 113.3665 71.649 ;
      RECT MASK 1 113.6865 70.8925 113.8065 71.649 ;
      RECT MASK 1 114.1265 70.8925 114.2465 71.649 ;
      RECT MASK 1 114.221 72.236 114.301 72.544 ;
      RECT MASK 1 114.387 72.236 114.467 72.544 ;
      RECT MASK 1 114.719 72.236 114.799 72.932 ;
      RECT MASK 1 115.051 72.236 115.131 72.932 ;
      RECT MASK 1 115.383 72.236 115.463 72.932 ;
      RECT MASK 1 115.715 72.236 115.795 72.932 ;
      RECT MASK 1 116.047 72.236 116.127 72.544 ;
      RECT MASK 1 116.379 72.236 116.459 72.544 ;
      RECT MASK 1 116.711 72.236 116.791 72.544 ;
      RECT MASK 1 117.043 72.236 117.123 72.544 ;
      RECT MASK 1 117.375 72.236 117.455 72.544 ;
      RECT MASK 1 117.707 72.236 117.787 72.544 ;
      RECT MASK 1 118.039 72.236 118.119 72.544 ;
      RECT MASK 1 118.371 72.236 118.451 72.544 ;
      RECT MASK 1 118.703 72.236 118.783 72.544 ;
      RECT MASK 1 119.035 72.236 119.115 72.544 ;
      RECT MASK 1 119.367 72.236 119.447 72.544 ;
      RECT MASK 1 119.699 72.236 119.779 72.544 ;
      RECT MASK 1 120.031 72.236 120.111 72.544 ;
      RECT MASK 1 120.363 72.236 120.443 72.544 ;
      RECT MASK 1 120.695 72.236 120.775 72.544 ;
      RECT MASK 1 121.027 72.236 121.107 72.544 ;
      RECT MASK 1 121.359 72.236 121.439 72.544 ;
      RECT MASK 1 121.691 72.236 121.771 72.544 ;
      RECT MASK 1 122.023 72.236 122.103 72.544 ;
      RECT MASK 1 122.355 72.236 122.435 72.544 ;
      RECT MASK 1 122.687 72.236 122.767 72.544 ;
      RECT MASK 1 123.019 72.236 123.099 72.544 ;
      RECT MASK 1 123.351 72.236 123.431 72.544 ;
      RECT MASK 1 123.683 72.236 123.763 72.544 ;
      RECT MASK 1 124.015 72.236 124.095 72.544 ;
      RECT MASK 1 124.181 72.236 124.261 72.544 ;
      RECT MASK 1 124.347 72.236 124.427 72.544 ;
      RECT MASK 1 124.513 72.236 124.593 72.544 ;
      RECT MASK 1 124.679 72.236 124.759 72.544 ;
      RECT MASK 1 124.845 72.236 124.925 72.544 ;
      RECT MASK 1 125.011 72.236 125.091 72.544 ;
      RECT MASK 1 125.177 72.236 125.257 72.544 ;
      RECT MASK 1 125.343 72.236 125.423 72.544 ;
      RECT MASK 1 125.675 72.236 125.755 72.544 ;
      RECT MASK 1 126.007 72.236 126.087 72.544 ;
      RECT MASK 1 126.339 72.236 126.419 72.544 ;
      RECT MASK 1 126.505 72.236 126.585 72.544 ;
      RECT MASK 1 126.671 72.236 126.751 72.544 ;
      RECT MASK 1 127.003 72.236 127.083 72.544 ;
      RECT MASK 1 127.169 72.236 127.249 72.544 ;
      RECT MASK 1 127.335 72.236 127.415 72.544 ;
      RECT MASK 1 127.667 72.236 127.747 72.544 ;
      RECT MASK 1 127.999 72.236 128.079 72.544 ;
      RECT MASK 1 128.331 72.236 128.411 72.544 ;
      RECT MASK 1 128.663 72.236 128.743 72.544 ;
      RECT MASK 1 113.869 72.26 113.989 77.818 ;
      RECT MASK 1 114.441 72.75 114.561 77.78 ;
      RECT MASK 1 116.095 73.196 116.175 80.458 ;
      RECT MASK 1 116.261 73.196 116.341 73.528 ;
      RECT MASK 1 116.593 73.196 116.673 73.528 ;
      RECT MASK 1 116.925 73.196 117.005 73.528 ;
      RECT MASK 1 117.257 73.196 117.337 73.528 ;
      RECT MASK 1 117.589 73.196 117.669 73.528 ;
      RECT MASK 1 117.921 73.196 118.001 73.528 ;
      RECT MASK 1 118.253 73.196 118.333 73.528 ;
      RECT MASK 1 118.585 73.196 118.665 73.528 ;
      RECT MASK 1 118.917 73.196 118.997 73.528 ;
      RECT MASK 1 119.249 73.196 119.329 73.528 ;
      RECT MASK 1 119.581 73.196 119.661 73.528 ;
      RECT MASK 1 119.913 73.196 119.993 73.528 ;
      RECT MASK 1 120.245 73.196 120.325 73.528 ;
      RECT MASK 1 120.577 73.196 120.657 73.528 ;
      RECT MASK 1 120.909 73.196 120.989 73.528 ;
      RECT MASK 1 121.241 73.196 121.321 73.528 ;
      RECT MASK 1 121.573 73.196 121.653 73.528 ;
      RECT MASK 1 121.905 73.196 121.985 73.528 ;
      RECT MASK 1 122.237 73.196 122.317 73.528 ;
      RECT MASK 1 122.569 73.196 122.649 73.528 ;
      RECT MASK 1 122.901 73.196 122.981 73.528 ;
      RECT MASK 1 123.233 73.196 123.313 73.528 ;
      RECT MASK 1 123.565 73.196 123.645 73.528 ;
      RECT MASK 1 123.897 73.196 123.977 73.528 ;
      RECT MASK 1 124.229 73.196 124.309 73.528 ;
      RECT MASK 1 124.395 73.196 124.475 73.528 ;
      RECT MASK 1 124.561 73.196 124.641 73.528 ;
      RECT MASK 1 124.893 73.196 124.973 73.528 ;
      RECT MASK 1 125.059 73.196 125.139 73.528 ;
      RECT MASK 1 125.225 73.196 125.305 73.528 ;
      RECT MASK 1 125.557 73.196 125.637 73.528 ;
      RECT MASK 1 125.889 73.196 125.969 73.528 ;
      RECT MASK 1 126.221 73.196 126.301 73.528 ;
      RECT MASK 1 126.387 73.196 126.467 80.4615 ;
      RECT MASK 1 116.261 73.958 116.341 74.242 ;
      RECT MASK 1 116.593 73.958 116.673 74.242 ;
      RECT MASK 1 116.925 73.958 117.005 74.242 ;
      RECT MASK 1 117.257 73.958 117.337 74.242 ;
      RECT MASK 1 117.589 73.958 117.669 74.242 ;
      RECT MASK 1 117.921 73.958 118.001 74.242 ;
      RECT MASK 1 118.253 73.958 118.333 74.242 ;
      RECT MASK 1 118.585 73.958 118.665 74.242 ;
      RECT MASK 1 118.917 73.958 118.997 74.242 ;
      RECT MASK 1 119.249 73.958 119.329 74.242 ;
      RECT MASK 1 119.581 73.958 119.661 74.242 ;
      RECT MASK 1 119.913 73.958 119.993 74.242 ;
      RECT MASK 1 120.245 73.958 120.325 74.242 ;
      RECT MASK 1 120.577 73.958 120.657 74.242 ;
      RECT MASK 1 120.909 73.958 120.989 74.242 ;
      RECT MASK 1 121.241 73.958 121.321 74.242 ;
      RECT MASK 1 121.573 73.958 121.653 74.242 ;
      RECT MASK 1 121.905 73.958 121.985 74.242 ;
      RECT MASK 1 122.237 73.958 122.317 74.242 ;
      RECT MASK 1 122.569 73.958 122.649 74.242 ;
      RECT MASK 1 122.901 73.958 122.981 74.242 ;
      RECT MASK 1 123.233 73.958 123.313 74.242 ;
      RECT MASK 1 123.565 73.958 123.645 74.242 ;
      RECT MASK 1 123.897 73.958 123.977 74.242 ;
      RECT MASK 1 124.229 73.958 124.309 74.242 ;
      RECT MASK 1 124.561 73.958 124.641 74.242 ;
      RECT MASK 1 124.893 73.958 124.973 74.242 ;
      RECT MASK 1 125.225 73.958 125.305 74.242 ;
      RECT MASK 1 125.557 73.958 125.637 74.242 ;
      RECT MASK 1 125.889 73.958 125.969 74.242 ;
      RECT MASK 1 126.221 73.958 126.301 74.242 ;
      RECT MASK 1 126.554 74.168 126.634 74.54 ;
      RECT MASK 1 116.261 74.736 116.341 75.022 ;
      RECT MASK 1 116.593 74.736 116.673 75.022 ;
      RECT MASK 1 116.925 74.736 117.005 75.022 ;
      RECT MASK 1 117.257 74.736 117.337 75.022 ;
      RECT MASK 1 117.589 74.736 117.669 75.022 ;
      RECT MASK 1 117.921 74.736 118.001 75.022 ;
      RECT MASK 1 118.253 74.736 118.333 75.022 ;
      RECT MASK 1 118.585 74.736 118.665 75.022 ;
      RECT MASK 1 118.917 74.736 118.997 75.022 ;
      RECT MASK 1 119.249 74.736 119.329 75.022 ;
      RECT MASK 1 119.581 74.736 119.661 75.022 ;
      RECT MASK 1 119.913 74.736 119.993 75.022 ;
      RECT MASK 1 120.245 74.736 120.325 75.022 ;
      RECT MASK 1 120.577 74.736 120.657 75.022 ;
      RECT MASK 1 120.909 74.736 120.989 75.022 ;
      RECT MASK 1 121.241 74.736 121.321 75.022 ;
      RECT MASK 1 121.573 74.736 121.653 75.022 ;
      RECT MASK 1 121.905 74.736 121.985 75.022 ;
      RECT MASK 1 122.237 74.736 122.317 75.022 ;
      RECT MASK 1 122.569 74.736 122.649 75.022 ;
      RECT MASK 1 122.901 74.736 122.981 75.022 ;
      RECT MASK 1 123.233 74.736 123.313 75.022 ;
      RECT MASK 1 123.565 74.736 123.645 75.022 ;
      RECT MASK 1 123.897 74.736 123.977 75.022 ;
      RECT MASK 1 124.229 74.736 124.309 75.022 ;
      RECT MASK 1 124.561 74.736 124.641 75.022 ;
      RECT MASK 1 124.893 74.736 124.973 75.022 ;
      RECT MASK 1 125.225 74.736 125.305 75.022 ;
      RECT MASK 1 125.557 74.736 125.637 75.022 ;
      RECT MASK 1 125.889 74.736 125.969 75.022 ;
      RECT MASK 1 126.221 74.736 126.301 75.022 ;
      RECT MASK 1 126.554 74.948 126.634 75.32 ;
      RECT MASK 1 116.261 75.507 116.341 75.802 ;
      RECT MASK 1 116.593 75.507 116.673 75.802 ;
      RECT MASK 1 116.925 75.507 117.005 75.802 ;
      RECT MASK 1 117.257 75.507 117.337 75.802 ;
      RECT MASK 1 117.589 75.507 117.669 75.802 ;
      RECT MASK 1 117.921 75.507 118.001 75.802 ;
      RECT MASK 1 118.253 75.507 118.333 75.802 ;
      RECT MASK 1 118.585 75.507 118.665 75.802 ;
      RECT MASK 1 118.917 75.507 118.997 75.802 ;
      RECT MASK 1 119.249 75.507 119.329 75.802 ;
      RECT MASK 1 119.581 75.507 119.661 75.802 ;
      RECT MASK 1 119.913 75.507 119.993 75.802 ;
      RECT MASK 1 120.245 75.507 120.325 75.802 ;
      RECT MASK 1 120.577 75.507 120.657 75.802 ;
      RECT MASK 1 120.909 75.507 120.989 75.802 ;
      RECT MASK 1 121.241 75.507 121.321 75.802 ;
      RECT MASK 1 121.573 75.507 121.653 75.802 ;
      RECT MASK 1 121.905 75.507 121.985 75.802 ;
      RECT MASK 1 122.237 75.507 122.317 75.802 ;
      RECT MASK 1 122.569 75.507 122.649 75.802 ;
      RECT MASK 1 122.901 75.507 122.981 75.802 ;
      RECT MASK 1 123.233 75.507 123.313 75.802 ;
      RECT MASK 1 123.565 75.507 123.645 75.802 ;
      RECT MASK 1 123.897 75.507 123.977 75.802 ;
      RECT MASK 1 124.229 75.507 124.309 75.802 ;
      RECT MASK 1 124.561 75.507 124.641 75.802 ;
      RECT MASK 1 124.893 75.507 124.973 75.802 ;
      RECT MASK 1 125.225 75.507 125.305 75.802 ;
      RECT MASK 1 125.557 75.507 125.637 75.802 ;
      RECT MASK 1 125.889 75.507 125.969 75.802 ;
      RECT MASK 1 126.221 75.507 126.301 75.802 ;
      RECT MASK 1 126.554 75.728 126.634 76.1 ;
      RECT MASK 1 116.261 76.297 116.341 76.589 ;
      RECT MASK 1 116.593 76.297 116.673 76.589 ;
      RECT MASK 1 116.925 76.297 117.005 76.589 ;
      RECT MASK 1 117.257 76.297 117.337 76.589 ;
      RECT MASK 1 117.589 76.297 117.669 76.589 ;
      RECT MASK 1 117.921 76.297 118.001 76.589 ;
      RECT MASK 1 118.253 76.297 118.333 76.589 ;
      RECT MASK 1 118.585 76.297 118.665 76.589 ;
      RECT MASK 1 118.917 76.297 118.997 76.589 ;
      RECT MASK 1 119.249 76.297 119.329 76.589 ;
      RECT MASK 1 119.581 76.297 119.661 76.589 ;
      RECT MASK 1 119.913 76.297 119.993 76.589 ;
      RECT MASK 1 120.245 76.297 120.325 76.589 ;
      RECT MASK 1 120.577 76.297 120.657 76.589 ;
      RECT MASK 1 120.909 76.297 120.989 76.589 ;
      RECT MASK 1 121.241 76.297 121.321 76.589 ;
      RECT MASK 1 121.573 76.297 121.653 76.589 ;
      RECT MASK 1 121.905 76.297 121.985 76.589 ;
      RECT MASK 1 122.237 76.297 122.317 76.589 ;
      RECT MASK 1 122.569 76.297 122.649 76.589 ;
      RECT MASK 1 122.901 76.297 122.981 76.589 ;
      RECT MASK 1 123.233 76.297 123.313 76.589 ;
      RECT MASK 1 123.565 76.297 123.645 76.589 ;
      RECT MASK 1 123.897 76.297 123.977 76.589 ;
      RECT MASK 1 124.229 76.297 124.309 76.589 ;
      RECT MASK 1 124.561 76.297 124.641 76.589 ;
      RECT MASK 1 124.893 76.297 124.973 76.589 ;
      RECT MASK 1 125.225 76.297 125.305 76.589 ;
      RECT MASK 1 125.557 76.297 125.637 76.589 ;
      RECT MASK 1 125.889 76.297 125.969 76.589 ;
      RECT MASK 1 126.221 76.297 126.301 76.589 ;
      RECT MASK 1 126.554 76.508 126.634 76.88 ;
      RECT MASK 1 116.261 77.081 116.341 77.366 ;
      RECT MASK 1 116.593 77.081 116.673 77.366 ;
      RECT MASK 1 116.925 77.081 117.005 77.366 ;
      RECT MASK 1 117.257 77.081 117.337 77.366 ;
      RECT MASK 1 117.589 77.081 117.669 77.366 ;
      RECT MASK 1 117.921 77.081 118.001 77.366 ;
      RECT MASK 1 118.253 77.081 118.333 77.366 ;
      RECT MASK 1 118.585 77.081 118.665 77.366 ;
      RECT MASK 1 118.917 77.081 118.997 77.366 ;
      RECT MASK 1 119.249 77.081 119.329 77.366 ;
      RECT MASK 1 119.581 77.081 119.661 77.366 ;
      RECT MASK 1 119.913 77.081 119.993 77.366 ;
      RECT MASK 1 120.245 77.081 120.325 77.366 ;
      RECT MASK 1 120.577 77.081 120.657 77.366 ;
      RECT MASK 1 120.909 77.081 120.989 77.366 ;
      RECT MASK 1 121.241 77.081 121.321 77.366 ;
      RECT MASK 1 121.573 77.081 121.653 77.366 ;
      RECT MASK 1 121.905 77.081 121.985 77.366 ;
      RECT MASK 1 122.237 77.081 122.317 77.366 ;
      RECT MASK 1 122.569 77.081 122.649 77.366 ;
      RECT MASK 1 122.901 77.081 122.981 77.366 ;
      RECT MASK 1 123.233 77.081 123.313 77.366 ;
      RECT MASK 1 123.565 77.081 123.645 77.366 ;
      RECT MASK 1 123.897 77.081 123.977 77.366 ;
      RECT MASK 1 124.229 77.081 124.309 77.366 ;
      RECT MASK 1 124.561 77.081 124.641 77.366 ;
      RECT MASK 1 124.893 77.081 124.973 77.366 ;
      RECT MASK 1 125.225 77.081 125.305 77.366 ;
      RECT MASK 1 125.557 77.081 125.637 77.366 ;
      RECT MASK 1 125.889 77.081 125.969 77.366 ;
      RECT MASK 1 126.221 77.081 126.301 77.366 ;
      RECT MASK 1 126.554 77.288 126.634 77.66 ;
      RECT MASK 1 2.005 77.486 2.085 77.818 ;
      RECT MASK 1 2.337 77.486 2.417 77.818 ;
      RECT MASK 1 2.669 77.486 2.749 77.818 ;
      RECT MASK 1 4.329 77.486 4.409 77.818 ;
      RECT MASK 1 4.661 77.486 4.741 77.818 ;
      RECT MASK 1 4.993 77.486 5.073 77.818 ;
      RECT MASK 1 5.325 77.486 5.405 77.818 ;
      RECT MASK 1 5.657 77.486 5.737 77.818 ;
      RECT MASK 1 5.989 77.486 6.069 77.818 ;
      RECT MASK 1 6.321 77.486 6.401 77.818 ;
      RECT MASK 1 6.653 77.486 6.733 77.818 ;
      RECT MASK 1 6.985 77.486 7.065 77.818 ;
      RECT MASK 1 7.317 77.486 7.397 77.818 ;
      RECT MASK 1 7.649 77.486 7.729 77.818 ;
      RECT MASK 1 7.981 77.486 8.061 77.818 ;
      RECT MASK 1 8.313 77.486 8.393 77.818 ;
      RECT MASK 1 8.645 77.486 8.725 77.818 ;
      RECT MASK 1 8.977 77.486 9.057 77.818 ;
      RECT MASK 1 9.309 77.486 9.389 77.818 ;
      RECT MASK 1 9.641 77.486 9.721 77.818 ;
      RECT MASK 1 9.973 77.486 10.053 77.818 ;
      RECT MASK 1 10.305 77.486 10.385 77.818 ;
      RECT MASK 1 10.637 77.486 10.717 77.818 ;
      RECT MASK 1 10.969 77.486 11.049 77.818 ;
      RECT MASK 1 11.301 77.486 11.381 77.818 ;
      RECT MASK 1 11.633 77.486 11.713 77.818 ;
      RECT MASK 1 11.965 77.486 12.045 77.818 ;
      RECT MASK 1 12.297 77.486 12.377 77.818 ;
      RECT MASK 1 12.629 77.486 12.709 77.818 ;
      RECT MASK 1 12.961 77.486 13.041 77.818 ;
      RECT MASK 1 13.293 77.486 13.373 77.818 ;
      RECT MASK 1 13.625 77.486 13.705 77.818 ;
      RECT MASK 1 13.957 77.486 14.037 77.818 ;
      RECT MASK 1 14.289 77.486 14.369 77.818 ;
      RECT MASK 1 14.621 77.486 14.701 77.818 ;
      RECT MASK 1 14.953 77.486 15.033 77.818 ;
      RECT MASK 1 15.285 77.486 15.365 77.818 ;
      RECT MASK 1 15.617 77.486 15.697 77.818 ;
      RECT MASK 1 15.949 77.486 16.029 77.818 ;
      RECT MASK 1 16.281 77.486 16.361 77.818 ;
      RECT MASK 1 16.613 77.486 16.693 77.818 ;
      RECT MASK 1 16.945 77.486 17.025 77.818 ;
      RECT MASK 1 17.277 77.486 17.357 77.818 ;
      RECT MASK 1 17.609 77.486 17.689 77.818 ;
      RECT MASK 1 17.941 77.486 18.021 77.818 ;
      RECT MASK 1 18.273 77.486 18.353 77.818 ;
      RECT MASK 1 18.605 77.486 18.685 77.818 ;
      RECT MASK 1 18.937 77.486 19.017 77.818 ;
      RECT MASK 1 19.269 77.486 19.349 77.818 ;
      RECT MASK 1 19.601 77.486 19.681 77.818 ;
      RECT MASK 1 19.933 77.486 20.013 77.818 ;
      RECT MASK 1 20.265 77.486 20.345 77.818 ;
      RECT MASK 1 20.597 77.486 20.677 77.818 ;
      RECT MASK 1 20.929 77.486 21.009 77.818 ;
      RECT MASK 1 21.261 77.486 21.341 77.818 ;
      RECT MASK 1 21.593 77.486 21.673 77.818 ;
      RECT MASK 1 21.925 77.486 22.005 77.818 ;
      RECT MASK 1 22.257 77.486 22.337 77.818 ;
      RECT MASK 1 22.589 77.486 22.669 77.818 ;
      RECT MASK 1 22.921 77.486 23.001 77.818 ;
      RECT MASK 1 23.253 77.486 23.333 77.818 ;
      RECT MASK 1 23.585 77.486 23.665 77.818 ;
      RECT MASK 1 23.917 77.486 23.997 77.818 ;
      RECT MASK 1 24.249 77.486 24.329 77.818 ;
      RECT MASK 1 24.581 77.486 24.661 77.818 ;
      RECT MASK 1 24.913 77.486 24.993 77.818 ;
      RECT MASK 1 25.245 77.486 25.325 77.818 ;
      RECT MASK 1 25.577 77.486 25.657 77.818 ;
      RECT MASK 1 25.909 77.486 25.989 77.818 ;
      RECT MASK 1 26.241 77.486 26.321 77.818 ;
      RECT MASK 1 26.573 77.486 26.653 77.818 ;
      RECT MASK 1 26.905 77.486 26.985 77.818 ;
      RECT MASK 1 27.237 77.486 27.317 77.818 ;
      RECT MASK 1 27.569 77.486 27.649 77.818 ;
      RECT MASK 1 27.901 77.486 27.981 77.818 ;
      RECT MASK 1 28.233 77.486 28.313 77.818 ;
      RECT MASK 1 28.565 77.486 28.645 77.818 ;
      RECT MASK 1 28.897 77.486 28.977 77.818 ;
      RECT MASK 1 29.229 77.486 29.309 77.818 ;
      RECT MASK 1 29.561 77.486 29.641 77.818 ;
      RECT MASK 1 29.893 77.486 29.973 77.818 ;
      RECT MASK 1 30.225 77.486 30.305 77.818 ;
      RECT MASK 1 30.557 77.486 30.637 77.818 ;
      RECT MASK 1 30.889 77.486 30.969 77.818 ;
      RECT MASK 1 31.221 77.486 31.301 77.818 ;
      RECT MASK 1 31.553 77.486 31.633 77.818 ;
      RECT MASK 1 31.885 77.486 31.965 77.818 ;
      RECT MASK 1 32.217 77.486 32.297 77.818 ;
      RECT MASK 1 32.549 77.486 32.629 77.818 ;
      RECT MASK 1 32.881 77.486 32.961 77.818 ;
      RECT MASK 1 33.213 77.486 33.293 77.818 ;
      RECT MASK 1 33.545 77.486 33.625 77.818 ;
      RECT MASK 1 33.877 77.486 33.957 77.818 ;
      RECT MASK 1 34.209 77.486 34.289 77.818 ;
      RECT MASK 1 34.541 77.486 34.621 77.818 ;
      RECT MASK 1 34.873 77.486 34.953 77.818 ;
      RECT MASK 1 35.205 77.486 35.285 77.818 ;
      RECT MASK 1 35.537 77.486 35.617 77.818 ;
      RECT MASK 1 35.869 77.486 35.949 77.818 ;
      RECT MASK 1 36.201 77.486 36.281 77.818 ;
      RECT MASK 1 36.533 77.486 36.613 77.818 ;
      RECT MASK 1 36.865 77.486 36.945 77.818 ;
      RECT MASK 1 37.197 77.486 37.277 77.818 ;
      RECT MASK 1 37.529 77.486 37.609 77.818 ;
      RECT MASK 1 37.861 77.486 37.941 77.818 ;
      RECT MASK 1 38.193 77.486 38.273 77.818 ;
      RECT MASK 1 38.525 77.486 38.605 77.818 ;
      RECT MASK 1 38.857 77.486 38.937 77.818 ;
      RECT MASK 1 39.189 77.486 39.269 77.818 ;
      RECT MASK 1 39.521 77.486 39.601 77.818 ;
      RECT MASK 1 39.853 77.486 39.933 77.818 ;
      RECT MASK 1 40.185 77.486 40.265 77.818 ;
      RECT MASK 1 40.517 77.486 40.597 77.818 ;
      RECT MASK 1 40.849 77.486 40.929 77.818 ;
      RECT MASK 1 41.181 77.486 41.261 77.818 ;
      RECT MASK 1 41.513 77.486 41.593 77.818 ;
      RECT MASK 1 41.845 77.486 41.925 77.818 ;
      RECT MASK 1 42.177 77.486 42.257 77.818 ;
      RECT MASK 1 42.509 77.486 42.589 77.818 ;
      RECT MASK 1 42.841 77.486 42.921 77.818 ;
      RECT MASK 1 43.173 77.486 43.253 77.818 ;
      RECT MASK 1 43.505 77.486 43.585 77.818 ;
      RECT MASK 1 43.837 77.486 43.917 77.818 ;
      RECT MASK 1 44.169 77.486 44.249 77.818 ;
      RECT MASK 1 44.501 77.486 44.581 77.818 ;
      RECT MASK 1 44.833 77.486 44.913 77.818 ;
      RECT MASK 1 45.165 77.486 45.245 77.818 ;
      RECT MASK 1 45.497 77.486 45.577 77.818 ;
      RECT MASK 1 45.829 77.486 45.909 77.818 ;
      RECT MASK 1 46.161 77.486 46.241 77.818 ;
      RECT MASK 1 46.493 77.486 46.573 77.818 ;
      RECT MASK 1 46.825 77.486 46.905 77.818 ;
      RECT MASK 1 47.157 77.486 47.237 77.818 ;
      RECT MASK 1 47.489 77.486 47.569 77.818 ;
      RECT MASK 1 47.821 77.486 47.901 77.818 ;
      RECT MASK 1 48.153 77.486 48.233 77.818 ;
      RECT MASK 1 48.485 77.486 48.565 77.818 ;
      RECT MASK 1 48.817 77.486 48.897 77.818 ;
      RECT MASK 1 49.149 77.486 49.229 77.818 ;
      RECT MASK 1 49.481 77.486 49.561 77.818 ;
      RECT MASK 1 49.813 77.486 49.893 77.818 ;
      RECT MASK 1 50.145 77.486 50.225 77.818 ;
      RECT MASK 1 50.477 77.486 50.557 77.818 ;
      RECT MASK 1 50.809 77.486 50.889 77.818 ;
      RECT MASK 1 51.141 77.486 51.221 77.818 ;
      RECT MASK 1 51.473 77.486 51.553 77.818 ;
      RECT MASK 1 51.805 77.486 51.885 77.818 ;
      RECT MASK 1 52.137 77.486 52.217 77.818 ;
      RECT MASK 1 52.469 77.486 52.549 77.818 ;
      RECT MASK 1 52.801 77.486 52.881 77.818 ;
      RECT MASK 1 53.133 77.486 53.213 77.818 ;
      RECT MASK 1 53.465 77.486 53.545 77.818 ;
      RECT MASK 1 53.797 77.486 53.877 77.818 ;
      RECT MASK 1 54.129 77.486 54.209 77.818 ;
      RECT MASK 1 54.461 77.486 54.541 77.818 ;
      RECT MASK 1 54.793 77.486 54.873 77.818 ;
      RECT MASK 1 55.125 77.486 55.205 77.818 ;
      RECT MASK 1 55.457 77.486 55.537 77.818 ;
      RECT MASK 1 55.789 77.486 55.869 77.818 ;
      RECT MASK 1 56.121 77.486 56.201 77.818 ;
      RECT MASK 1 56.453 77.486 56.533 77.818 ;
      RECT MASK 1 56.785 77.486 56.865 77.818 ;
      RECT MASK 1 57.117 77.486 57.197 77.818 ;
      RECT MASK 1 57.449 77.486 57.529 77.818 ;
      RECT MASK 1 57.781 77.486 57.861 77.818 ;
      RECT MASK 1 58.113 77.486 58.193 77.818 ;
      RECT MASK 1 58.445 77.486 58.525 77.818 ;
      RECT MASK 1 58.777 77.486 58.857 77.818 ;
      RECT MASK 1 59.109 77.486 59.189 77.818 ;
      RECT MASK 1 59.441 77.486 59.521 77.818 ;
      RECT MASK 1 59.773 77.486 59.853 77.818 ;
      RECT MASK 1 60.105 77.486 60.185 77.818 ;
      RECT MASK 1 60.437 77.486 60.517 77.818 ;
      RECT MASK 1 60.769 77.486 60.849 77.818 ;
      RECT MASK 1 61.101 77.486 61.181 77.818 ;
      RECT MASK 1 61.433 77.486 61.513 77.818 ;
      RECT MASK 1 61.765 77.486 61.845 77.818 ;
      RECT MASK 1 62.097 77.486 62.177 77.818 ;
      RECT MASK 1 62.429 77.486 62.509 77.818 ;
      RECT MASK 1 62.761 77.486 62.841 77.818 ;
      RECT MASK 1 63.093 77.486 63.173 77.818 ;
      RECT MASK 1 63.425 77.486 63.505 77.818 ;
      RECT MASK 1 63.757 77.486 63.837 77.818 ;
      RECT MASK 1 64.089 77.486 64.169 77.818 ;
      RECT MASK 1 64.421 77.486 64.501 77.818 ;
      RECT MASK 1 64.753 77.486 64.833 77.818 ;
      RECT MASK 1 65.085 77.486 65.165 77.818 ;
      RECT MASK 1 65.417 77.486 65.497 77.818 ;
      RECT MASK 1 65.749 77.486 65.829 77.818 ;
      RECT MASK 1 66.081 77.486 66.161 77.818 ;
      RECT MASK 1 66.413 77.486 66.493 77.818 ;
      RECT MASK 1 66.745 77.486 66.825 77.818 ;
      RECT MASK 1 67.077 77.486 67.157 77.818 ;
      RECT MASK 1 67.409 77.486 67.489 77.818 ;
      RECT MASK 1 67.741 77.486 67.821 77.818 ;
      RECT MASK 1 68.073 77.486 68.153 77.818 ;
      RECT MASK 1 68.405 77.486 68.485 77.818 ;
      RECT MASK 1 68.737 77.486 68.817 77.818 ;
      RECT MASK 1 69.069 77.486 69.149 77.818 ;
      RECT MASK 1 69.401 77.486 69.481 77.818 ;
      RECT MASK 1 69.733 77.486 69.813 77.818 ;
      RECT MASK 1 70.065 77.486 70.145 77.818 ;
      RECT MASK 1 70.397 77.486 70.477 77.818 ;
      RECT MASK 1 70.729 77.486 70.809 77.818 ;
      RECT MASK 1 71.061 77.486 71.141 77.818 ;
      RECT MASK 1 71.393 77.486 71.473 77.818 ;
      RECT MASK 1 71.725 77.486 71.805 77.818 ;
      RECT MASK 1 72.057 77.486 72.137 77.818 ;
      RECT MASK 1 72.389 77.486 72.469 77.818 ;
      RECT MASK 1 72.721 77.486 72.801 77.818 ;
      RECT MASK 1 73.053 77.486 73.133 77.818 ;
      RECT MASK 1 73.385 77.486 73.465 77.818 ;
      RECT MASK 1 73.717 77.486 73.797 77.818 ;
      RECT MASK 1 74.049 77.486 74.129 77.818 ;
      RECT MASK 1 74.381 77.486 74.461 77.818 ;
      RECT MASK 1 74.713 77.486 74.793 77.818 ;
      RECT MASK 1 75.045 77.486 75.125 77.818 ;
      RECT MASK 1 75.377 77.486 75.457 77.818 ;
      RECT MASK 1 75.709 77.486 75.789 77.818 ;
      RECT MASK 1 76.041 77.486 76.121 77.818 ;
      RECT MASK 1 76.373 77.486 76.453 77.818 ;
      RECT MASK 1 76.705 77.486 76.785 77.818 ;
      RECT MASK 1 77.037 77.486 77.117 77.818 ;
      RECT MASK 1 77.369 77.486 77.449 77.818 ;
      RECT MASK 1 77.701 77.486 77.781 77.818 ;
      RECT MASK 1 78.033 77.486 78.113 77.818 ;
      RECT MASK 1 78.365 77.486 78.445 77.818 ;
      RECT MASK 1 78.697 77.486 78.777 77.818 ;
      RECT MASK 1 79.029 77.486 79.109 77.818 ;
      RECT MASK 1 79.361 77.486 79.441 77.818 ;
      RECT MASK 1 79.693 77.486 79.773 77.818 ;
      RECT MASK 1 80.025 77.486 80.105 77.818 ;
      RECT MASK 1 80.357 77.486 80.437 77.818 ;
      RECT MASK 1 80.689 77.486 80.769 77.818 ;
      RECT MASK 1 81.021 77.486 81.101 77.818 ;
      RECT MASK 1 81.353 77.486 81.433 77.818 ;
      RECT MASK 1 81.685 77.486 81.765 77.818 ;
      RECT MASK 1 82.017 77.486 82.097 77.818 ;
      RECT MASK 1 82.349 77.486 82.429 77.818 ;
      RECT MASK 1 82.681 77.486 82.761 77.818 ;
      RECT MASK 1 83.013 77.486 83.093 77.818 ;
      RECT MASK 1 83.345 77.486 83.425 77.818 ;
      RECT MASK 1 83.677 77.486 83.757 77.818 ;
      RECT MASK 1 84.009 77.486 84.089 77.818 ;
      RECT MASK 1 84.341 77.486 84.421 77.818 ;
      RECT MASK 1 84.673 77.486 84.753 77.818 ;
      RECT MASK 1 85.005 77.486 85.085 77.818 ;
      RECT MASK 1 85.337 77.486 85.417 77.818 ;
      RECT MASK 1 85.669 77.486 85.749 77.818 ;
      RECT MASK 1 86.001 77.486 86.081 77.818 ;
      RECT MASK 1 86.333 77.486 86.413 77.818 ;
      RECT MASK 1 86.665 77.486 86.745 77.818 ;
      RECT MASK 1 86.997 77.486 87.077 77.818 ;
      RECT MASK 1 87.329 77.486 87.409 77.818 ;
      RECT MASK 1 87.661 77.486 87.741 77.818 ;
      RECT MASK 1 87.993 77.486 88.073 77.818 ;
      RECT MASK 1 88.325 77.486 88.405 77.818 ;
      RECT MASK 1 88.657 77.486 88.737 77.818 ;
      RECT MASK 1 88.989 77.486 89.069 77.818 ;
      RECT MASK 1 89.321 77.486 89.401 77.818 ;
      RECT MASK 1 89.653 77.486 89.733 77.818 ;
      RECT MASK 1 89.985 77.486 90.065 77.818 ;
      RECT MASK 1 90.317 77.486 90.397 77.818 ;
      RECT MASK 1 90.649 77.486 90.729 77.818 ;
      RECT MASK 1 90.981 77.486 91.061 77.818 ;
      RECT MASK 1 91.313 77.486 91.393 77.818 ;
      RECT MASK 1 91.645 77.486 91.725 77.818 ;
      RECT MASK 1 91.977 77.486 92.057 77.818 ;
      RECT MASK 1 92.309 77.486 92.389 77.818 ;
      RECT MASK 1 92.641 77.486 92.721 77.818 ;
      RECT MASK 1 92.973 77.486 93.053 77.818 ;
      RECT MASK 1 93.305 77.486 93.385 77.818 ;
      RECT MASK 1 93.637 77.486 93.717 77.818 ;
      RECT MASK 1 93.969 77.486 94.049 77.818 ;
      RECT MASK 1 94.301 77.486 94.381 77.818 ;
      RECT MASK 1 94.633 77.486 94.713 77.818 ;
      RECT MASK 1 94.965 77.486 95.045 77.818 ;
      RECT MASK 1 95.297 77.486 95.377 77.818 ;
      RECT MASK 1 95.629 77.486 95.709 77.818 ;
      RECT MASK 1 95.961 77.486 96.041 77.818 ;
      RECT MASK 1 96.293 77.486 96.373 77.818 ;
      RECT MASK 1 96.625 77.486 96.705 77.818 ;
      RECT MASK 1 96.957 77.486 97.037 77.818 ;
      RECT MASK 1 97.289 77.486 97.369 77.818 ;
      RECT MASK 1 97.621 77.486 97.701 77.818 ;
      RECT MASK 1 97.953 77.486 98.033 77.818 ;
      RECT MASK 1 98.285 77.486 98.365 77.818 ;
      RECT MASK 1 98.617 77.486 98.697 77.818 ;
      RECT MASK 1 98.949 77.486 99.029 77.818 ;
      RECT MASK 1 99.281 77.486 99.361 77.818 ;
      RECT MASK 1 99.613 77.486 99.693 77.818 ;
      RECT MASK 1 99.945 77.486 100.025 77.818 ;
      RECT MASK 1 100.277 77.486 100.357 77.818 ;
      RECT MASK 1 100.609 77.486 100.689 77.818 ;
      RECT MASK 1 100.941 77.486 101.021 77.818 ;
      RECT MASK 1 101.273 77.486 101.353 77.818 ;
      RECT MASK 1 101.605 77.486 101.685 77.818 ;
      RECT MASK 1 101.937 77.486 102.017 77.818 ;
      RECT MASK 1 102.269 77.486 102.349 77.818 ;
      RECT MASK 1 102.601 77.486 102.681 77.818 ;
      RECT MASK 1 102.933 77.486 103.013 77.818 ;
      RECT MASK 1 103.265 77.486 103.345 77.818 ;
      RECT MASK 1 103.597 77.486 103.677 77.818 ;
      RECT MASK 1 103.929 77.486 104.009 77.818 ;
      RECT MASK 1 104.261 77.486 104.341 77.818 ;
      RECT MASK 1 104.593 77.486 104.673 77.818 ;
      RECT MASK 1 104.925 77.486 105.005 77.818 ;
      RECT MASK 1 105.257 77.486 105.337 77.818 ;
      RECT MASK 1 105.589 77.486 105.669 77.818 ;
      RECT MASK 1 105.921 77.486 106.001 77.818 ;
      RECT MASK 1 106.253 77.486 106.333 77.818 ;
      RECT MASK 1 106.585 77.486 106.665 77.818 ;
      RECT MASK 1 106.917 77.486 106.997 77.818 ;
      RECT MASK 1 107.249 77.486 107.329 77.818 ;
      RECT MASK 1 107.581 77.486 107.661 77.818 ;
      RECT MASK 1 107.913 77.486 107.993 77.818 ;
      RECT MASK 1 108.245 77.486 108.325 77.818 ;
      RECT MASK 1 108.577 77.486 108.657 77.818 ;
      RECT MASK 1 108.909 77.486 108.989 77.818 ;
      RECT MASK 1 109.241 77.486 109.321 77.818 ;
      RECT MASK 1 109.573 77.486 109.653 77.818 ;
      RECT MASK 1 109.905 77.486 109.985 77.818 ;
      RECT MASK 1 110.237 77.486 110.317 77.818 ;
      RECT MASK 1 110.569 77.486 110.649 77.818 ;
      RECT MASK 1 110.901 77.486 110.981 77.818 ;
      RECT MASK 1 112.229 77.486 112.309 77.818 ;
      RECT MASK 1 112.561 77.486 112.641 77.818 ;
      RECT MASK 1 112.893 77.486 112.973 77.818 ;
      RECT MASK 1 113.225 77.486 113.305 77.818 ;
      RECT MASK 1 113.557 77.486 113.637 77.818 ;
      RECT MASK 1 116.261 77.855 116.341 78.157 ;
      RECT MASK 1 116.593 77.855 116.673 78.157 ;
      RECT MASK 1 116.925 77.855 117.005 78.157 ;
      RECT MASK 1 117.257 77.855 117.337 78.157 ;
      RECT MASK 1 117.589 77.855 117.669 78.157 ;
      RECT MASK 1 117.921 77.855 118.001 78.157 ;
      RECT MASK 1 118.253 77.855 118.333 78.157 ;
      RECT MASK 1 118.585 77.855 118.665 78.157 ;
      RECT MASK 1 118.917 77.855 118.997 78.157 ;
      RECT MASK 1 119.249 77.855 119.329 78.157 ;
      RECT MASK 1 119.581 77.855 119.661 78.157 ;
      RECT MASK 1 119.913 77.855 119.993 78.157 ;
      RECT MASK 1 120.245 77.855 120.325 78.157 ;
      RECT MASK 1 120.577 77.855 120.657 78.157 ;
      RECT MASK 1 120.909 77.855 120.989 78.157 ;
      RECT MASK 1 121.241 77.855 121.321 78.157 ;
      RECT MASK 1 121.573 77.855 121.653 78.157 ;
      RECT MASK 1 121.905 77.855 121.985 78.157 ;
      RECT MASK 1 122.237 77.855 122.317 78.157 ;
      RECT MASK 1 122.569 77.855 122.649 78.157 ;
      RECT MASK 1 122.901 77.855 122.981 78.157 ;
      RECT MASK 1 123.233 77.855 123.313 78.157 ;
      RECT MASK 1 123.565 77.855 123.645 78.157 ;
      RECT MASK 1 123.897 77.855 123.977 78.157 ;
      RECT MASK 1 124.229 77.855 124.309 78.157 ;
      RECT MASK 1 124.561 77.855 124.641 78.157 ;
      RECT MASK 1 124.893 77.855 124.973 78.157 ;
      RECT MASK 1 125.225 77.855 125.305 78.157 ;
      RECT MASK 1 125.557 77.855 125.637 78.157 ;
      RECT MASK 1 125.889 77.855 125.969 78.157 ;
      RECT MASK 1 126.221 77.855 126.301 78.157 ;
      RECT MASK 1 6.329 77.9995 6.389 80.28 ;
      RECT MASK 1 77.965 78.005 78.025 80.28 ;
      RECT MASK 1 11.785 78.0125 11.845 80.28 ;
      RECT MASK 1 63.423 78.0125 63.483 80.245 ;
      RECT MASK 1 64.729 78.0125 64.789 80.28 ;
      RECT MASK 1 89.895 78.0165 89.955 80.28 ;
      RECT MASK 1 91.201 78.0165 91.261 80.28 ;
      RECT MASK 1 36.951 78.02 37.011 80.28 ;
      RECT MASK 1 38.257 78.02 38.317 80.28 ;
      RECT MASK 1 10.479 78.022 10.539 80.28 ;
      RECT MASK 1 43.569 78.022 43.629 80.28 ;
      RECT MASK 1 44.875 78.022 44.935 80.28 ;
      RECT MASK 1 96.513 78.022 96.573 80.28 ;
      RECT MASK 1 97.819 78.022 97.879 80.28 ;
      RECT MASK 1 56.805 78.023 56.865 80.28 ;
      RECT MASK 1 58.111 78.023 58.171 80.28 ;
      RECT MASK 1 83.277 78.0235 83.337 80.28 ;
      RECT MASK 1 84.583 78.0235 84.643 80.28 ;
      RECT MASK 1 18.403 78.024 18.463 80.28 ;
      RECT MASK 1 30.333 78.0255 30.393 80.28 ;
      RECT MASK 1 31.639 78.0255 31.699 80.28 ;
      RECT MASK 1 76.659 78.0255 76.719 80.28 ;
      RECT MASK 1 50.187 78.0275 50.247 80.28 ;
      RECT MASK 1 51.493 78.0275 51.553 80.28 ;
      RECT MASK 1 103.131 78.0275 103.191 80.28 ;
      RECT MASK 1 104.437 78.0275 104.497 80.28 ;
      RECT MASK 1 6.993 78.03 7.053 78.3 ;
      RECT MASK 1 7.325 78.03 7.385 78.3 ;
      RECT MASK 1 7.657 78.03 7.717 78.3 ;
      RECT MASK 1 8.155 78.03 8.215 78.3 ;
      RECT MASK 1 8.487 78.03 8.547 78.3 ;
      RECT MASK 1 8.819 78.03 8.879 78.3 ;
      RECT MASK 1 9.317 78.03 9.377 78.3 ;
      RECT MASK 1 9.649 78.03 9.709 78.3 ;
      RECT MASK 1 9.981 78.03 10.041 78.3 ;
      RECT MASK 1 12.449 78.03 12.509 78.3 ;
      RECT MASK 1 12.781 78.03 12.841 78.3 ;
      RECT MASK 1 13.113 78.03 13.173 78.3 ;
      RECT MASK 1 13.611 78.03 13.671 78.3 ;
      RECT MASK 1 13.943 78.03 14.003 78.3 ;
      RECT MASK 1 14.275 78.03 14.335 78.3 ;
      RECT MASK 1 14.773 78.03 14.833 78.3 ;
      RECT MASK 1 15.105 78.03 15.165 78.3 ;
      RECT MASK 1 15.437 78.03 15.497 78.3 ;
      RECT MASK 1 15.935 78.03 15.995 78.3 ;
      RECT MASK 1 16.267 78.03 16.327 78.3 ;
      RECT MASK 1 16.599 78.03 16.659 78.3 ;
      RECT MASK 1 17.667 78.03 17.727 80.25 ;
      RECT MASK 1 17.999 78.03 18.059 80.25 ;
      RECT MASK 1 19.067 78.03 19.127 78.3 ;
      RECT MASK 1 19.399 78.03 19.459 78.3 ;
      RECT MASK 1 19.731 78.03 19.791 78.3 ;
      RECT MASK 1 20.229 78.03 20.289 78.3 ;
      RECT MASK 1 20.561 78.03 20.621 78.3 ;
      RECT MASK 1 20.893 78.03 20.953 78.3 ;
      RECT MASK 1 21.391 78.03 21.451 78.3 ;
      RECT MASK 1 21.723 78.03 21.783 78.3 ;
      RECT MASK 1 22.055 78.03 22.115 78.3 ;
      RECT MASK 1 22.553 78.03 22.613 78.3 ;
      RECT MASK 1 22.885 78.03 22.945 78.3 ;
      RECT MASK 1 23.217 78.03 23.277 78.3 ;
      RECT MASK 1 25.685 78.03 25.745 78.3 ;
      RECT MASK 1 26.017 78.03 26.077 78.3 ;
      RECT MASK 1 26.349 78.03 26.409 78.3 ;
      RECT MASK 1 26.847 78.03 26.907 78.3 ;
      RECT MASK 1 27.179 78.03 27.239 78.3 ;
      RECT MASK 1 27.511 78.03 27.571 78.3 ;
      RECT MASK 1 28.009 78.03 28.069 78.3 ;
      RECT MASK 1 28.341 78.03 28.401 78.3 ;
      RECT MASK 1 28.673 78.03 28.733 78.3 ;
      RECT MASK 1 29.171 78.03 29.231 78.3 ;
      RECT MASK 1 29.503 78.03 29.563 78.3 ;
      RECT MASK 1 29.835 78.03 29.895 78.3 ;
      RECT MASK 1 32.303 78.03 32.363 78.3 ;
      RECT MASK 1 32.635 78.03 32.695 78.3 ;
      RECT MASK 1 32.967 78.03 33.027 78.3 ;
      RECT MASK 1 33.465 78.03 33.525 78.3 ;
      RECT MASK 1 33.797 78.03 33.857 78.3 ;
      RECT MASK 1 34.129 78.03 34.189 78.3 ;
      RECT MASK 1 34.627 78.03 34.687 78.3 ;
      RECT MASK 1 34.959 78.03 35.019 78.3 ;
      RECT MASK 1 35.291 78.03 35.351 78.3 ;
      RECT MASK 1 35.789 78.03 35.849 78.3 ;
      RECT MASK 1 36.121 78.03 36.181 78.3 ;
      RECT MASK 1 36.453 78.03 36.513 78.3 ;
      RECT MASK 1 38.921 78.03 38.981 78.3 ;
      RECT MASK 1 39.253 78.03 39.313 78.3 ;
      RECT MASK 1 39.585 78.03 39.645 78.3 ;
      RECT MASK 1 40.083 78.03 40.143 78.3 ;
      RECT MASK 1 40.415 78.03 40.475 78.3 ;
      RECT MASK 1 40.747 78.03 40.807 78.3 ;
      RECT MASK 1 41.245 78.03 41.305 78.3 ;
      RECT MASK 1 41.577 78.03 41.637 78.3 ;
      RECT MASK 1 41.909 78.03 41.969 78.3 ;
      RECT MASK 1 42.407 78.03 42.467 78.3 ;
      RECT MASK 1 42.739 78.03 42.799 78.3 ;
      RECT MASK 1 43.071 78.03 43.131 78.3 ;
      RECT MASK 1 45.539 78.03 45.599 78.3 ;
      RECT MASK 1 45.871 78.03 45.931 78.3 ;
      RECT MASK 1 46.203 78.03 46.263 78.3 ;
      RECT MASK 1 46.701 78.03 46.761 78.3 ;
      RECT MASK 1 47.033 78.03 47.093 78.3 ;
      RECT MASK 1 47.365 78.03 47.425 78.3 ;
      RECT MASK 1 47.863 78.03 47.923 78.3 ;
      RECT MASK 1 48.195 78.03 48.255 78.3 ;
      RECT MASK 1 48.527 78.03 48.587 78.3 ;
      RECT MASK 1 49.025 78.03 49.085 78.3 ;
      RECT MASK 1 49.357 78.03 49.417 78.3 ;
      RECT MASK 1 49.689 78.03 49.749 78.3 ;
      RECT MASK 1 52.157 78.03 52.217 78.3 ;
      RECT MASK 1 52.489 78.03 52.549 78.3 ;
      RECT MASK 1 52.821 78.03 52.881 78.3 ;
      RECT MASK 1 53.319 78.03 53.379 78.3 ;
      RECT MASK 1 53.651 78.03 53.711 78.3 ;
      RECT MASK 1 53.983 78.03 54.043 78.3 ;
      RECT MASK 1 54.481 78.03 54.541 78.3 ;
      RECT MASK 1 54.813 78.03 54.873 78.3 ;
      RECT MASK 1 55.145 78.03 55.205 78.3 ;
      RECT MASK 1 55.643 78.03 55.703 78.3 ;
      RECT MASK 1 55.975 78.03 56.035 78.3 ;
      RECT MASK 1 56.307 78.03 56.367 78.3 ;
      RECT MASK 1 58.775 78.03 58.835 78.3 ;
      RECT MASK 1 59.107 78.03 59.167 78.3 ;
      RECT MASK 1 59.439 78.03 59.499 78.3 ;
      RECT MASK 1 59.937 78.03 59.997 78.3 ;
      RECT MASK 1 60.269 78.03 60.329 78.3 ;
      RECT MASK 1 60.601 78.03 60.661 78.3 ;
      RECT MASK 1 61.099 78.03 61.159 78.3 ;
      RECT MASK 1 61.431 78.03 61.491 78.3 ;
      RECT MASK 1 61.763 78.03 61.823 78.3 ;
      RECT MASK 1 62.261 78.03 62.321 78.3 ;
      RECT MASK 1 62.593 78.03 62.653 78.3 ;
      RECT MASK 1 62.925 78.03 62.985 78.3 ;
      RECT MASK 1 65.393 78.03 65.453 78.3 ;
      RECT MASK 1 65.725 78.03 65.785 78.3 ;
      RECT MASK 1 66.057 78.03 66.117 78.3 ;
      RECT MASK 1 66.555 78.03 66.615 78.3 ;
      RECT MASK 1 66.887 78.03 66.947 78.3 ;
      RECT MASK 1 67.219 78.03 67.279 78.3 ;
      RECT MASK 1 67.717 78.03 67.777 78.3 ;
      RECT MASK 1 68.049 78.03 68.109 78.3 ;
      RECT MASK 1 68.381 78.03 68.441 78.3 ;
      RECT MASK 1 68.879 78.03 68.939 78.3 ;
      RECT MASK 1 69.211 78.03 69.271 78.3 ;
      RECT MASK 1 69.543 78.03 69.603 78.3 ;
      RECT MASK 1 72.011 78.03 72.071 78.3 ;
      RECT MASK 1 72.343 78.03 72.403 78.3 ;
      RECT MASK 1 72.675 78.03 72.735 78.3 ;
      RECT MASK 1 73.173 78.03 73.233 78.3 ;
      RECT MASK 1 73.505 78.03 73.565 78.3 ;
      RECT MASK 1 73.837 78.03 73.897 78.3 ;
      RECT MASK 1 74.335 78.03 74.395 78.3 ;
      RECT MASK 1 74.667 78.03 74.727 78.3 ;
      RECT MASK 1 74.999 78.03 75.059 78.3 ;
      RECT MASK 1 75.497 78.03 75.557 78.3 ;
      RECT MASK 1 75.829 78.03 75.889 78.3 ;
      RECT MASK 1 76.161 78.03 76.221 78.3 ;
      RECT MASK 1 78.629 78.03 78.689 78.3 ;
      RECT MASK 1 78.961 78.03 79.021 78.3 ;
      RECT MASK 1 79.293 78.03 79.353 78.3 ;
      RECT MASK 1 79.791 78.03 79.851 78.3 ;
      RECT MASK 1 80.123 78.03 80.183 78.3 ;
      RECT MASK 1 80.455 78.03 80.515 78.3 ;
      RECT MASK 1 80.953 78.03 81.013 78.3 ;
      RECT MASK 1 81.285 78.03 81.345 78.3 ;
      RECT MASK 1 81.617 78.03 81.677 78.3 ;
      RECT MASK 1 82.115 78.03 82.175 78.3 ;
      RECT MASK 1 82.447 78.03 82.507 78.3 ;
      RECT MASK 1 82.779 78.03 82.839 78.3 ;
      RECT MASK 1 85.247 78.03 85.307 78.3 ;
      RECT MASK 1 85.579 78.03 85.639 78.3 ;
      RECT MASK 1 85.911 78.03 85.971 78.3 ;
      RECT MASK 1 86.409 78.03 86.469 78.3 ;
      RECT MASK 1 86.741 78.03 86.801 78.3 ;
      RECT MASK 1 87.073 78.03 87.133 78.3 ;
      RECT MASK 1 87.571 78.03 87.631 78.3 ;
      RECT MASK 1 87.903 78.03 87.963 78.3 ;
      RECT MASK 1 88.235 78.03 88.295 78.3 ;
      RECT MASK 1 88.733 78.03 88.793 78.3 ;
      RECT MASK 1 89.065 78.03 89.125 78.3 ;
      RECT MASK 1 89.397 78.03 89.457 78.3 ;
      RECT MASK 1 91.865 78.03 91.925 78.3 ;
      RECT MASK 1 92.197 78.03 92.257 78.3 ;
      RECT MASK 1 92.529 78.03 92.589 78.3 ;
      RECT MASK 1 93.027 78.03 93.087 78.3 ;
      RECT MASK 1 93.359 78.03 93.419 78.3 ;
      RECT MASK 1 93.691 78.03 93.751 78.3 ;
      RECT MASK 1 94.189 78.03 94.249 78.3 ;
      RECT MASK 1 94.521 78.03 94.581 78.3 ;
      RECT MASK 1 94.853 78.03 94.913 78.3 ;
      RECT MASK 1 95.351 78.03 95.411 78.3 ;
      RECT MASK 1 95.683 78.03 95.743 78.3 ;
      RECT MASK 1 96.015 78.03 96.075 78.3 ;
      RECT MASK 1 98.483 78.03 98.543 78.3 ;
      RECT MASK 1 98.815 78.03 98.875 78.3 ;
      RECT MASK 1 99.147 78.03 99.207 78.3 ;
      RECT MASK 1 99.645 78.03 99.705 78.3 ;
      RECT MASK 1 99.977 78.03 100.037 78.3 ;
      RECT MASK 1 100.309 78.03 100.369 78.3 ;
      RECT MASK 1 100.807 78.03 100.867 78.3 ;
      RECT MASK 1 101.139 78.03 101.199 78.3 ;
      RECT MASK 1 101.471 78.03 101.531 78.3 ;
      RECT MASK 1 101.969 78.03 102.029 78.3 ;
      RECT MASK 1 102.301 78.03 102.361 78.3 ;
      RECT MASK 1 102.633 78.03 102.693 78.3 ;
      RECT MASK 1 105.101 78.03 105.161 78.3 ;
      RECT MASK 1 105.433 78.03 105.493 78.3 ;
      RECT MASK 1 105.765 78.03 105.825 78.3 ;
      RECT MASK 1 106.263 78.03 106.323 78.3 ;
      RECT MASK 1 106.595 78.03 106.655 78.3 ;
      RECT MASK 1 106.927 78.03 106.987 78.3 ;
      RECT MASK 1 107.425 78.03 107.485 78.3 ;
      RECT MASK 1 107.757 78.03 107.817 78.3 ;
      RECT MASK 1 108.089 78.03 108.149 78.3 ;
      RECT MASK 1 108.587 78.03 108.647 78.3 ;
      RECT MASK 1 108.919 78.03 108.979 78.3 ;
      RECT MASK 1 109.251 78.03 109.311 78.3 ;
      RECT MASK 1 11.049 78.0305 11.109 80.25 ;
      RECT MASK 1 11.381 78.0305 11.441 80.25 ;
      RECT MASK 1 24.285 78.0305 24.345 80.25 ;
      RECT MASK 1 24.617 78.0305 24.677 80.25 ;
      RECT MASK 1 30.903 78.0305 30.963 80.25 ;
      RECT MASK 1 31.235 78.0305 31.295 80.25 ;
      RECT MASK 1 37.521 78.0305 37.581 80.25 ;
      RECT MASK 1 37.853 78.0305 37.913 80.25 ;
      RECT MASK 1 44.139 78.0305 44.199 80.25 ;
      RECT MASK 1 44.471 78.0305 44.531 80.25 ;
      RECT MASK 1 50.757 78.0305 50.817 80.25 ;
      RECT MASK 1 51.089 78.0305 51.149 80.25 ;
      RECT MASK 1 57.375 78.0305 57.435 80.25 ;
      RECT MASK 1 57.707 78.0305 57.767 80.25 ;
      RECT MASK 1 63.993 78.0305 64.053 80.25 ;
      RECT MASK 1 64.325 78.0305 64.385 80.25 ;
      RECT MASK 1 70.611 78.0305 70.671 80.25 ;
      RECT MASK 1 70.943 78.0305 71.003 80.25 ;
      RECT MASK 1 77.229 78.0305 77.289 80.25 ;
      RECT MASK 1 77.561 78.0305 77.621 80.25 ;
      RECT MASK 1 83.847 78.0305 83.907 80.25 ;
      RECT MASK 1 84.179 78.0305 84.239 80.25 ;
      RECT MASK 1 90.465 78.0305 90.525 80.25 ;
      RECT MASK 1 90.797 78.0305 90.857 80.25 ;
      RECT MASK 1 97.083 78.0305 97.143 80.25 ;
      RECT MASK 1 97.415 78.0305 97.475 80.25 ;
      RECT MASK 1 103.701 78.0305 103.761 80.25 ;
      RECT MASK 1 104.033 78.0305 104.093 80.25 ;
      RECT MASK 1 17.097 78.035 17.157 80.245 ;
      RECT MASK 1 23.715 78.035 23.775 80.245 ;
      RECT MASK 1 25.021 78.035 25.081 80.245 ;
      RECT MASK 1 70.041 78.035 70.101 80.28 ;
      RECT MASK 1 71.347 78.035 71.407 80.28 ;
      RECT MASK 1 109.749 78.035 109.809 80.245 ;
      RECT MASK 1 126.554 78.068 126.634 78.44 ;
      RECT MASK 1 1.263 78.44 1.363 96.411 ;
      RECT MASK 1 5.247 78.44 5.347 96.411 ;
      RECT MASK 1 6.983 78.586 7.063 81.8885 ;
      RECT MASK 1 7.315 78.586 7.395 81.8885 ;
      RECT MASK 1 8.145 78.586 8.225 81.8885 ;
      RECT MASK 1 8.477 78.586 8.557 81.8885 ;
      RECT MASK 1 9.307 78.586 9.387 81.8885 ;
      RECT MASK 1 9.639 78.586 9.719 81.8885 ;
      RECT MASK 1 12.439 78.586 12.519 81.8885 ;
      RECT MASK 1 12.771 78.586 12.851 81.8885 ;
      RECT MASK 1 13.601 78.586 13.681 81.8885 ;
      RECT MASK 1 13.933 78.586 14.013 81.8885 ;
      RECT MASK 1 14.763 78.586 14.843 81.8885 ;
      RECT MASK 1 15.095 78.586 15.175 81.8885 ;
      RECT MASK 1 15.925 78.586 16.005 81.8885 ;
      RECT MASK 1 16.257 78.586 16.337 81.8885 ;
      RECT MASK 1 19.057 78.586 19.137 81.8885 ;
      RECT MASK 1 19.389 78.586 19.469 81.8885 ;
      RECT MASK 1 20.219 78.586 20.299 81.8885 ;
      RECT MASK 1 20.551 78.586 20.631 81.8885 ;
      RECT MASK 1 21.381 78.586 21.461 81.8885 ;
      RECT MASK 1 21.713 78.586 21.793 81.8885 ;
      RECT MASK 1 22.543 78.586 22.623 81.8885 ;
      RECT MASK 1 22.875 78.586 22.955 81.8885 ;
      RECT MASK 1 25.675 78.586 25.755 81.8885 ;
      RECT MASK 1 26.007 78.586 26.087 81.8885 ;
      RECT MASK 1 26.837 78.586 26.917 81.8885 ;
      RECT MASK 1 27.169 78.586 27.249 81.8885 ;
      RECT MASK 1 27.999 78.586 28.079 81.8885 ;
      RECT MASK 1 28.331 78.586 28.411 81.8885 ;
      RECT MASK 1 29.161 78.586 29.241 81.8885 ;
      RECT MASK 1 29.493 78.586 29.573 81.8885 ;
      RECT MASK 1 32.293 78.586 32.373 81.8885 ;
      RECT MASK 1 32.625 78.586 32.705 81.8885 ;
      RECT MASK 1 33.455 78.586 33.535 81.8885 ;
      RECT MASK 1 33.787 78.586 33.867 81.8885 ;
      RECT MASK 1 34.617 78.586 34.697 81.8885 ;
      RECT MASK 1 34.949 78.586 35.029 81.8885 ;
      RECT MASK 1 35.779 78.586 35.859 81.8885 ;
      RECT MASK 1 36.111 78.586 36.191 81.8885 ;
      RECT MASK 1 38.911 78.586 38.991 81.8885 ;
      RECT MASK 1 39.243 78.586 39.323 81.8885 ;
      RECT MASK 1 40.073 78.586 40.153 81.8885 ;
      RECT MASK 1 40.405 78.586 40.485 81.8885 ;
      RECT MASK 1 41.235 78.586 41.315 81.8885 ;
      RECT MASK 1 41.567 78.586 41.647 81.8885 ;
      RECT MASK 1 42.397 78.586 42.477 81.8885 ;
      RECT MASK 1 42.729 78.586 42.809 81.8885 ;
      RECT MASK 1 45.529 78.586 45.609 81.8885 ;
      RECT MASK 1 45.861 78.586 45.941 81.8885 ;
      RECT MASK 1 46.691 78.586 46.771 81.8885 ;
      RECT MASK 1 47.023 78.586 47.103 81.8885 ;
      RECT MASK 1 47.853 78.586 47.933 81.8885 ;
      RECT MASK 1 48.185 78.586 48.265 81.8885 ;
      RECT MASK 1 49.015 78.586 49.095 81.8885 ;
      RECT MASK 1 49.347 78.586 49.427 81.8885 ;
      RECT MASK 1 52.147 78.586 52.227 81.8885 ;
      RECT MASK 1 52.479 78.586 52.559 81.8885 ;
      RECT MASK 1 53.309 78.586 53.389 81.8885 ;
      RECT MASK 1 53.641 78.586 53.721 81.8885 ;
      RECT MASK 1 54.471 78.586 54.551 81.8885 ;
      RECT MASK 1 54.803 78.586 54.883 81.8885 ;
      RECT MASK 1 55.633 78.586 55.713 81.8885 ;
      RECT MASK 1 55.965 78.586 56.045 81.8885 ;
      RECT MASK 1 58.765 78.586 58.845 81.8885 ;
      RECT MASK 1 59.097 78.586 59.177 81.8885 ;
      RECT MASK 1 59.927 78.586 60.007 81.8885 ;
      RECT MASK 1 60.259 78.586 60.339 81.8885 ;
      RECT MASK 1 61.089 78.586 61.169 81.8885 ;
      RECT MASK 1 61.421 78.586 61.501 81.8885 ;
      RECT MASK 1 62.251 78.586 62.331 81.8885 ;
      RECT MASK 1 62.583 78.586 62.663 81.8885 ;
      RECT MASK 1 65.383 78.586 65.463 81.8885 ;
      RECT MASK 1 65.715 78.586 65.795 81.8885 ;
      RECT MASK 1 66.545 78.586 66.625 81.8885 ;
      RECT MASK 1 66.877 78.586 66.957 81.8885 ;
      RECT MASK 1 67.707 78.586 67.787 81.8885 ;
      RECT MASK 1 68.039 78.586 68.119 81.8885 ;
      RECT MASK 1 68.869 78.586 68.949 81.8885 ;
      RECT MASK 1 69.201 78.586 69.281 81.8885 ;
      RECT MASK 1 72.001 78.586 72.081 81.8885 ;
      RECT MASK 1 72.333 78.586 72.413 81.8885 ;
      RECT MASK 1 73.163 78.586 73.243 81.8885 ;
      RECT MASK 1 73.495 78.586 73.575 81.8885 ;
      RECT MASK 1 74.325 78.586 74.405 81.8885 ;
      RECT MASK 1 74.657 78.586 74.737 81.8885 ;
      RECT MASK 1 75.487 78.586 75.567 81.8885 ;
      RECT MASK 1 75.819 78.586 75.899 81.8885 ;
      RECT MASK 1 78.619 78.586 78.699 81.8885 ;
      RECT MASK 1 78.951 78.586 79.031 81.8885 ;
      RECT MASK 1 79.781 78.586 79.861 81.8885 ;
      RECT MASK 1 80.113 78.586 80.193 81.8885 ;
      RECT MASK 1 80.943 78.586 81.023 81.8885 ;
      RECT MASK 1 81.275 78.586 81.355 81.8885 ;
      RECT MASK 1 82.105 78.586 82.185 81.8885 ;
      RECT MASK 1 82.437 78.586 82.517 81.8885 ;
      RECT MASK 1 85.237 78.586 85.317 81.8885 ;
      RECT MASK 1 85.569 78.586 85.649 81.8885 ;
      RECT MASK 1 86.399 78.586 86.479 81.8885 ;
      RECT MASK 1 86.731 78.586 86.811 81.8885 ;
      RECT MASK 1 87.561 78.586 87.641 81.8885 ;
      RECT MASK 1 87.893 78.586 87.973 81.8885 ;
      RECT MASK 1 88.723 78.586 88.803 81.8885 ;
      RECT MASK 1 89.055 78.586 89.135 81.8885 ;
      RECT MASK 1 91.855 78.586 91.935 81.8885 ;
      RECT MASK 1 92.187 78.586 92.267 81.8885 ;
      RECT MASK 1 93.017 78.586 93.097 81.8885 ;
      RECT MASK 1 93.349 78.586 93.429 81.8885 ;
      RECT MASK 1 94.179 78.586 94.259 81.8885 ;
      RECT MASK 1 94.511 78.586 94.591 81.8885 ;
      RECT MASK 1 95.341 78.586 95.421 81.8885 ;
      RECT MASK 1 95.673 78.586 95.753 81.8885 ;
      RECT MASK 1 98.473 78.586 98.553 81.8885 ;
      RECT MASK 1 98.805 78.586 98.885 81.8885 ;
      RECT MASK 1 99.635 78.586 99.715 81.8885 ;
      RECT MASK 1 99.967 78.586 100.047 81.8885 ;
      RECT MASK 1 100.797 78.586 100.877 81.8885 ;
      RECT MASK 1 101.129 78.586 101.209 81.8885 ;
      RECT MASK 1 101.959 78.586 102.039 81.8885 ;
      RECT MASK 1 102.291 78.586 102.371 81.8885 ;
      RECT MASK 1 105.091 78.586 105.171 81.8885 ;
      RECT MASK 1 105.423 78.586 105.503 81.8885 ;
      RECT MASK 1 106.253 78.586 106.333 81.8885 ;
      RECT MASK 1 106.585 78.586 106.665 81.8885 ;
      RECT MASK 1 107.415 78.586 107.495 81.8885 ;
      RECT MASK 1 107.747 78.586 107.827 81.8885 ;
      RECT MASK 1 108.577 78.586 108.657 81.8885 ;
      RECT MASK 1 108.909 78.586 108.989 81.8885 ;
      RECT MASK 1 116.261 78.635 116.341 78.937 ;
      RECT MASK 1 116.593 78.635 116.673 78.937 ;
      RECT MASK 1 116.925 78.635 117.005 78.937 ;
      RECT MASK 1 117.257 78.635 117.337 78.937 ;
      RECT MASK 1 117.589 78.635 117.669 78.937 ;
      RECT MASK 1 117.921 78.635 118.001 78.937 ;
      RECT MASK 1 118.253 78.635 118.333 78.937 ;
      RECT MASK 1 118.585 78.635 118.665 78.937 ;
      RECT MASK 1 118.917 78.635 118.997 78.937 ;
      RECT MASK 1 119.249 78.635 119.329 78.937 ;
      RECT MASK 1 119.581 78.635 119.661 78.937 ;
      RECT MASK 1 119.913 78.635 119.993 78.937 ;
      RECT MASK 1 120.245 78.635 120.325 78.937 ;
      RECT MASK 1 120.577 78.635 120.657 78.937 ;
      RECT MASK 1 120.909 78.635 120.989 78.937 ;
      RECT MASK 1 121.241 78.635 121.321 78.937 ;
      RECT MASK 1 121.573 78.635 121.653 78.937 ;
      RECT MASK 1 121.905 78.635 121.985 78.937 ;
      RECT MASK 1 122.237 78.635 122.317 78.937 ;
      RECT MASK 1 122.569 78.635 122.649 78.937 ;
      RECT MASK 1 122.901 78.635 122.981 78.937 ;
      RECT MASK 1 123.233 78.635 123.313 78.937 ;
      RECT MASK 1 123.565 78.635 123.645 78.937 ;
      RECT MASK 1 123.897 78.635 123.977 78.937 ;
      RECT MASK 1 124.229 78.635 124.309 78.937 ;
      RECT MASK 1 124.561 78.635 124.641 78.937 ;
      RECT MASK 1 124.893 78.635 124.973 78.937 ;
      RECT MASK 1 125.225 78.635 125.305 78.937 ;
      RECT MASK 1 125.557 78.635 125.637 78.937 ;
      RECT MASK 1 125.889 78.635 125.969 78.937 ;
      RECT MASK 1 126.221 78.635 126.301 78.937 ;
      RECT MASK 1 111.211 78.785 111.271 80.512 ;
      RECT MASK 1 111.543 78.785 111.603 79.045 ;
      RECT MASK 1 111.875 78.785 111.935 79.045 ;
      RECT MASK 1 112.207 78.785 112.267 79.045 ;
      RECT MASK 1 112.539 78.785 112.599 79.045 ;
      RECT MASK 1 112.871 78.785 112.931 79.045 ;
      RECT MASK 1 113.203 78.785 113.263 80.512 ;
      RECT MASK 1 126.554 78.848 126.634 79.22 ;
      RECT MASK 1 7.657 78.981 7.717 82.34 ;
      RECT MASK 1 8.819 78.981 8.879 82.34 ;
      RECT MASK 1 9.981 78.981 10.041 82.34 ;
      RECT MASK 1 13.113 78.981 13.173 82.34 ;
      RECT MASK 1 14.275 78.981 14.335 82.34 ;
      RECT MASK 1 15.437 78.981 15.497 82.34 ;
      RECT MASK 1 16.599 78.981 16.659 82.34 ;
      RECT MASK 1 19.731 78.981 19.791 82.34 ;
      RECT MASK 1 20.893 78.981 20.953 82.34 ;
      RECT MASK 1 22.055 78.981 22.115 82.34 ;
      RECT MASK 1 23.217 78.981 23.277 82.34 ;
      RECT MASK 1 26.349 78.981 26.409 82.34 ;
      RECT MASK 1 27.511 78.981 27.571 82.34 ;
      RECT MASK 1 28.673 78.981 28.733 82.34 ;
      RECT MASK 1 29.835 78.981 29.895 82.34 ;
      RECT MASK 1 32.967 78.981 33.027 82.34 ;
      RECT MASK 1 34.129 78.981 34.189 82.34 ;
      RECT MASK 1 35.291 78.981 35.351 82.34 ;
      RECT MASK 1 36.453 78.981 36.513 82.34 ;
      RECT MASK 1 39.585 78.981 39.645 82.34 ;
      RECT MASK 1 40.747 78.981 40.807 82.34 ;
      RECT MASK 1 41.909 78.981 41.969 82.34 ;
      RECT MASK 1 43.071 78.981 43.131 82.34 ;
      RECT MASK 1 46.203 78.981 46.263 82.34 ;
      RECT MASK 1 47.365 78.981 47.425 82.34 ;
      RECT MASK 1 48.527 78.981 48.587 82.34 ;
      RECT MASK 1 49.689 78.981 49.749 82.34 ;
      RECT MASK 1 52.821 78.981 52.881 82.34 ;
      RECT MASK 1 53.983 78.981 54.043 82.34 ;
      RECT MASK 1 55.145 78.981 55.205 82.34 ;
      RECT MASK 1 56.307 78.981 56.367 82.34 ;
      RECT MASK 1 59.439 78.981 59.499 82.34 ;
      RECT MASK 1 60.601 78.981 60.661 82.34 ;
      RECT MASK 1 61.763 78.981 61.823 82.34 ;
      RECT MASK 1 62.925 78.981 62.985 82.34 ;
      RECT MASK 1 66.057 78.981 66.117 82.34 ;
      RECT MASK 1 67.219 78.981 67.279 82.34 ;
      RECT MASK 1 68.381 78.981 68.441 82.34 ;
      RECT MASK 1 69.543 78.981 69.603 82.34 ;
      RECT MASK 1 72.675 78.981 72.735 82.34 ;
      RECT MASK 1 73.837 78.981 73.897 82.34 ;
      RECT MASK 1 74.999 78.981 75.059 82.34 ;
      RECT MASK 1 76.161 78.981 76.221 82.34 ;
      RECT MASK 1 79.293 78.981 79.353 82.34 ;
      RECT MASK 1 80.455 78.981 80.515 82.34 ;
      RECT MASK 1 81.617 78.981 81.677 82.34 ;
      RECT MASK 1 82.779 78.981 82.839 82.34 ;
      RECT MASK 1 85.911 78.981 85.971 82.34 ;
      RECT MASK 1 87.073 78.981 87.133 82.34 ;
      RECT MASK 1 88.235 78.981 88.295 82.34 ;
      RECT MASK 1 89.397 78.981 89.457 82.34 ;
      RECT MASK 1 92.529 78.981 92.589 82.34 ;
      RECT MASK 1 93.691 78.981 93.751 82.34 ;
      RECT MASK 1 94.853 78.981 94.913 82.34 ;
      RECT MASK 1 96.015 78.981 96.075 82.34 ;
      RECT MASK 1 99.147 78.981 99.207 82.34 ;
      RECT MASK 1 100.309 78.981 100.369 82.34 ;
      RECT MASK 1 101.471 78.981 101.531 82.34 ;
      RECT MASK 1 102.633 78.981 102.693 82.34 ;
      RECT MASK 1 105.765 78.981 105.825 82.34 ;
      RECT MASK 1 106.927 78.981 106.987 82.34 ;
      RECT MASK 1 108.089 78.981 108.149 82.34 ;
      RECT MASK 1 109.251 78.981 109.311 82.34 ;
      RECT MASK 1 2.067 79.05 2.127 95.882 ;
      RECT MASK 1 2.341 79.05 2.401 95.88 ;
      RECT MASK 1 2.615 79.05 2.675 95.88 ;
      RECT MASK 1 2.889 79.05 2.949 95.88 ;
      RECT MASK 1 3.163 79.05 3.223 95.88 ;
      RECT MASK 1 3.437 79.05 3.497 95.88 ;
      RECT MASK 1 3.711 79.05 3.771 95.88 ;
      RECT MASK 1 3.985 79.05 4.045 95.88 ;
      RECT MASK 1 4.259 79.05 4.319 95.88 ;
      RECT MASK 1 4.533 79.05 4.593 95.882 ;
      RECT MASK 1 111.958 79.29 112.018 79.559 ;
      RECT MASK 1 112.622 79.29 112.682 79.559 ;
      RECT MASK 1 116.261 79.415 116.341 79.717 ;
      RECT MASK 1 116.593 79.415 116.673 79.717 ;
      RECT MASK 1 116.925 79.415 117.005 79.717 ;
      RECT MASK 1 117.257 79.415 117.337 79.717 ;
      RECT MASK 1 117.589 79.415 117.669 79.717 ;
      RECT MASK 1 117.921 79.415 118.001 79.717 ;
      RECT MASK 1 118.253 79.415 118.333 79.717 ;
      RECT MASK 1 118.585 79.415 118.665 79.717 ;
      RECT MASK 1 118.917 79.415 118.997 79.717 ;
      RECT MASK 1 119.249 79.415 119.329 79.717 ;
      RECT MASK 1 119.581 79.415 119.661 79.717 ;
      RECT MASK 1 119.913 79.415 119.993 79.717 ;
      RECT MASK 1 120.245 79.415 120.325 79.717 ;
      RECT MASK 1 120.577 79.415 120.657 79.717 ;
      RECT MASK 1 120.909 79.415 120.989 79.717 ;
      RECT MASK 1 121.241 79.415 121.321 79.717 ;
      RECT MASK 1 121.573 79.415 121.653 79.717 ;
      RECT MASK 1 121.905 79.415 121.985 79.717 ;
      RECT MASK 1 122.237 79.415 122.317 79.717 ;
      RECT MASK 1 122.569 79.415 122.649 79.717 ;
      RECT MASK 1 122.901 79.415 122.981 79.717 ;
      RECT MASK 1 123.233 79.415 123.313 79.717 ;
      RECT MASK 1 123.565 79.415 123.645 79.717 ;
      RECT MASK 1 123.897 79.415 123.977 79.717 ;
      RECT MASK 1 124.229 79.415 124.309 79.717 ;
      RECT MASK 1 124.561 79.415 124.641 79.717 ;
      RECT MASK 1 124.893 79.415 124.973 79.717 ;
      RECT MASK 1 125.225 79.415 125.305 79.717 ;
      RECT MASK 1 125.557 79.415 125.637 79.717 ;
      RECT MASK 1 125.889 79.415 125.969 79.717 ;
      RECT MASK 1 126.221 79.415 126.301 79.717 ;
      RECT MASK 1 10.23 79.57 10.29 79.79 ;
      RECT MASK 1 12.034 79.57 12.094 79.79 ;
      RECT MASK 1 16.848 79.57 16.908 79.79 ;
      RECT MASK 1 18.652 79.57 18.712 79.79 ;
      RECT MASK 1 23.466 79.57 23.526 79.79 ;
      RECT MASK 1 25.27 79.57 25.33 79.79 ;
      RECT MASK 1 30.084 79.57 30.144 79.79 ;
      RECT MASK 1 31.888 79.57 31.948 79.79 ;
      RECT MASK 1 36.702 79.57 36.762 79.79 ;
      RECT MASK 1 38.506 79.57 38.566 79.79 ;
      RECT MASK 1 43.32 79.57 43.38 79.79 ;
      RECT MASK 1 45.124 79.57 45.184 79.79 ;
      RECT MASK 1 49.938 79.57 49.998 79.79 ;
      RECT MASK 1 51.742 79.57 51.802 79.79 ;
      RECT MASK 1 56.556 79.57 56.616 79.79 ;
      RECT MASK 1 58.36 79.57 58.42 79.79 ;
      RECT MASK 1 63.174 79.57 63.234 79.79 ;
      RECT MASK 1 64.978 79.57 65.038 79.79 ;
      RECT MASK 1 69.792 79.57 69.852 79.79 ;
      RECT MASK 1 71.596 79.57 71.656 79.79 ;
      RECT MASK 1 76.41 79.57 76.47 79.79 ;
      RECT MASK 1 78.214 79.57 78.274 79.79 ;
      RECT MASK 1 83.028 79.57 83.088 79.79 ;
      RECT MASK 1 84.832 79.57 84.892 79.79 ;
      RECT MASK 1 89.646 79.57 89.706 79.79 ;
      RECT MASK 1 91.45 79.57 91.51 79.79 ;
      RECT MASK 1 96.264 79.57 96.324 79.79 ;
      RECT MASK 1 98.068 79.57 98.128 79.79 ;
      RECT MASK 1 102.882 79.57 102.942 79.79 ;
      RECT MASK 1 104.686 79.57 104.746 79.79 ;
      RECT MASK 1 109.5 79.57 109.56 79.79 ;
      RECT MASK 1 112.456 79.579 112.516 81.511 ;
      RECT MASK 1 126.554 79.628 126.634 80 ;
      RECT MASK 1 111.958 79.679 112.018 81.611 ;
      RECT MASK 1 116.261 80.126 116.341 80.458 ;
      RECT MASK 1 116.593 80.126 116.673 80.458 ;
      RECT MASK 1 116.925 80.126 117.005 80.458 ;
      RECT MASK 1 117.257 80.126 117.337 80.458 ;
      RECT MASK 1 117.589 80.126 117.669 80.458 ;
      RECT MASK 1 117.921 80.126 118.001 80.458 ;
      RECT MASK 1 118.253 80.126 118.333 80.458 ;
      RECT MASK 1 118.585 80.126 118.665 80.458 ;
      RECT MASK 1 118.917 80.126 118.997 80.458 ;
      RECT MASK 1 119.249 80.126 119.329 80.458 ;
      RECT MASK 1 119.581 80.126 119.661 80.458 ;
      RECT MASK 1 119.913 80.126 119.993 80.458 ;
      RECT MASK 1 120.245 80.126 120.325 80.458 ;
      RECT MASK 1 120.577 80.126 120.657 80.458 ;
      RECT MASK 1 120.909 80.126 120.989 80.458 ;
      RECT MASK 1 121.241 80.126 121.321 80.458 ;
      RECT MASK 1 121.573 80.126 121.653 80.458 ;
      RECT MASK 1 121.905 80.126 121.985 80.458 ;
      RECT MASK 1 122.237 80.126 122.317 80.458 ;
      RECT MASK 1 122.569 80.126 122.649 80.458 ;
      RECT MASK 1 122.901 80.126 122.981 80.458 ;
      RECT MASK 1 123.233 80.126 123.313 80.458 ;
      RECT MASK 1 123.565 80.126 123.645 80.458 ;
      RECT MASK 1 123.897 80.126 123.977 80.458 ;
      RECT MASK 1 124.229 80.126 124.309 80.458 ;
      RECT MASK 1 124.561 80.126 124.641 80.458 ;
      RECT MASK 1 124.893 80.126 124.973 80.458 ;
      RECT MASK 1 125.225 80.126 125.305 80.458 ;
      RECT MASK 1 125.557 80.126 125.637 80.458 ;
      RECT MASK 1 125.889 80.126 125.969 80.458 ;
      RECT MASK 1 126.221 80.126 126.301 80.458 ;
      RECT MASK 1 6.329 80.423 6.389 82.645 ;
      RECT MASK 1 58.277 80.43 58.337 84.169 ;
      RECT MASK 1 11.785 80.4335 11.845 82.645 ;
      RECT MASK 1 17.097 80.4335 17.157 82.645 ;
      RECT MASK 1 58.111 80.4335 58.171 84.164 ;
      RECT MASK 1 63.423 80.4335 63.483 84.164 ;
      RECT MASK 1 103.131 80.4335 103.191 82.645 ;
      RECT MASK 1 109.749 80.4335 109.809 82.645 ;
      RECT MASK 1 10.479 80.435 10.539 82.645 ;
      RECT MASK 1 11.049 80.4655 11.109 84.157 ;
      RECT MASK 1 11.381 80.4655 11.441 84.157 ;
      RECT MASK 1 17.667 80.4655 17.727 84.157 ;
      RECT MASK 1 17.999 80.4655 18.059 84.157 ;
      RECT MASK 1 24.285 80.4655 24.345 84.157 ;
      RECT MASK 1 24.617 80.4655 24.677 84.157 ;
      RECT MASK 1 30.903 80.4655 30.963 84.157 ;
      RECT MASK 1 31.235 80.4655 31.295 84.157 ;
      RECT MASK 1 37.521 80.4655 37.581 84.157 ;
      RECT MASK 1 37.853 80.4655 37.913 84.157 ;
      RECT MASK 1 44.139 80.4655 44.199 84.157 ;
      RECT MASK 1 44.471 80.4655 44.531 84.157 ;
      RECT MASK 1 50.757 80.4655 50.817 84.157 ;
      RECT MASK 1 51.089 80.4655 51.149 84.157 ;
      RECT MASK 1 57.375 80.4655 57.435 84.157 ;
      RECT MASK 1 57.707 80.4655 57.767 84.157 ;
      RECT MASK 1 63.993 80.4655 64.053 84.157 ;
      RECT MASK 1 64.325 80.4655 64.385 84.157 ;
      RECT MASK 1 70.611 80.4655 70.671 84.157 ;
      RECT MASK 1 70.943 80.4655 71.003 84.157 ;
      RECT MASK 1 77.229 80.4655 77.289 84.157 ;
      RECT MASK 1 77.561 80.4655 77.621 84.157 ;
      RECT MASK 1 83.847 80.4655 83.907 84.157 ;
      RECT MASK 1 84.179 80.4655 84.239 84.157 ;
      RECT MASK 1 90.465 80.4655 90.525 84.157 ;
      RECT MASK 1 90.797 80.4655 90.857 84.157 ;
      RECT MASK 1 97.083 80.4655 97.143 84.157 ;
      RECT MASK 1 97.415 80.4655 97.475 84.157 ;
      RECT MASK 1 103.701 80.4655 103.761 84.157 ;
      RECT MASK 1 104.033 80.4655 104.093 84.157 ;
      RECT MASK 1 111.211 80.708 111.271 82.405 ;
      RECT MASK 1 113.203 80.708 113.263 82.405 ;
      RECT MASK 1 128.41 81.229 128.51 107.66 ;
      RECT MASK 1 115.628 81.23 115.728 87.081 ;
      RECT MASK 1 10.23 81.294 10.29 81.514 ;
      RECT MASK 1 12.034 81.294 12.094 81.514 ;
      RECT MASK 1 16.848 81.294 16.908 81.514 ;
      RECT MASK 1 18.652 81.294 18.712 81.514 ;
      RECT MASK 1 23.466 81.294 23.526 81.514 ;
      RECT MASK 1 25.27 81.294 25.33 81.514 ;
      RECT MASK 1 30.084 81.294 30.144 81.514 ;
      RECT MASK 1 31.888 81.294 31.948 81.514 ;
      RECT MASK 1 36.702 81.294 36.762 81.514 ;
      RECT MASK 1 38.506 81.294 38.566 81.514 ;
      RECT MASK 1 43.32 81.294 43.38 81.514 ;
      RECT MASK 1 45.124 81.294 45.184 81.514 ;
      RECT MASK 1 49.938 81.294 49.998 81.514 ;
      RECT MASK 1 51.742 81.294 51.802 81.514 ;
      RECT MASK 1 56.556 81.294 56.616 81.514 ;
      RECT MASK 1 60.767 81.294 60.827 81.514 ;
      RECT MASK 1 63.174 81.294 63.234 81.514 ;
      RECT MASK 1 64.978 81.294 65.038 81.514 ;
      RECT MASK 1 69.792 81.294 69.852 81.514 ;
      RECT MASK 1 71.596 81.294 71.656 81.514 ;
      RECT MASK 1 76.41 81.294 76.47 81.514 ;
      RECT MASK 1 78.214 81.294 78.274 81.514 ;
      RECT MASK 1 83.028 81.294 83.088 81.514 ;
      RECT MASK 1 84.832 81.294 84.892 81.514 ;
      RECT MASK 1 89.646 81.294 89.706 81.514 ;
      RECT MASK 1 91.45 81.294 91.51 81.514 ;
      RECT MASK 1 96.264 81.294 96.324 81.514 ;
      RECT MASK 1 98.068 81.294 98.128 81.514 ;
      RECT MASK 1 102.882 81.294 102.942 81.514 ;
      RECT MASK 1 104.686 81.294 104.746 81.514 ;
      RECT MASK 1 109.5 81.294 109.56 81.514 ;
      RECT MASK 1 103.361 81.302 103.421 82.929 ;
      RECT MASK 1 112.456 81.631 112.516 81.925 ;
      RECT MASK 1 116.462 81.82 116.522 86.7 ;
      RECT MASK 1 116.736 81.84 116.796 96.66 ;
      RECT MASK 1 117.01 81.84 117.07 96.66 ;
      RECT MASK 1 117.284 81.84 117.344 96.66 ;
      RECT MASK 1 117.558 81.84 117.618 96.66 ;
      RECT MASK 1 117.832 81.84 117.892 96.66 ;
      RECT MASK 1 118.106 81.84 118.166 96.66 ;
      RECT MASK 1 118.38 81.84 118.44 96.66 ;
      RECT MASK 1 118.654 81.84 118.714 96.66 ;
      RECT MASK 1 118.928 81.84 118.988 96.66 ;
      RECT MASK 1 119.202 81.84 119.262 96.66 ;
      RECT MASK 1 119.476 81.84 119.536 96.66 ;
      RECT MASK 1 119.75 81.84 119.81 96.66 ;
      RECT MASK 1 120.024 81.84 120.084 96.66 ;
      RECT MASK 1 120.298 81.84 120.358 96.66 ;
      RECT MASK 1 120.572 81.84 120.632 96.66 ;
      RECT MASK 1 120.846 81.84 120.906 96.66 ;
      RECT MASK 1 121.12 81.84 121.18 96.66 ;
      RECT MASK 1 121.394 81.84 121.454 96.66 ;
      RECT MASK 1 121.668 81.84 121.728 96.66 ;
      RECT MASK 1 121.942 81.84 122.002 96.66 ;
      RECT MASK 1 122.216 81.84 122.276 96.66 ;
      RECT MASK 1 122.49 81.84 122.55 96.66 ;
      RECT MASK 1 122.764 81.84 122.824 96.66 ;
      RECT MASK 1 123.038 81.84 123.098 96.66 ;
      RECT MASK 1 123.312 81.84 123.372 96.66 ;
      RECT MASK 1 123.586 81.84 123.646 96.66 ;
      RECT MASK 1 123.86 81.84 123.92 96.66 ;
      RECT MASK 1 124.134 81.84 124.194 96.66 ;
      RECT MASK 1 124.408 81.84 124.468 96.66 ;
      RECT MASK 1 124.682 81.84 124.742 96.66 ;
      RECT MASK 1 124.956 81.84 125.016 96.66 ;
      RECT MASK 1 125.23 81.84 125.29 96.66 ;
      RECT MASK 1 125.504 81.84 125.564 96.66 ;
      RECT MASK 1 125.778 81.84 125.838 96.66 ;
      RECT MASK 1 126.052 81.84 126.112 96.66 ;
      RECT MASK 1 126.326 81.84 126.386 96.66 ;
      RECT MASK 1 126.6 81.84 126.66 96.66 ;
      RECT MASK 1 126.874 81.84 126.934 96.66 ;
      RECT MASK 1 127.148 81.84 127.208 96.66 ;
      RECT MASK 1 127.422 81.84 127.482 96.66 ;
      RECT MASK 1 127.696 81.84 127.756 86.7 ;
      RECT MASK 1 63.257 81.893 63.317 84.157 ;
      RECT MASK 1 58.609 82.013 58.669 82.675 ;
      RECT MASK 1 59.024 82.013 59.084 84.157 ;
      RECT MASK 1 59.771 82.013 59.831 82.675 ;
      RECT MASK 1 60.933 82.013 60.993 82.675 ;
      RECT MASK 1 62.095 82.013 62.155 82.675 ;
      RECT MASK 1 60.141 82.133 60.291 84.157 ;
      RECT MASK 1 61.303 82.133 61.453 84.157 ;
      RECT MASK 1 62.465 82.133 62.615 84.157 ;
      RECT MASK 1 111.543 82.145 111.603 82.405 ;
      RECT MASK 1 111.875 82.145 111.935 82.405 ;
      RECT MASK 1 112.207 82.145 112.267 82.405 ;
      RECT MASK 1 112.539 82.145 112.599 82.405 ;
      RECT MASK 1 112.871 82.145 112.931 82.405 ;
      RECT MASK 1 6.827 82.38 6.887 82.65 ;
      RECT MASK 1 7.989 82.38 8.049 82.65 ;
      RECT MASK 1 9.151 82.38 9.211 82.65 ;
      RECT MASK 1 12.283 82.38 12.343 82.65 ;
      RECT MASK 1 13.445 82.38 13.505 82.65 ;
      RECT MASK 1 14.607 82.38 14.667 82.65 ;
      RECT MASK 1 15.769 82.38 15.829 82.65 ;
      RECT MASK 1 18.901 82.38 18.961 82.65 ;
      RECT MASK 1 20.063 82.38 20.123 82.65 ;
      RECT MASK 1 21.225 82.38 21.285 82.65 ;
      RECT MASK 1 22.387 82.38 22.447 82.65 ;
      RECT MASK 1 25.519 82.38 25.579 82.65 ;
      RECT MASK 1 26.681 82.38 26.741 82.65 ;
      RECT MASK 1 27.843 82.38 27.903 82.65 ;
      RECT MASK 1 29.005 82.38 29.065 82.65 ;
      RECT MASK 1 32.137 82.38 32.197 82.65 ;
      RECT MASK 1 33.299 82.38 33.359 82.65 ;
      RECT MASK 1 34.461 82.38 34.521 82.65 ;
      RECT MASK 1 35.623 82.38 35.683 82.65 ;
      RECT MASK 1 38.755 82.38 38.815 82.65 ;
      RECT MASK 1 39.917 82.38 39.977 82.65 ;
      RECT MASK 1 41.079 82.38 41.139 82.65 ;
      RECT MASK 1 42.241 82.38 42.301 82.65 ;
      RECT MASK 1 45.373 82.38 45.433 82.65 ;
      RECT MASK 1 46.535 82.38 46.595 82.65 ;
      RECT MASK 1 47.697 82.38 47.757 82.65 ;
      RECT MASK 1 48.859 82.38 48.919 82.65 ;
      RECT MASK 1 51.991 82.38 52.051 82.65 ;
      RECT MASK 1 53.153 82.38 53.213 82.65 ;
      RECT MASK 1 54.315 82.38 54.375 82.65 ;
      RECT MASK 1 55.477 82.38 55.537 82.65 ;
      RECT MASK 1 65.227 82.38 65.287 82.65 ;
      RECT MASK 1 66.389 82.38 66.449 82.65 ;
      RECT MASK 1 67.551 82.38 67.611 82.65 ;
      RECT MASK 1 68.713 82.38 68.773 82.65 ;
      RECT MASK 1 71.845 82.38 71.905 82.65 ;
      RECT MASK 1 73.007 82.38 73.067 82.65 ;
      RECT MASK 1 74.169 82.38 74.229 82.65 ;
      RECT MASK 1 75.331 82.38 75.391 82.65 ;
      RECT MASK 1 78.463 82.38 78.523 82.65 ;
      RECT MASK 1 79.625 82.38 79.685 82.65 ;
      RECT MASK 1 80.787 82.38 80.847 82.65 ;
      RECT MASK 1 81.949 82.38 82.009 82.65 ;
      RECT MASK 1 85.081 82.38 85.141 82.65 ;
      RECT MASK 1 86.243 82.38 86.303 82.65 ;
      RECT MASK 1 87.405 82.38 87.465 82.65 ;
      RECT MASK 1 88.567 82.38 88.627 82.65 ;
      RECT MASK 1 91.699 82.38 91.759 82.65 ;
      RECT MASK 1 92.861 82.38 92.921 82.65 ;
      RECT MASK 1 94.023 82.38 94.083 82.65 ;
      RECT MASK 1 95.185 82.38 95.245 82.65 ;
      RECT MASK 1 98.317 82.38 98.377 82.65 ;
      RECT MASK 1 99.479 82.38 99.539 82.65 ;
      RECT MASK 1 100.641 82.38 100.701 82.65 ;
      RECT MASK 1 101.803 82.38 101.863 82.65 ;
      RECT MASK 1 104.935 82.38 104.995 82.65 ;
      RECT MASK 1 106.097 82.38 106.157 82.65 ;
      RECT MASK 1 107.259 82.38 107.319 82.65 ;
      RECT MASK 1 108.421 82.38 108.481 82.65 ;
      RECT MASK 1 59.356 82.475 59.416 83.189 ;
      RECT MASK 1 60.498 82.475 60.598 83.189 ;
      RECT MASK 1 61.66 82.475 61.76 83.189 ;
      RECT MASK 1 62.822 82.475 62.922 83.189 ;
      RECT MASK 1 6.329 82.77 6.389 84.164 ;
      RECT MASK 1 10.479 82.77 10.539 84.164 ;
      RECT MASK 1 11.785 82.77 11.845 84.164 ;
      RECT MASK 1 17.097 82.77 17.157 84.164 ;
      RECT MASK 1 18.403 82.77 18.463 84.164 ;
      RECT MASK 1 23.715 82.77 23.775 84.164 ;
      RECT MASK 1 25.021 82.77 25.081 84.164 ;
      RECT MASK 1 30.333 82.77 30.393 84.164 ;
      RECT MASK 1 31.639 82.77 31.699 84.164 ;
      RECT MASK 1 36.951 82.77 37.011 84.164 ;
      RECT MASK 1 38.257 82.77 38.317 84.164 ;
      RECT MASK 1 43.569 82.77 43.629 84.164 ;
      RECT MASK 1 44.875 82.77 44.935 84.164 ;
      RECT MASK 1 50.187 82.77 50.247 84.164 ;
      RECT MASK 1 51.493 82.77 51.553 84.164 ;
      RECT MASK 1 56.805 82.77 56.865 84.164 ;
      RECT MASK 1 64.729 82.77 64.789 84.164 ;
      RECT MASK 1 70.041 82.77 70.101 84.164 ;
      RECT MASK 1 71.347 82.77 71.407 84.164 ;
      RECT MASK 1 76.659 82.77 76.719 84.164 ;
      RECT MASK 1 77.965 82.77 78.025 84.164 ;
      RECT MASK 1 83.277 82.77 83.337 84.164 ;
      RECT MASK 1 84.583 82.77 84.643 84.164 ;
      RECT MASK 1 89.895 82.77 89.955 84.164 ;
      RECT MASK 1 91.201 82.77 91.261 84.164 ;
      RECT MASK 1 96.513 82.77 96.573 84.164 ;
      RECT MASK 1 97.819 82.77 97.879 84.164 ;
      RECT MASK 1 103.131 82.77 103.191 84.164 ;
      RECT MASK 1 104.437 82.77 104.497 84.164 ;
      RECT MASK 1 109.749 82.77 109.809 84.164 ;
      RECT MASK 1 6.91 82.895 6.97 83.189 ;
      RECT MASK 1 7.574 82.895 7.634 83.189 ;
      RECT MASK 1 8.072 82.895 8.132 83.189 ;
      RECT MASK 1 8.736 82.895 8.796 83.189 ;
      RECT MASK 1 9.234 82.895 9.294 83.189 ;
      RECT MASK 1 9.898 82.895 9.958 83.189 ;
      RECT MASK 1 12.366 82.895 12.426 83.189 ;
      RECT MASK 1 13.03 82.895 13.09 83.189 ;
      RECT MASK 1 13.528 82.895 13.588 83.189 ;
      RECT MASK 1 14.192 82.895 14.252 83.189 ;
      RECT MASK 1 14.69 82.895 14.75 83.189 ;
      RECT MASK 1 15.354 82.895 15.414 83.189 ;
      RECT MASK 1 15.852 82.895 15.912 83.189 ;
      RECT MASK 1 16.516 82.895 16.576 83.189 ;
      RECT MASK 1 18.984 82.895 19.044 83.189 ;
      RECT MASK 1 19.648 82.895 19.708 83.189 ;
      RECT MASK 1 20.146 82.895 20.206 83.189 ;
      RECT MASK 1 20.81 82.895 20.87 83.189 ;
      RECT MASK 1 21.308 82.895 21.368 83.189 ;
      RECT MASK 1 21.972 82.895 22.032 83.189 ;
      RECT MASK 1 22.47 82.895 22.53 83.189 ;
      RECT MASK 1 23.134 82.895 23.194 83.189 ;
      RECT MASK 1 25.602 82.895 25.662 83.189 ;
      RECT MASK 1 26.266 82.895 26.326 83.189 ;
      RECT MASK 1 26.764 82.895 26.824 83.189 ;
      RECT MASK 1 27.428 82.895 27.488 83.189 ;
      RECT MASK 1 27.926 82.895 27.986 83.189 ;
      RECT MASK 1 28.59 82.895 28.65 83.189 ;
      RECT MASK 1 29.088 82.895 29.148 83.189 ;
      RECT MASK 1 29.752 82.895 29.812 83.189 ;
      RECT MASK 1 32.22 82.895 32.28 83.189 ;
      RECT MASK 1 32.884 82.895 32.944 83.189 ;
      RECT MASK 1 33.382 82.895 33.442 83.189 ;
      RECT MASK 1 34.046 82.895 34.106 83.189 ;
      RECT MASK 1 34.544 82.895 34.604 83.189 ;
      RECT MASK 1 35.208 82.895 35.268 83.189 ;
      RECT MASK 1 35.706 82.895 35.766 83.189 ;
      RECT MASK 1 36.37 82.895 36.43 83.189 ;
      RECT MASK 1 38.838 82.895 38.898 83.189 ;
      RECT MASK 1 39.502 82.895 39.562 83.189 ;
      RECT MASK 1 40 82.895 40.06 83.189 ;
      RECT MASK 1 40.664 82.895 40.724 83.189 ;
      RECT MASK 1 41.162 82.895 41.222 83.189 ;
      RECT MASK 1 41.826 82.895 41.886 83.189 ;
      RECT MASK 1 42.324 82.895 42.384 83.189 ;
      RECT MASK 1 42.988 82.895 43.048 83.189 ;
      RECT MASK 1 45.456 82.895 45.516 83.189 ;
      RECT MASK 1 46.12 82.895 46.18 83.189 ;
      RECT MASK 1 46.618 82.895 46.678 83.189 ;
      RECT MASK 1 47.282 82.895 47.342 83.189 ;
      RECT MASK 1 47.78 82.895 47.84 83.189 ;
      RECT MASK 1 48.444 82.895 48.504 83.189 ;
      RECT MASK 1 48.942 82.895 49.002 83.189 ;
      RECT MASK 1 49.606 82.895 49.666 83.189 ;
      RECT MASK 1 52.074 82.895 52.134 83.189 ;
      RECT MASK 1 52.738 82.895 52.798 83.189 ;
      RECT MASK 1 53.236 82.895 53.296 83.189 ;
      RECT MASK 1 53.9 82.895 53.96 83.189 ;
      RECT MASK 1 54.398 82.895 54.458 83.189 ;
      RECT MASK 1 55.062 82.895 55.122 83.189 ;
      RECT MASK 1 55.56 82.895 55.62 83.189 ;
      RECT MASK 1 56.224 82.895 56.284 83.189 ;
      RECT MASK 1 58.568 82.895 58.608 84.169 ;
      RECT MASK 1 58.692 82.895 58.752 83.189 ;
      RECT MASK 1 59.5 82.895 59.54 84.022 ;
      RECT MASK 1 59.73 82.895 59.77 84.022 ;
      RECT MASK 1 59.854 82.895 59.914 83.189 ;
      RECT MASK 1 61.016 82.895 61.076 83.189 ;
      RECT MASK 1 62.178 82.895 62.238 83.189 ;
      RECT MASK 1 65.31 82.895 65.37 83.189 ;
      RECT MASK 1 65.974 82.895 66.034 83.189 ;
      RECT MASK 1 66.472 82.895 66.532 83.189 ;
      RECT MASK 1 67.136 82.895 67.196 83.189 ;
      RECT MASK 1 67.634 82.895 67.694 83.189 ;
      RECT MASK 1 68.298 82.895 68.358 83.189 ;
      RECT MASK 1 68.796 82.895 68.856 83.189 ;
      RECT MASK 1 69.46 82.895 69.52 83.189 ;
      RECT MASK 1 71.928 82.895 71.988 83.189 ;
      RECT MASK 1 72.592 82.895 72.652 83.189 ;
      RECT MASK 1 73.09 82.895 73.15 83.189 ;
      RECT MASK 1 73.754 82.895 73.814 83.189 ;
      RECT MASK 1 74.252 82.895 74.312 83.189 ;
      RECT MASK 1 74.916 82.895 74.976 83.189 ;
      RECT MASK 1 75.414 82.895 75.474 83.189 ;
      RECT MASK 1 76.078 82.895 76.138 83.189 ;
      RECT MASK 1 78.546 82.895 78.606 83.189 ;
      RECT MASK 1 79.21 82.895 79.27 83.189 ;
      RECT MASK 1 79.708 82.895 79.768 83.189 ;
      RECT MASK 1 80.372 82.895 80.432 83.189 ;
      RECT MASK 1 80.87 82.895 80.93 83.189 ;
      RECT MASK 1 81.534 82.895 81.594 83.189 ;
      RECT MASK 1 82.032 82.895 82.092 83.189 ;
      RECT MASK 1 82.696 82.895 82.756 83.189 ;
      RECT MASK 1 85.164 82.895 85.224 83.189 ;
      RECT MASK 1 85.828 82.895 85.888 83.189 ;
      RECT MASK 1 86.326 82.895 86.386 83.189 ;
      RECT MASK 1 86.99 82.895 87.05 83.189 ;
      RECT MASK 1 87.488 82.895 87.548 83.189 ;
      RECT MASK 1 88.152 82.895 88.212 83.189 ;
      RECT MASK 1 88.65 82.895 88.71 83.189 ;
      RECT MASK 1 89.314 82.895 89.374 83.189 ;
      RECT MASK 1 91.782 82.895 91.842 83.189 ;
      RECT MASK 1 92.446 82.895 92.506 83.189 ;
      RECT MASK 1 92.944 82.895 93.004 83.189 ;
      RECT MASK 1 93.608 82.895 93.668 83.189 ;
      RECT MASK 1 94.106 82.895 94.166 83.189 ;
      RECT MASK 1 94.77 82.895 94.83 83.189 ;
      RECT MASK 1 95.268 82.895 95.328 83.189 ;
      RECT MASK 1 95.932 82.895 95.992 83.189 ;
      RECT MASK 1 98.4 82.895 98.46 83.189 ;
      RECT MASK 1 99.064 82.895 99.124 83.189 ;
      RECT MASK 1 99.562 82.895 99.622 83.189 ;
      RECT MASK 1 100.226 82.895 100.286 83.189 ;
      RECT MASK 1 100.724 82.895 100.784 83.189 ;
      RECT MASK 1 101.388 82.895 101.448 83.189 ;
      RECT MASK 1 101.886 82.895 101.946 83.189 ;
      RECT MASK 1 102.55 82.895 102.61 83.189 ;
      RECT MASK 1 105.018 82.895 105.078 83.189 ;
      RECT MASK 1 105.682 82.895 105.742 83.189 ;
      RECT MASK 1 106.18 82.895 106.24 83.189 ;
      RECT MASK 1 106.844 82.895 106.904 83.189 ;
      RECT MASK 1 107.342 82.895 107.402 83.189 ;
      RECT MASK 1 108.006 82.895 108.066 83.189 ;
      RECT MASK 1 108.504 82.895 108.564 83.189 ;
      RECT MASK 1 109.168 82.895 109.228 83.189 ;
      RECT MASK 1 6.91 83.309 6.97 85.141 ;
      RECT MASK 1 7.574 83.309 7.634 85.141 ;
      RECT MASK 1 8.072 83.309 8.132 85.141 ;
      RECT MASK 1 8.736 83.309 8.796 85.141 ;
      RECT MASK 1 9.234 83.309 9.294 85.141 ;
      RECT MASK 1 9.898 83.309 9.958 85.141 ;
      RECT MASK 1 12.366 83.309 12.426 85.141 ;
      RECT MASK 1 13.03 83.309 13.09 85.141 ;
      RECT MASK 1 13.528 83.309 13.588 85.141 ;
      RECT MASK 1 14.192 83.309 14.252 85.141 ;
      RECT MASK 1 14.69 83.309 14.75 85.141 ;
      RECT MASK 1 15.354 83.309 15.414 85.141 ;
      RECT MASK 1 15.852 83.309 15.912 85.141 ;
      RECT MASK 1 16.516 83.309 16.576 85.141 ;
      RECT MASK 1 18.984 83.309 19.044 85.141 ;
      RECT MASK 1 19.648 83.309 19.708 85.141 ;
      RECT MASK 1 20.146 83.309 20.206 85.141 ;
      RECT MASK 1 20.81 83.309 20.87 85.141 ;
      RECT MASK 1 21.308 83.309 21.368 85.141 ;
      RECT MASK 1 21.972 83.309 22.032 85.141 ;
      RECT MASK 1 22.47 83.309 22.53 85.141 ;
      RECT MASK 1 23.134 83.309 23.194 85.141 ;
      RECT MASK 1 25.602 83.309 25.662 85.141 ;
      RECT MASK 1 26.266 83.309 26.326 85.141 ;
      RECT MASK 1 26.764 83.309 26.824 85.141 ;
      RECT MASK 1 27.428 83.309 27.488 85.141 ;
      RECT MASK 1 27.926 83.309 27.986 85.141 ;
      RECT MASK 1 28.59 83.309 28.65 85.141 ;
      RECT MASK 1 29.088 83.309 29.148 85.141 ;
      RECT MASK 1 29.752 83.309 29.812 85.141 ;
      RECT MASK 1 32.22 83.309 32.28 85.141 ;
      RECT MASK 1 32.884 83.309 32.944 85.141 ;
      RECT MASK 1 33.382 83.309 33.442 85.141 ;
      RECT MASK 1 34.046 83.309 34.106 85.141 ;
      RECT MASK 1 34.544 83.309 34.604 85.141 ;
      RECT MASK 1 35.208 83.309 35.268 85.141 ;
      RECT MASK 1 35.706 83.309 35.766 85.141 ;
      RECT MASK 1 36.37 83.309 36.43 85.141 ;
      RECT MASK 1 38.838 83.309 38.898 85.141 ;
      RECT MASK 1 39.502 83.309 39.562 85.141 ;
      RECT MASK 1 40 83.309 40.06 85.141 ;
      RECT MASK 1 40.664 83.309 40.724 85.141 ;
      RECT MASK 1 41.162 83.309 41.222 85.141 ;
      RECT MASK 1 41.826 83.309 41.886 85.141 ;
      RECT MASK 1 42.324 83.309 42.384 85.141 ;
      RECT MASK 1 42.988 83.309 43.048 85.141 ;
      RECT MASK 1 45.456 83.309 45.516 85.141 ;
      RECT MASK 1 46.12 83.309 46.18 85.141 ;
      RECT MASK 1 46.618 83.309 46.678 85.141 ;
      RECT MASK 1 47.282 83.309 47.342 85.141 ;
      RECT MASK 1 47.78 83.309 47.84 85.141 ;
      RECT MASK 1 48.444 83.309 48.504 85.141 ;
      RECT MASK 1 48.942 83.309 49.002 85.141 ;
      RECT MASK 1 49.606 83.309 49.666 85.141 ;
      RECT MASK 1 52.074 83.309 52.134 85.141 ;
      RECT MASK 1 52.738 83.309 52.798 85.141 ;
      RECT MASK 1 53.236 83.309 53.296 85.141 ;
      RECT MASK 1 53.9 83.309 53.96 85.141 ;
      RECT MASK 1 54.398 83.309 54.458 85.141 ;
      RECT MASK 1 55.062 83.309 55.122 85.141 ;
      RECT MASK 1 55.56 83.309 55.62 85.141 ;
      RECT MASK 1 56.224 83.309 56.284 85.141 ;
      RECT MASK 1 58.692 83.309 58.752 85.141 ;
      RECT MASK 1 59.356 83.309 59.416 85.141 ;
      RECT MASK 1 59.854 83.309 59.914 85.141 ;
      RECT MASK 1 60.518 83.309 60.578 85.141 ;
      RECT MASK 1 61.016 83.309 61.076 85.141 ;
      RECT MASK 1 61.68 83.309 61.74 85.141 ;
      RECT MASK 1 62.178 83.309 62.238 85.141 ;
      RECT MASK 1 62.842 83.309 62.902 85.141 ;
      RECT MASK 1 65.31 83.309 65.37 85.141 ;
      RECT MASK 1 65.974 83.309 66.034 85.141 ;
      RECT MASK 1 66.472 83.309 66.532 85.141 ;
      RECT MASK 1 67.136 83.309 67.196 85.141 ;
      RECT MASK 1 67.634 83.309 67.694 85.141 ;
      RECT MASK 1 68.298 83.309 68.358 85.141 ;
      RECT MASK 1 68.796 83.309 68.856 85.141 ;
      RECT MASK 1 69.46 83.309 69.52 85.141 ;
      RECT MASK 1 71.928 83.309 71.988 85.141 ;
      RECT MASK 1 72.592 83.309 72.652 85.141 ;
      RECT MASK 1 73.09 83.309 73.15 85.141 ;
      RECT MASK 1 73.754 83.309 73.814 85.141 ;
      RECT MASK 1 74.252 83.309 74.312 85.141 ;
      RECT MASK 1 74.916 83.309 74.976 85.141 ;
      RECT MASK 1 75.414 83.309 75.474 85.141 ;
      RECT MASK 1 76.078 83.309 76.138 85.141 ;
      RECT MASK 1 78.546 83.309 78.606 85.141 ;
      RECT MASK 1 79.21 83.309 79.27 85.141 ;
      RECT MASK 1 79.708 83.309 79.768 85.141 ;
      RECT MASK 1 80.372 83.309 80.432 85.141 ;
      RECT MASK 1 80.87 83.309 80.93 85.141 ;
      RECT MASK 1 81.534 83.309 81.594 85.141 ;
      RECT MASK 1 82.032 83.309 82.092 85.141 ;
      RECT MASK 1 82.696 83.309 82.756 85.141 ;
      RECT MASK 1 85.164 83.309 85.224 85.141 ;
      RECT MASK 1 85.828 83.309 85.888 85.141 ;
      RECT MASK 1 86.326 83.309 86.386 85.141 ;
      RECT MASK 1 86.99 83.309 87.05 85.141 ;
      RECT MASK 1 87.488 83.309 87.548 85.141 ;
      RECT MASK 1 88.152 83.309 88.212 85.141 ;
      RECT MASK 1 88.65 83.309 88.71 85.141 ;
      RECT MASK 1 89.314 83.309 89.374 85.141 ;
      RECT MASK 1 91.782 83.309 91.842 85.141 ;
      RECT MASK 1 92.446 83.309 92.506 85.141 ;
      RECT MASK 1 92.944 83.309 93.004 85.141 ;
      RECT MASK 1 93.608 83.309 93.668 85.141 ;
      RECT MASK 1 94.106 83.309 94.166 85.141 ;
      RECT MASK 1 94.77 83.309 94.83 85.141 ;
      RECT MASK 1 95.268 83.309 95.328 85.141 ;
      RECT MASK 1 95.932 83.309 95.992 85.141 ;
      RECT MASK 1 98.4 83.309 98.46 85.141 ;
      RECT MASK 1 99.064 83.309 99.124 85.141 ;
      RECT MASK 1 99.562 83.309 99.622 85.141 ;
      RECT MASK 1 100.226 83.309 100.286 85.141 ;
      RECT MASK 1 100.724 83.309 100.784 85.141 ;
      RECT MASK 1 101.388 83.309 101.448 85.141 ;
      RECT MASK 1 101.886 83.309 101.946 85.141 ;
      RECT MASK 1 102.55 83.309 102.61 85.141 ;
      RECT MASK 1 105.018 83.309 105.078 85.141 ;
      RECT MASK 1 105.682 83.309 105.742 85.141 ;
      RECT MASK 1 106.18 83.309 106.24 85.141 ;
      RECT MASK 1 106.844 83.309 106.904 85.141 ;
      RECT MASK 1 107.342 83.309 107.402 85.141 ;
      RECT MASK 1 108.006 83.309 108.066 85.141 ;
      RECT MASK 1 108.504 83.309 108.564 85.141 ;
      RECT MASK 1 109.168 83.309 109.228 85.141 ;
      RECT MASK 1 6.329 84.308 6.389 86.056 ;
      RECT MASK 1 10.479 84.308 10.539 86.056 ;
      RECT MASK 1 11.049 84.308 11.109 86.0585 ;
      RECT MASK 1 11.381 84.308 11.441 86.0585 ;
      RECT MASK 1 11.785 84.308 11.845 86.056 ;
      RECT MASK 1 17.097 84.308 17.157 86.056 ;
      RECT MASK 1 17.667 84.308 17.727 86.0585 ;
      RECT MASK 1 17.999 84.308 18.059 86.0585 ;
      RECT MASK 1 18.403 84.308 18.463 86.056 ;
      RECT MASK 1 23.715 84.308 23.775 86.056 ;
      RECT MASK 1 24.285 84.308 24.345 86.0585 ;
      RECT MASK 1 24.617 84.308 24.677 86.0585 ;
      RECT MASK 1 25.021 84.308 25.081 86.056 ;
      RECT MASK 1 30.333 84.308 30.393 86.056 ;
      RECT MASK 1 30.903 84.308 30.963 86.0585 ;
      RECT MASK 1 31.235 84.308 31.295 86.0585 ;
      RECT MASK 1 31.639 84.308 31.699 86.056 ;
      RECT MASK 1 36.951 84.308 37.011 86.056 ;
      RECT MASK 1 37.521 84.308 37.581 86.0585 ;
      RECT MASK 1 37.853 84.308 37.913 86.0585 ;
      RECT MASK 1 38.257 84.308 38.317 86.056 ;
      RECT MASK 1 43.569 84.308 43.629 86.056 ;
      RECT MASK 1 44.139 84.308 44.199 86.0585 ;
      RECT MASK 1 44.471 84.308 44.531 86.0585 ;
      RECT MASK 1 44.875 84.308 44.935 86.056 ;
      RECT MASK 1 50.187 84.308 50.247 86.056 ;
      RECT MASK 1 50.757 84.308 50.817 86.0585 ;
      RECT MASK 1 51.089 84.308 51.149 86.0585 ;
      RECT MASK 1 51.493 84.308 51.553 86.056 ;
      RECT MASK 1 56.805 84.308 56.865 86.056 ;
      RECT MASK 1 57.375 84.308 57.435 86.0585 ;
      RECT MASK 1 57.707 84.308 57.767 86.0585 ;
      RECT MASK 1 58.111 84.308 58.171 86.056 ;
      RECT MASK 1 63.423 84.308 63.483 86.056 ;
      RECT MASK 1 63.993 84.308 64.053 86.0585 ;
      RECT MASK 1 64.325 84.308 64.385 86.0585 ;
      RECT MASK 1 64.729 84.308 64.789 86.056 ;
      RECT MASK 1 70.041 84.308 70.101 86.056 ;
      RECT MASK 1 70.611 84.308 70.671 86.0585 ;
      RECT MASK 1 70.943 84.308 71.003 86.0585 ;
      RECT MASK 1 71.347 84.308 71.407 86.056 ;
      RECT MASK 1 76.659 84.308 76.719 86.056 ;
      RECT MASK 1 77.229 84.308 77.289 86.0585 ;
      RECT MASK 1 77.561 84.308 77.621 86.0585 ;
      RECT MASK 1 77.965 84.308 78.025 86.056 ;
      RECT MASK 1 83.277 84.308 83.337 86.056 ;
      RECT MASK 1 83.847 84.308 83.907 86.0585 ;
      RECT MASK 1 84.179 84.308 84.239 86.0585 ;
      RECT MASK 1 84.583 84.308 84.643 86.056 ;
      RECT MASK 1 89.895 84.308 89.955 86.056 ;
      RECT MASK 1 90.465 84.308 90.525 86.0585 ;
      RECT MASK 1 90.797 84.308 90.857 86.0585 ;
      RECT MASK 1 91.201 84.308 91.261 86.056 ;
      RECT MASK 1 96.513 84.308 96.573 86.056 ;
      RECT MASK 1 97.083 84.308 97.143 86.0585 ;
      RECT MASK 1 97.415 84.308 97.475 86.0585 ;
      RECT MASK 1 97.819 84.308 97.879 86.056 ;
      RECT MASK 1 103.131 84.308 103.191 86.056 ;
      RECT MASK 1 103.701 84.308 103.761 86.0585 ;
      RECT MASK 1 104.033 84.308 104.093 86.0585 ;
      RECT MASK 1 104.437 84.308 104.497 86.056 ;
      RECT MASK 1 109.749 84.308 109.809 86.056 ;
      RECT MASK 1 6.91 85.261 6.97 86.056 ;
      RECT MASK 1 7.574 85.261 7.634 86.056 ;
      RECT MASK 1 8.072 85.261 8.132 86.056 ;
      RECT MASK 1 8.736 85.261 8.796 86.055 ;
      RECT MASK 1 9.234 85.261 9.294 86.056 ;
      RECT MASK 1 9.898 85.261 9.958 86.056 ;
      RECT MASK 1 12.366 85.261 12.426 86.056 ;
      RECT MASK 1 13.03 85.261 13.09 86.056 ;
      RECT MASK 1 13.528 85.261 13.588 86.056 ;
      RECT MASK 1 14.192 85.261 14.252 86.056 ;
      RECT MASK 1 14.69 85.261 14.75 86.056 ;
      RECT MASK 1 15.354 85.261 15.414 86.055 ;
      RECT MASK 1 15.852 85.261 15.912 86.056 ;
      RECT MASK 1 16.516 85.261 16.576 86.056 ;
      RECT MASK 1 18.984 85.261 19.044 86.056 ;
      RECT MASK 1 19.648 85.261 19.708 86.056 ;
      RECT MASK 1 20.146 85.261 20.206 86.056 ;
      RECT MASK 1 20.81 85.261 20.87 86.056 ;
      RECT MASK 1 21.308 85.261 21.368 86.056 ;
      RECT MASK 1 21.972 85.261 22.032 86.055 ;
      RECT MASK 1 22.47 85.261 22.53 86.056 ;
      RECT MASK 1 23.134 85.261 23.194 86.056 ;
      RECT MASK 1 25.602 85.261 25.662 86.056 ;
      RECT MASK 1 26.266 85.261 26.326 86.056 ;
      RECT MASK 1 26.764 85.261 26.824 86.056 ;
      RECT MASK 1 27.428 85.261 27.488 86.056 ;
      RECT MASK 1 27.926 85.261 27.986 86.056 ;
      RECT MASK 1 28.59 85.261 28.65 86.055 ;
      RECT MASK 1 29.088 85.261 29.148 86.056 ;
      RECT MASK 1 29.752 85.261 29.812 86.056 ;
      RECT MASK 1 32.22 85.261 32.28 86.056 ;
      RECT MASK 1 32.884 85.261 32.944 86.056 ;
      RECT MASK 1 33.382 85.261 33.442 86.056 ;
      RECT MASK 1 34.046 85.261 34.106 86.056 ;
      RECT MASK 1 34.544 85.261 34.604 86.056 ;
      RECT MASK 1 35.208 85.261 35.268 86.055 ;
      RECT MASK 1 35.706 85.261 35.766 86.056 ;
      RECT MASK 1 36.37 85.261 36.43 86.056 ;
      RECT MASK 1 38.838 85.261 38.898 86.056 ;
      RECT MASK 1 39.502 85.261 39.562 86.056 ;
      RECT MASK 1 40 85.261 40.06 86.056 ;
      RECT MASK 1 40.664 85.261 40.724 86.056 ;
      RECT MASK 1 41.162 85.261 41.222 86.056 ;
      RECT MASK 1 41.826 85.261 41.886 86.055 ;
      RECT MASK 1 42.324 85.261 42.384 86.056 ;
      RECT MASK 1 42.988 85.261 43.048 86.056 ;
      RECT MASK 1 45.456 85.261 45.516 86.056 ;
      RECT MASK 1 46.12 85.261 46.18 86.056 ;
      RECT MASK 1 46.618 85.261 46.678 86.056 ;
      RECT MASK 1 47.282 85.261 47.342 86.056 ;
      RECT MASK 1 47.78 85.261 47.84 86.056 ;
      RECT MASK 1 48.444 85.261 48.504 86.055 ;
      RECT MASK 1 48.942 85.261 49.002 86.056 ;
      RECT MASK 1 49.606 85.261 49.666 86.056 ;
      RECT MASK 1 52.074 85.261 52.134 86.056 ;
      RECT MASK 1 52.738 85.261 52.798 86.056 ;
      RECT MASK 1 53.236 85.261 53.296 86.056 ;
      RECT MASK 1 53.9 85.261 53.96 86.056 ;
      RECT MASK 1 54.398 85.261 54.458 86.056 ;
      RECT MASK 1 55.062 85.261 55.122 86.055 ;
      RECT MASK 1 55.56 85.261 55.62 86.056 ;
      RECT MASK 1 56.224 85.261 56.284 86.056 ;
      RECT MASK 1 58.692 85.261 58.752 86.056 ;
      RECT MASK 1 59.356 85.261 59.416 86.056 ;
      RECT MASK 1 59.854 85.261 59.914 86.056 ;
      RECT MASK 1 60.518 85.261 60.578 86.056 ;
      RECT MASK 1 61.016 85.261 61.076 86.056 ;
      RECT MASK 1 61.68 85.261 61.74 86.055 ;
      RECT MASK 1 62.178 85.261 62.238 86.056 ;
      RECT MASK 1 62.842 85.261 62.902 86.056 ;
      RECT MASK 1 65.31 85.261 65.37 86.056 ;
      RECT MASK 1 65.974 85.261 66.034 86.056 ;
      RECT MASK 1 66.472 85.261 66.532 86.056 ;
      RECT MASK 1 67.136 85.261 67.196 86.056 ;
      RECT MASK 1 67.634 85.261 67.694 86.056 ;
      RECT MASK 1 68.298 85.261 68.358 86.055 ;
      RECT MASK 1 68.796 85.261 68.856 86.056 ;
      RECT MASK 1 69.46 85.261 69.52 86.056 ;
      RECT MASK 1 71.928 85.261 71.988 86.056 ;
      RECT MASK 1 72.592 85.261 72.652 86.056 ;
      RECT MASK 1 73.09 85.261 73.15 86.056 ;
      RECT MASK 1 73.754 85.261 73.814 86.056 ;
      RECT MASK 1 74.252 85.261 74.312 86.056 ;
      RECT MASK 1 74.916 85.261 74.976 86.055 ;
      RECT MASK 1 75.414 85.261 75.474 86.056 ;
      RECT MASK 1 76.078 85.261 76.138 86.056 ;
      RECT MASK 1 78.546 85.261 78.606 86.056 ;
      RECT MASK 1 79.21 85.261 79.27 86.056 ;
      RECT MASK 1 79.708 85.261 79.768 86.056 ;
      RECT MASK 1 80.372 85.261 80.432 86.056 ;
      RECT MASK 1 80.87 85.261 80.93 86.056 ;
      RECT MASK 1 81.534 85.261 81.594 86.055 ;
      RECT MASK 1 82.032 85.261 82.092 86.056 ;
      RECT MASK 1 82.696 85.261 82.756 86.056 ;
      RECT MASK 1 85.164 85.261 85.224 86.056 ;
      RECT MASK 1 85.828 85.261 85.888 86.056 ;
      RECT MASK 1 86.326 85.261 86.386 86.056 ;
      RECT MASK 1 86.99 85.261 87.05 86.056 ;
      RECT MASK 1 87.488 85.261 87.548 86.056 ;
      RECT MASK 1 88.152 85.261 88.212 86.055 ;
      RECT MASK 1 88.65 85.261 88.71 86.056 ;
      RECT MASK 1 89.314 85.261 89.374 86.056 ;
      RECT MASK 1 91.782 85.261 91.842 86.056 ;
      RECT MASK 1 92.446 85.261 92.506 86.056 ;
      RECT MASK 1 92.944 85.261 93.004 86.056 ;
      RECT MASK 1 93.608 85.261 93.668 86.056 ;
      RECT MASK 1 94.106 85.261 94.166 86.056 ;
      RECT MASK 1 94.77 85.261 94.83 86.055 ;
      RECT MASK 1 95.268 85.261 95.328 86.056 ;
      RECT MASK 1 95.932 85.261 95.992 86.056 ;
      RECT MASK 1 98.4 85.261 98.46 86.056 ;
      RECT MASK 1 99.064 85.261 99.124 86.056 ;
      RECT MASK 1 99.562 85.261 99.622 86.056 ;
      RECT MASK 1 100.226 85.261 100.286 86.056 ;
      RECT MASK 1 100.724 85.261 100.784 86.056 ;
      RECT MASK 1 101.388 85.261 101.448 86.055 ;
      RECT MASK 1 101.886 85.261 101.946 86.056 ;
      RECT MASK 1 102.55 85.261 102.61 86.056 ;
      RECT MASK 1 105.018 85.261 105.078 86.056 ;
      RECT MASK 1 105.682 85.261 105.742 86.056 ;
      RECT MASK 1 106.18 85.261 106.24 86.056 ;
      RECT MASK 1 106.844 85.261 106.904 86.056 ;
      RECT MASK 1 107.342 85.261 107.402 86.056 ;
      RECT MASK 1 108.006 85.261 108.066 86.055 ;
      RECT MASK 1 108.504 85.261 108.564 86.056 ;
      RECT MASK 1 109.168 85.261 109.228 86.056 ;
      RECT MASK 1 22.218 85.4905 22.278 86.055 ;
      RECT MASK 1 28.836 85.4905 28.896 86.055 ;
      RECT MASK 1 35.454 85.4905 35.514 86.055 ;
      RECT MASK 1 42.072 85.4905 42.132 86.055 ;
      RECT MASK 1 48.69 85.4905 48.75 86.055 ;
      RECT MASK 1 55.308 85.4905 55.368 86.055 ;
      RECT MASK 1 61.926 85.4905 61.986 86.055 ;
      RECT MASK 1 68.544 85.4905 68.604 86.055 ;
      RECT MASK 1 75.162 85.4905 75.222 86.055 ;
      RECT MASK 1 81.78 85.4905 81.84 86.055 ;
      RECT MASK 1 88.398 85.4905 88.458 86.055 ;
      RECT MASK 1 95.016 85.4905 95.076 86.055 ;
      RECT MASK 1 101.634 85.4905 101.694 86.055 ;
      RECT MASK 1 108.252 85.4905 108.312 86.055 ;
      RECT MASK 1 20.478 85.4915 20.538 86.056 ;
      RECT MASK 1 21.056 85.4915 21.116 86.056 ;
      RECT MASK 1 21.64 85.4915 21.7 86.056 ;
      RECT MASK 1 22.802 85.4915 22.862 86.056 ;
      RECT MASK 1 23.434 85.4915 23.494 86.056 ;
      RECT MASK 1 27.096 85.4915 27.156 86.056 ;
      RECT MASK 1 27.674 85.4915 27.734 86.056 ;
      RECT MASK 1 28.258 85.4915 28.318 86.056 ;
      RECT MASK 1 29.42 85.4915 29.48 86.056 ;
      RECT MASK 1 30.052 85.4915 30.112 86.056 ;
      RECT MASK 1 33.714 85.4915 33.774 86.056 ;
      RECT MASK 1 34.292 85.4915 34.352 86.056 ;
      RECT MASK 1 34.876 85.4915 34.936 86.056 ;
      RECT MASK 1 36.038 85.4915 36.098 86.056 ;
      RECT MASK 1 36.67 85.4915 36.73 86.056 ;
      RECT MASK 1 40.332 85.4915 40.392 86.056 ;
      RECT MASK 1 40.91 85.4915 40.97 86.056 ;
      RECT MASK 1 41.494 85.4915 41.554 86.056 ;
      RECT MASK 1 42.656 85.4915 42.716 86.056 ;
      RECT MASK 1 43.288 85.4915 43.348 86.056 ;
      RECT MASK 1 46.95 85.4915 47.01 86.056 ;
      RECT MASK 1 47.528 85.4915 47.588 86.056 ;
      RECT MASK 1 48.112 85.4915 48.172 86.056 ;
      RECT MASK 1 49.274 85.4915 49.334 86.056 ;
      RECT MASK 1 49.906 85.4915 49.966 86.056 ;
      RECT MASK 1 53.568 85.4915 53.628 86.056 ;
      RECT MASK 1 54.146 85.4915 54.206 86.056 ;
      RECT MASK 1 54.73 85.4915 54.79 86.056 ;
      RECT MASK 1 55.892 85.4915 55.952 86.056 ;
      RECT MASK 1 56.524 85.4915 56.584 86.056 ;
      RECT MASK 1 60.186 85.4915 60.246 86.056 ;
      RECT MASK 1 60.764 85.4915 60.824 86.056 ;
      RECT MASK 1 61.348 85.4915 61.408 86.056 ;
      RECT MASK 1 62.51 85.4915 62.57 86.056 ;
      RECT MASK 1 63.142 85.4915 63.202 86.056 ;
      RECT MASK 1 66.804 85.4915 66.864 86.056 ;
      RECT MASK 1 67.382 85.4915 67.442 86.056 ;
      RECT MASK 1 67.966 85.4915 68.026 86.056 ;
      RECT MASK 1 69.128 85.4915 69.188 86.056 ;
      RECT MASK 1 69.76 85.4915 69.82 86.056 ;
      RECT MASK 1 73.422 85.4915 73.482 86.056 ;
      RECT MASK 1 74 85.4915 74.06 86.056 ;
      RECT MASK 1 74.584 85.4915 74.644 86.056 ;
      RECT MASK 1 75.746 85.4915 75.806 86.056 ;
      RECT MASK 1 76.378 85.4915 76.438 86.056 ;
      RECT MASK 1 80.04 85.4915 80.1 86.056 ;
      RECT MASK 1 80.618 85.4915 80.678 86.056 ;
      RECT MASK 1 81.202 85.4915 81.262 86.056 ;
      RECT MASK 1 82.364 85.4915 82.424 86.056 ;
      RECT MASK 1 82.996 85.4915 83.056 86.056 ;
      RECT MASK 1 86.658 85.4915 86.718 86.056 ;
      RECT MASK 1 87.236 85.4915 87.296 86.056 ;
      RECT MASK 1 87.82 85.4915 87.88 86.056 ;
      RECT MASK 1 88.982 85.4915 89.042 86.056 ;
      RECT MASK 1 89.614 85.4915 89.674 86.056 ;
      RECT MASK 1 93.276 85.4915 93.336 86.056 ;
      RECT MASK 1 93.854 85.4915 93.914 86.056 ;
      RECT MASK 1 94.438 85.4915 94.498 86.056 ;
      RECT MASK 1 95.6 85.4915 95.66 86.056 ;
      RECT MASK 1 96.232 85.4915 96.292 86.056 ;
      RECT MASK 1 99.894 85.4915 99.954 86.056 ;
      RECT MASK 1 100.472 85.4915 100.532 86.056 ;
      RECT MASK 1 101.056 85.4915 101.116 86.056 ;
      RECT MASK 1 102.218 85.4915 102.278 86.056 ;
      RECT MASK 1 102.85 85.4915 102.91 86.056 ;
      RECT MASK 1 106.512 85.4915 106.572 86.056 ;
      RECT MASK 1 107.09 85.4915 107.15 86.056 ;
      RECT MASK 1 107.674 85.4915 107.734 86.056 ;
      RECT MASK 1 108.836 85.4915 108.896 86.056 ;
      RECT MASK 1 109.468 85.4915 109.528 86.056 ;
      RECT MASK 1 18.6935 85.5 18.7535 86.056 ;
      RECT MASK 1 19.316 85.5 19.376 86.056 ;
      RECT MASK 1 25.3115 85.5 25.3715 86.056 ;
      RECT MASK 1 25.934 85.5 25.994 86.056 ;
      RECT MASK 1 31.9295 85.5 31.9895 86.056 ;
      RECT MASK 1 32.552 85.5 32.612 86.056 ;
      RECT MASK 1 38.5475 85.5 38.6075 86.056 ;
      RECT MASK 1 39.17 85.5 39.23 86.056 ;
      RECT MASK 1 45.1655 85.5 45.2255 86.056 ;
      RECT MASK 1 45.788 85.5 45.848 86.056 ;
      RECT MASK 1 51.7835 85.5 51.8435 86.056 ;
      RECT MASK 1 52.406 85.5 52.466 86.056 ;
      RECT MASK 1 58.4015 85.5 58.4615 86.056 ;
      RECT MASK 1 59.024 85.5 59.084 86.056 ;
      RECT MASK 1 65.0195 85.5 65.0795 86.056 ;
      RECT MASK 1 65.642 85.5 65.702 86.056 ;
      RECT MASK 1 71.6375 85.5 71.6975 86.056 ;
      RECT MASK 1 72.26 85.5 72.32 86.056 ;
      RECT MASK 1 78.2555 85.5 78.3155 86.056 ;
      RECT MASK 1 78.878 85.5 78.938 86.056 ;
      RECT MASK 1 84.8735 85.5 84.9335 86.056 ;
      RECT MASK 1 85.496 85.5 85.556 86.056 ;
      RECT MASK 1 91.4915 85.5 91.5515 86.056 ;
      RECT MASK 1 92.114 85.5 92.174 86.056 ;
      RECT MASK 1 98.1095 85.5 98.1695 86.056 ;
      RECT MASK 1 98.732 85.5 98.792 86.056 ;
      RECT MASK 1 104.7275 85.5 104.7875 86.056 ;
      RECT MASK 1 105.35 85.5 105.41 86.056 ;
      RECT MASK 1 72.062 86.242 72.202 95.438 ;
      RECT MASK 1 103.38 86.242 103.52 95.438 ;
      RECT MASK 1 69.9 86.255 69.96 86.515 ;
      RECT MASK 1 70.149 86.255 70.209 86.515 ;
      RECT MASK 1 70.398 86.255 70.458 86.965 ;
      RECT MASK 1 70.647 86.255 70.707 86.965 ;
      RECT MASK 1 70.896 86.255 70.956 86.965 ;
      RECT MASK 1 71.145 86.255 71.205 86.965 ;
      RECT MASK 1 71.394 86.255 71.454 86.965 ;
      RECT MASK 1 71.643 86.255 71.703 86.965 ;
      RECT MASK 1 103.879 86.255 103.939 86.965 ;
      RECT MASK 1 104.128 86.255 104.188 86.965 ;
      RECT MASK 1 104.377 86.255 104.437 86.965 ;
      RECT MASK 1 104.626 86.255 104.686 86.965 ;
      RECT MASK 1 104.875 86.255 104.935 86.965 ;
      RECT MASK 1 105.124 86.255 105.184 86.965 ;
      RECT MASK 1 105.373 86.255 105.433 86.515 ;
      RECT MASK 1 105.622 86.255 105.682 86.515 ;
      RECT MASK 1 33.51 86.345 33.57 86.605 ;
      RECT MASK 1 33.759 86.345 33.819 86.605 ;
      RECT MASK 1 34.008 86.345 34.068 87.055 ;
      RECT MASK 1 34.257 86.345 34.317 87.055 ;
      RECT MASK 1 34.506 86.345 34.566 87.055 ;
      RECT MASK 1 34.755 86.345 34.815 87.055 ;
      RECT MASK 1 35.004 86.345 35.064 87.055 ;
      RECT MASK 1 35.253 86.345 35.313 87.055 ;
      RECT MASK 1 67.572 86.345 67.632 87.055 ;
      RECT MASK 1 67.821 86.345 67.881 87.055 ;
      RECT MASK 1 68.07 86.345 68.13 87.055 ;
      RECT MASK 1 68.319 86.345 68.379 87.055 ;
      RECT MASK 1 68.568 86.345 68.628 87.055 ;
      RECT MASK 1 68.817 86.345 68.877 86.605 ;
      RECT MASK 1 69.066 86.345 69.126 86.605 ;
      RECT MASK 1 35.672 86.35 35.812 95.33 ;
      RECT MASK 1 66.99 86.35 67.13 95.33 ;
      RECT MASK 1 36.1535 86.469 66.6485 86.569 ;
      RECT MASK 1 72.5435 86.469 103.0385 86.569 ;
      RECT MASK 1 69.797 86.6735 69.897 95.0065 ;
      RECT MASK 1 105.685 86.6735 105.785 95.0065 ;
      RECT MASK 1 33.407 86.7635 33.507 94.9165 ;
      RECT MASK 1 69.129 86.7635 69.229 94.9165 ;
      RECT MASK 1 70.129 87.1235 70.229 94.5565 ;
      RECT MASK 1 105.353 87.1235 105.453 94.5565 ;
      RECT MASK 1 36.326 87.147 66.476 87.207 ;
      RECT MASK 1 72.716 87.147 102.866 87.207 ;
      RECT MASK 1 17.061 87.19 17.161 94.37 ;
      RECT MASK 1 8.195 87.201 8.295 90.966 ;
      RECT MASK 1 12.677 87.201 12.777 94.359 ;
      RECT MASK 1 17.627 87.201 17.727 94.359 ;
      RECT MASK 1 22.109 87.201 22.209 94.359 ;
      RECT MASK 1 8.547 87.21 8.607 87.49 ;
      RECT MASK 1 8.879 87.21 8.939 87.49 ;
      RECT MASK 1 9.211 87.21 9.271 87.49 ;
      RECT MASK 1 9.543 87.21 9.603 87.49 ;
      RECT MASK 1 9.875 87.21 9.935 87.49 ;
      RECT MASK 1 10.207 87.21 10.267 87.49 ;
      RECT MASK 1 10.539 87.21 10.599 87.49 ;
      RECT MASK 1 10.871 87.21 10.931 87.49 ;
      RECT MASK 1 11.203 87.21 11.263 87.49 ;
      RECT MASK 1 11.535 87.21 11.595 87.49 ;
      RECT MASK 1 11.867 87.21 11.927 87.49 ;
      RECT MASK 1 12.199 87.21 12.259 87.49 ;
      RECT MASK 1 13.595 87.21 13.655 87.49 ;
      RECT MASK 1 13.927 87.21 13.987 87.49 ;
      RECT MASK 1 14.259 87.21 14.319 87.49 ;
      RECT MASK 1 14.757 87.21 14.817 87.49 ;
      RECT MASK 1 15.089 87.21 15.149 87.49 ;
      RECT MASK 1 15.421 87.21 15.481 87.49 ;
      RECT MASK 1 15.753 87.21 15.813 87.49 ;
      RECT MASK 1 16.085 87.21 16.145 87.49 ;
      RECT MASK 1 16.417 87.21 16.477 87.49 ;
      RECT MASK 1 16.749 87.21 16.809 87.49 ;
      RECT MASK 1 18.145 87.21 18.205 87.49 ;
      RECT MASK 1 18.477 87.21 18.537 87.49 ;
      RECT MASK 1 18.809 87.21 18.869 87.49 ;
      RECT MASK 1 19.141 87.21 19.201 87.49 ;
      RECT MASK 1 19.473 87.21 19.533 87.49 ;
      RECT MASK 1 19.805 87.21 19.865 87.49 ;
      RECT MASK 1 20.137 87.21 20.197 87.49 ;
      RECT MASK 1 20.469 87.21 20.529 87.49 ;
      RECT MASK 1 20.801 87.21 20.861 87.49 ;
      RECT MASK 1 21.133 87.21 21.193 87.49 ;
      RECT MASK 1 21.465 87.21 21.525 87.49 ;
      RECT MASK 1 21.797 87.21 21.857 87.49 ;
      RECT MASK 1 33.739 87.2135 33.839 94.4665 ;
      RECT MASK 1 68.797 87.2135 68.897 94.4665 ;
      RECT MASK 1 6.009 87.215 6.069 88.942 ;
      RECT MASK 1 7.005 87.215 7.065 88.942 ;
      RECT MASK 1 107.494 87.23 107.594 97.101 ;
      RECT MASK 1 25.66 87.237 30.63 87.297 ;
      RECT MASK 1 34.365 87.3 34.465 94.38 ;
      RECT MASK 1 34.697 87.3 34.797 94.38 ;
      RECT MASK 1 35.029 87.3 35.129 94.38 ;
      RECT MASK 1 67.839 87.3 67.939 94.38 ;
      RECT MASK 1 68.171 87.3 68.271 94.38 ;
      RECT MASK 1 70.755 87.3 70.855 94.38 ;
      RECT MASK 1 71.087 87.3 71.187 94.38 ;
      RECT MASK 1 71.419 87.3 71.519 94.38 ;
      RECT MASK 1 104.063 87.3 104.163 94.38 ;
      RECT MASK 1 104.395 87.3 104.495 94.38 ;
      RECT MASK 1 104.727 87.3 104.827 94.38 ;
      RECT MASK 1 36.326 87.399 66.476 87.459 ;
      RECT MASK 1 72.716 87.399 102.866 87.459 ;
      RECT MASK 1 8.7785 87.66 8.8785 90.24 ;
      RECT MASK 1 9.1305 87.66 9.1905 88.912 ;
      RECT MASK 1 9.4625 87.66 9.5225 88.912 ;
      RECT MASK 1 9.7945 87.66 9.8545 88.912 ;
      RECT MASK 1 10.1265 87.66 10.1865 88.912 ;
      RECT MASK 1 10.4585 87.66 10.5185 88.912 ;
      RECT MASK 1 10.7905 87.66 10.8505 88.912 ;
      RECT MASK 1 11.1225 87.66 11.1825 88.912 ;
      RECT MASK 1 11.4545 87.66 11.5145 88.912 ;
      RECT MASK 1 11.7865 87.66 11.8465 88.912 ;
      RECT MASK 1 13.8265 87.66 13.9265 90.24 ;
      RECT MASK 1 14.1585 87.66 14.2585 88.39 ;
      RECT MASK 1 14.4905 87.66 14.5905 88.39 ;
      RECT MASK 1 14.8225 87.66 14.9225 88.39 ;
      RECT MASK 1 15.1545 87.66 15.2545 88.39 ;
      RECT MASK 1 15.4865 87.66 15.5865 88.39 ;
      RECT MASK 1 15.8185 87.66 15.9185 88.39 ;
      RECT MASK 1 16.1505 87.66 16.2505 88.39 ;
      RECT MASK 1 16.4825 87.66 16.5825 90.24 ;
      RECT MASK 1 18.2105 87.66 18.3105 90.24 ;
      RECT MASK 1 18.7285 87.66 18.7885 88.912 ;
      RECT MASK 1 21.0525 87.66 21.1125 88.912 ;
      RECT MASK 1 21.5305 87.66 21.6305 90.24 ;
      RECT MASK 1 6.424 87.72 6.484 87.989 ;
      RECT MASK 1 108.242 87.72 108.302 96.66 ;
      RECT MASK 1 108.516 87.72 108.576 96.66 ;
      RECT MASK 1 108.79 87.72 108.85 96.66 ;
      RECT MASK 1 109.064 87.72 109.124 96.66 ;
      RECT MASK 1 109.338 87.72 109.398 96.66 ;
      RECT MASK 1 109.612 87.72 109.672 96.66 ;
      RECT MASK 1 109.886 87.72 109.946 96.66 ;
      RECT MASK 1 110.16 87.72 110.22 96.66 ;
      RECT MASK 1 110.434 87.72 110.494 96.66 ;
      RECT MASK 1 110.708 87.72 110.768 96.66 ;
      RECT MASK 1 110.982 87.72 111.042 96.66 ;
      RECT MASK 1 111.256 87.72 111.316 96.66 ;
      RECT MASK 1 111.53 87.72 111.59 96.66 ;
      RECT MASK 1 111.804 87.72 111.864 96.66 ;
      RECT MASK 1 112.078 87.72 112.138 96.66 ;
      RECT MASK 1 112.352 87.72 112.412 96.66 ;
      RECT MASK 1 112.626 87.72 112.686 96.66 ;
      RECT MASK 1 112.9 87.72 112.96 96.66 ;
      RECT MASK 1 113.174 87.72 113.234 96.66 ;
      RECT MASK 1 113.448 87.72 113.508 96.66 ;
      RECT MASK 1 113.722 87.72 113.782 96.66 ;
      RECT MASK 1 113.996 87.72 114.056 96.66 ;
      RECT MASK 1 114.27 87.72 114.33 96.66 ;
      RECT MASK 1 114.544 87.72 114.604 96.66 ;
      RECT MASK 1 114.818 87.72 114.878 96.66 ;
      RECT MASK 1 115.092 87.72 115.152 96.66 ;
      RECT MASK 1 115.366 87.72 115.426 96.66 ;
      RECT MASK 1 115.64 87.72 115.7 96.66 ;
      RECT MASK 1 115.914 87.72 115.974 96.66 ;
      RECT MASK 1 116.188 87.72 116.248 96.66 ;
      RECT MASK 1 116.462 87.72 116.522 96.66 ;
      RECT MASK 1 127.696 87.72 127.756 96.66 ;
      RECT MASK 1 25.66 87.821 25.945 87.881 ;
      RECT MASK 1 26.204 87.821 30.086 87.881 ;
      RECT MASK 1 30.345 87.821 30.63 87.881 ;
      RECT MASK 1 36.326 88.047 36.778 88.107 ;
      RECT MASK 1 37.048 88.047 65.754 88.107 ;
      RECT MASK 1 66.024 88.047 66.476 88.107 ;
      RECT MASK 1 72.716 88.047 73.168 88.107 ;
      RECT MASK 1 73.438 88.047 102.144 88.107 ;
      RECT MASK 1 102.414 88.047 102.866 88.107 ;
      RECT MASK 1 25.66 88.083 25.944 88.143 ;
      RECT MASK 1 26.205 88.083 30.085 88.143 ;
      RECT MASK 1 30.346 88.083 30.63 88.143 ;
      RECT MASK 1 6.424 88.109 6.484 90.041 ;
      RECT MASK 1 36.326 88.299 36.778 88.359 ;
      RECT MASK 1 37.048 88.299 65.754 88.359 ;
      RECT MASK 1 66.024 88.299 66.476 88.359 ;
      RECT MASK 1 72.716 88.299 73.168 88.359 ;
      RECT MASK 1 73.438 88.299 102.144 88.359 ;
      RECT MASK 1 102.414 88.299 102.866 88.359 ;
      RECT MASK 1 19.0605 88.3735 19.1205 88.912 ;
      RECT MASK 1 19.3925 88.3735 19.4525 88.912 ;
      RECT MASK 1 19.7245 88.3735 19.7845 88.912 ;
      RECT MASK 1 20.0565 88.3735 20.1165 88.912 ;
      RECT MASK 1 20.3885 88.3735 20.4485 88.912 ;
      RECT MASK 1 20.7205 88.3735 20.7805 88.912 ;
      RECT MASK 1 14.1785 88.595 14.2385 88.912 ;
      RECT MASK 1 14.5105 88.595 14.5705 88.912 ;
      RECT MASK 1 14.8425 88.595 14.9025 88.912 ;
      RECT MASK 1 15.1745 88.595 15.2345 88.912 ;
      RECT MASK 1 15.5065 88.595 15.5665 88.912 ;
      RECT MASK 1 15.8385 88.595 15.8985 88.912 ;
      RECT MASK 1 16.1705 88.595 16.2305 88.912 ;
      RECT MASK 1 25.66 88.677 30.63 88.737 ;
      RECT MASK 1 36.326 88.947 66.476 89.007 ;
      RECT MASK 1 72.716 88.947 102.866 89.007 ;
      RECT MASK 1 7.637 89.005 7.697 93.927 ;
      RECT MASK 1 9.2135 89.05 9.2735 89.33 ;
      RECT MASK 1 11.5375 89.05 11.5975 89.33 ;
      RECT MASK 1 11.8695 89.05 11.9295 89.33 ;
      RECT MASK 1 14.2615 89.05 14.3215 89.33 ;
      RECT MASK 1 15.9215 89.05 15.9815 89.33 ;
      RECT MASK 1 16.2535 89.05 16.3135 89.33 ;
      RECT MASK 1 18.4795 89.05 18.5395 89.33 ;
      RECT MASK 1 18.8115 89.05 18.8715 89.33 ;
      RECT MASK 1 21.1355 89.05 21.1955 89.33 ;
      RECT MASK 1 9.8775 89.0915 9.9375 89.2865 ;
      RECT MASK 1 10.2095 89.0915 10.2695 89.2865 ;
      RECT MASK 1 10.5415 89.0915 10.6015 89.2865 ;
      RECT MASK 1 10.8735 89.0915 10.9335 89.2865 ;
      RECT MASK 1 11.2055 89.0915 11.2655 89.2865 ;
      RECT MASK 1 14.9255 89.0915 14.9855 89.2865 ;
      RECT MASK 1 15.2575 89.0915 15.3175 89.2865 ;
      RECT MASK 1 19.1435 89.0915 19.2035 89.2865 ;
      RECT MASK 1 19.4755 89.0915 19.5355 89.2865 ;
      RECT MASK 1 19.8075 89.0915 19.8675 89.2865 ;
      RECT MASK 1 20.1395 89.0915 20.1995 89.2865 ;
      RECT MASK 1 20.4715 89.0915 20.5315 89.2865 ;
      RECT MASK 1 6.009 89.138 6.069 92.422 ;
      RECT MASK 1 7.005 89.138 7.065 92.422 ;
      RECT MASK 1 36.326 89.199 66.476 89.259 ;
      RECT MASK 1 72.716 89.199 102.866 89.259 ;
      RECT MASK 1 18.7285 89.455 18.7885 90.24 ;
      RECT MASK 1 19.0605 89.455 19.1205 89.8075 ;
      RECT MASK 1 19.3925 89.455 19.4525 89.8075 ;
      RECT MASK 1 19.7245 89.455 19.7845 89.8075 ;
      RECT MASK 1 20.0565 89.455 20.1165 89.8075 ;
      RECT MASK 1 20.3885 89.455 20.4485 89.8075 ;
      RECT MASK 1 20.7205 89.455 20.7805 89.8075 ;
      RECT MASK 1 21.0525 89.455 21.1125 90.24 ;
      RECT MASK 1 9.1305 89.468 9.1905 90.24 ;
      RECT MASK 1 9.4625 89.468 9.5225 90.24 ;
      RECT MASK 1 9.7945 89.468 9.8545 90.24 ;
      RECT MASK 1 10.1265 89.468 10.1865 90.24 ;
      RECT MASK 1 10.4585 89.468 10.5185 90.24 ;
      RECT MASK 1 10.7905 89.468 10.8505 90.24 ;
      RECT MASK 1 11.1225 89.468 11.1825 90.24 ;
      RECT MASK 1 11.4545 89.468 11.5145 90.24 ;
      RECT MASK 1 11.7865 89.468 11.8465 90.24 ;
      RECT MASK 1 14.1785 89.468 14.2385 89.692 ;
      RECT MASK 1 14.5105 89.468 14.5705 89.692 ;
      RECT MASK 1 14.8425 89.468 14.9025 89.692 ;
      RECT MASK 1 15.1745 89.468 15.2345 89.692 ;
      RECT MASK 1 15.5065 89.468 15.5665 89.692 ;
      RECT MASK 1 15.8385 89.468 15.8985 89.692 ;
      RECT MASK 1 16.1705 89.468 16.2305 89.692 ;
      RECT MASK 1 25.66 89.577 30.63 89.637 ;
      RECT MASK 1 36.326 89.847 36.778 89.907 ;
      RECT MASK 1 37.048 89.847 65.754 89.907 ;
      RECT MASK 1 66.024 89.847 66.476 89.907 ;
      RECT MASK 1 72.716 89.847 73.168 89.907 ;
      RECT MASK 1 73.438 89.847 102.144 89.907 ;
      RECT MASK 1 102.414 89.847 102.866 89.907 ;
      RECT MASK 1 14.1585 89.905 14.2585 90.25 ;
      RECT MASK 1 14.4905 89.905 14.5905 90.25 ;
      RECT MASK 1 14.8225 89.905 14.9225 90.25 ;
      RECT MASK 1 15.1545 89.905 15.2545 90.25 ;
      RECT MASK 1 15.4865 89.905 15.5865 90.25 ;
      RECT MASK 1 15.8185 89.905 15.9185 90.25 ;
      RECT MASK 1 16.1505 89.905 16.2505 90.25 ;
      RECT MASK 1 36.326 90.099 36.778 90.159 ;
      RECT MASK 1 37.048 90.099 65.754 90.159 ;
      RECT MASK 1 66.024 90.099 66.476 90.159 ;
      RECT MASK 1 72.716 90.099 73.168 90.159 ;
      RECT MASK 1 73.438 90.099 102.144 90.159 ;
      RECT MASK 1 102.414 90.099 102.866 90.159 ;
      RECT MASK 1 25.66 90.161 25.945 90.221 ;
      RECT MASK 1 26.204 90.161 30.086 90.221 ;
      RECT MASK 1 30.345 90.161 30.63 90.221 ;
      RECT MASK 1 6.77 90.334 6.83 90.87 ;
      RECT MASK 1 8.547 90.42 8.607 90.7 ;
      RECT MASK 1 8.879 90.42 8.939 90.7 ;
      RECT MASK 1 9.211 90.42 9.271 90.7 ;
      RECT MASK 1 9.543 90.42 9.603 90.7 ;
      RECT MASK 1 9.875 90.42 9.935 90.7 ;
      RECT MASK 1 10.207 90.42 10.267 90.7 ;
      RECT MASK 1 10.539 90.42 10.599 90.7 ;
      RECT MASK 1 10.871 90.42 10.931 90.7 ;
      RECT MASK 1 11.203 90.42 11.263 90.7 ;
      RECT MASK 1 11.535 90.42 11.595 90.7 ;
      RECT MASK 1 11.867 90.42 11.927 90.7 ;
      RECT MASK 1 12.199 90.42 12.259 90.7 ;
      RECT MASK 1 13.595 90.42 13.655 90.7 ;
      RECT MASK 1 13.927 90.42 13.987 90.7 ;
      RECT MASK 1 14.259 90.42 14.319 90.7 ;
      RECT MASK 1 14.757 90.42 14.817 90.7 ;
      RECT MASK 1 15.089 90.42 15.149 90.7 ;
      RECT MASK 1 15.421 90.42 15.481 90.7 ;
      RECT MASK 1 15.753 90.42 15.813 90.7 ;
      RECT MASK 1 16.085 90.42 16.145 90.7 ;
      RECT MASK 1 16.417 90.42 16.477 90.7 ;
      RECT MASK 1 16.749 90.42 16.809 90.7 ;
      RECT MASK 1 18.145 90.42 18.205 90.7 ;
      RECT MASK 1 18.477 90.42 18.537 90.7 ;
      RECT MASK 1 18.809 90.42 18.869 90.7 ;
      RECT MASK 1 19.141 90.42 19.201 90.7 ;
      RECT MASK 1 19.473 90.42 19.533 90.7 ;
      RECT MASK 1 19.805 90.42 19.865 90.7 ;
      RECT MASK 1 20.137 90.42 20.197 90.7 ;
      RECT MASK 1 20.469 90.42 20.529 90.7 ;
      RECT MASK 1 20.801 90.42 20.861 90.7 ;
      RECT MASK 1 21.133 90.42 21.193 90.7 ;
      RECT MASK 1 21.465 90.42 21.525 90.7 ;
      RECT MASK 1 21.797 90.42 21.857 90.7 ;
      RECT MASK 1 25.66 90.423 25.944 90.483 ;
      RECT MASK 1 26.205 90.423 30.085 90.483 ;
      RECT MASK 1 30.346 90.423 30.63 90.483 ;
      RECT MASK 1 36.326 90.747 66.476 90.807 ;
      RECT MASK 1 72.716 90.747 102.866 90.807 ;
      RECT MASK 1 8.547 90.86 8.607 91.14 ;
      RECT MASK 1 8.879 90.86 8.939 91.14 ;
      RECT MASK 1 9.211 90.86 9.271 91.14 ;
      RECT MASK 1 9.543 90.86 9.603 91.14 ;
      RECT MASK 1 9.875 90.86 9.935 91.14 ;
      RECT MASK 1 10.207 90.86 10.267 91.14 ;
      RECT MASK 1 10.539 90.86 10.599 91.14 ;
      RECT MASK 1 10.871 90.86 10.931 91.14 ;
      RECT MASK 1 11.203 90.86 11.263 91.14 ;
      RECT MASK 1 11.535 90.86 11.595 91.14 ;
      RECT MASK 1 11.867 90.86 11.927 91.14 ;
      RECT MASK 1 12.199 90.86 12.259 91.14 ;
      RECT MASK 1 13.595 90.86 13.655 91.14 ;
      RECT MASK 1 13.927 90.86 13.987 91.14 ;
      RECT MASK 1 14.259 90.86 14.319 91.14 ;
      RECT MASK 1 14.757 90.86 14.817 91.14 ;
      RECT MASK 1 15.089 90.86 15.149 91.14 ;
      RECT MASK 1 15.421 90.86 15.481 91.14 ;
      RECT MASK 1 15.753 90.86 15.813 91.14 ;
      RECT MASK 1 16.085 90.86 16.145 91.14 ;
      RECT MASK 1 16.417 90.86 16.477 91.14 ;
      RECT MASK 1 16.749 90.86 16.809 91.14 ;
      RECT MASK 1 18.145 90.86 18.205 91.14 ;
      RECT MASK 1 18.477 90.86 18.537 91.14 ;
      RECT MASK 1 18.809 90.86 18.869 91.14 ;
      RECT MASK 1 19.141 90.86 19.201 91.14 ;
      RECT MASK 1 19.473 90.86 19.533 91.14 ;
      RECT MASK 1 19.805 90.86 19.865 91.14 ;
      RECT MASK 1 20.137 90.86 20.197 91.14 ;
      RECT MASK 1 20.469 90.86 20.529 91.14 ;
      RECT MASK 1 20.801 90.86 20.861 91.14 ;
      RECT MASK 1 21.133 90.86 21.193 91.14 ;
      RECT MASK 1 21.465 90.86 21.525 91.14 ;
      RECT MASK 1 21.797 90.86 21.857 91.14 ;
      RECT MASK 1 7.863 90.8615 7.963 94.359 ;
      RECT MASK 1 36.326 90.999 66.476 91.059 ;
      RECT MASK 1 72.716 90.999 102.866 91.059 ;
      RECT MASK 1 25.66 91.017 30.63 91.077 ;
      RECT MASK 1 6.424 91.205 6.484 91.499 ;
      RECT MASK 1 14.1585 91.31 14.2585 91.655 ;
      RECT MASK 1 14.4905 91.31 14.5905 91.655 ;
      RECT MASK 1 14.8225 91.31 14.9225 91.655 ;
      RECT MASK 1 15.1545 91.31 15.2545 91.655 ;
      RECT MASK 1 15.4865 91.31 15.5865 91.655 ;
      RECT MASK 1 15.8185 91.31 15.9185 91.655 ;
      RECT MASK 1 16.1505 91.31 16.2505 91.655 ;
      RECT MASK 1 8.451 91.32 8.551 93.9 ;
      RECT MASK 1 8.803 91.32 8.863 92.092 ;
      RECT MASK 1 9.135 91.32 9.195 92.092 ;
      RECT MASK 1 9.467 91.32 9.527 92.092 ;
      RECT MASK 1 9.799 91.32 9.859 92.092 ;
      RECT MASK 1 10.131 91.32 10.191 92.092 ;
      RECT MASK 1 10.463 91.32 10.523 92.092 ;
      RECT MASK 1 10.795 91.32 10.855 92.092 ;
      RECT MASK 1 11.127 91.32 11.187 92.092 ;
      RECT MASK 1 11.459 91.32 11.519 92.092 ;
      RECT MASK 1 13.8265 91.32 13.9265 93.9 ;
      RECT MASK 1 16.4825 91.32 16.5825 93.9 ;
      RECT MASK 1 18.2105 91.32 18.3105 93.9 ;
      RECT MASK 1 18.7285 91.32 18.7885 92.105 ;
      RECT MASK 1 21.0525 91.32 21.1125 92.105 ;
      RECT MASK 1 21.5305 91.32 21.6305 93.9 ;
      RECT MASK 1 6.424 91.619 6.484 93.551 ;
      RECT MASK 1 36.326 91.647 36.778 91.707 ;
      RECT MASK 1 37.048 91.647 65.754 91.707 ;
      RECT MASK 1 66.024 91.647 66.476 91.707 ;
      RECT MASK 1 72.716 91.647 73.168 91.707 ;
      RECT MASK 1 73.438 91.647 102.144 91.707 ;
      RECT MASK 1 102.414 91.647 102.866 91.707 ;
      RECT MASK 1 19.0605 91.7525 19.1205 92.105 ;
      RECT MASK 1 19.3925 91.7525 19.4525 92.105 ;
      RECT MASK 1 19.7245 91.7525 19.7845 92.105 ;
      RECT MASK 1 20.0565 91.7525 20.1165 92.105 ;
      RECT MASK 1 20.3885 91.7525 20.4485 92.105 ;
      RECT MASK 1 20.7205 91.7525 20.7805 92.105 ;
      RECT MASK 1 14.1785 91.868 14.2385 92.092 ;
      RECT MASK 1 14.5105 91.868 14.5705 92.092 ;
      RECT MASK 1 14.8425 91.868 14.9025 92.095 ;
      RECT MASK 1 15.1745 91.868 15.2345 92.095 ;
      RECT MASK 1 15.5065 91.868 15.5665 92.095 ;
      RECT MASK 1 15.8385 91.868 15.8985 92.092 ;
      RECT MASK 1 16.1705 91.868 16.2305 92.092 ;
      RECT MASK 1 36.326 91.899 36.778 91.959 ;
      RECT MASK 1 37.048 91.899 65.754 91.959 ;
      RECT MASK 1 66.024 91.899 66.476 91.959 ;
      RECT MASK 1 72.716 91.899 73.168 91.959 ;
      RECT MASK 1 73.438 91.899 102.144 91.959 ;
      RECT MASK 1 102.414 91.899 102.866 91.959 ;
      RECT MASK 1 25.237 92.149 31.053 92.289 ;
      RECT MASK 1 8.886 92.23 8.946 92.51 ;
      RECT MASK 1 11.21 92.23 11.27 92.51 ;
      RECT MASK 1 11.542 92.23 11.602 92.51 ;
      RECT MASK 1 14.2615 92.23 14.3215 92.51 ;
      RECT MASK 1 15.9215 92.23 15.9815 92.51 ;
      RECT MASK 1 16.2535 92.23 16.3135 92.51 ;
      RECT MASK 1 18.4795 92.23 18.5395 92.51 ;
      RECT MASK 1 18.8115 92.23 18.8715 92.51 ;
      RECT MASK 1 21.1355 92.23 21.1955 92.51 ;
      RECT MASK 1 9.882 92.2735 9.942 92.4685 ;
      RECT MASK 1 10.214 92.2735 10.274 92.4685 ;
      RECT MASK 1 10.546 92.2735 10.606 92.4685 ;
      RECT MASK 1 10.878 92.2735 10.938 92.4685 ;
      RECT MASK 1 14.9255 92.2735 14.9855 92.4685 ;
      RECT MASK 1 15.2575 92.2735 15.3175 92.4685 ;
      RECT MASK 1 19.1435 92.2735 19.2035 92.4685 ;
      RECT MASK 1 19.4755 92.2735 19.5355 92.4685 ;
      RECT MASK 1 19.8075 92.2735 19.8675 92.4685 ;
      RECT MASK 1 20.1395 92.2735 20.1995 92.4685 ;
      RECT MASK 1 20.4715 92.2735 20.5315 92.4685 ;
      RECT MASK 1 36.326 92.547 66.476 92.607 ;
      RECT MASK 1 72.716 92.547 102.866 92.607 ;
      RECT MASK 1 6.009 92.618 6.069 94.345 ;
      RECT MASK 1 7.005 92.618 7.065 94.345 ;
      RECT MASK 1 8.803 92.648 8.863 93.9 ;
      RECT MASK 1 9.135 92.648 9.195 93.9 ;
      RECT MASK 1 9.467 92.648 9.527 93.9 ;
      RECT MASK 1 9.799 92.648 9.859 93.9 ;
      RECT MASK 1 10.131 92.648 10.191 93.9 ;
      RECT MASK 1 10.463 92.648 10.523 93.9 ;
      RECT MASK 1 10.795 92.648 10.855 93.9 ;
      RECT MASK 1 11.127 92.648 11.187 93.9 ;
      RECT MASK 1 11.459 92.648 11.519 93.9 ;
      RECT MASK 1 14.1785 92.648 14.2385 92.965 ;
      RECT MASK 1 14.5105 92.648 14.5705 92.965 ;
      RECT MASK 1 14.8425 92.648 14.9025 92.965 ;
      RECT MASK 1 15.1745 92.648 15.2345 92.965 ;
      RECT MASK 1 15.5065 92.648 15.5665 92.965 ;
      RECT MASK 1 15.8385 92.648 15.8985 92.965 ;
      RECT MASK 1 16.1705 92.648 16.2305 92.965 ;
      RECT MASK 1 18.7285 92.648 18.7885 93.9 ;
      RECT MASK 1 19.0605 92.648 19.1205 93.1865 ;
      RECT MASK 1 19.3925 92.648 19.4525 93.1865 ;
      RECT MASK 1 19.7245 92.648 19.7845 93.1865 ;
      RECT MASK 1 20.0565 92.648 20.1165 93.1865 ;
      RECT MASK 1 20.3885 92.648 20.4485 93.1865 ;
      RECT MASK 1 20.7205 92.648 20.7805 93.1865 ;
      RECT MASK 1 21.0525 92.648 21.1125 93.9 ;
      RECT MASK 1 36.326 92.799 66.476 92.859 ;
      RECT MASK 1 72.716 92.799 102.866 92.859 ;
      RECT MASK 1 14.1585 93.17 14.2585 93.9 ;
      RECT MASK 1 14.4905 93.17 14.5905 93.9 ;
      RECT MASK 1 14.8225 93.17 14.9225 93.9 ;
      RECT MASK 1 15.1545 93.17 15.2545 93.9 ;
      RECT MASK 1 15.4865 93.17 15.5865 93.9 ;
      RECT MASK 1 15.8185 93.17 15.9185 93.9 ;
      RECT MASK 1 16.1505 93.17 16.2505 93.9 ;
      RECT MASK 1 36.326 93.447 36.778 93.507 ;
      RECT MASK 1 37.048 93.447 65.754 93.507 ;
      RECT MASK 1 66.024 93.447 66.476 93.507 ;
      RECT MASK 1 72.716 93.447 73.168 93.507 ;
      RECT MASK 1 73.438 93.447 102.144 93.507 ;
      RECT MASK 1 102.414 93.447 102.866 93.507 ;
      RECT MASK 1 6.59 93.571 6.65 93.84 ;
      RECT MASK 1 36.326 93.699 36.778 93.759 ;
      RECT MASK 1 37.048 93.699 65.754 93.759 ;
      RECT MASK 1 66.024 93.699 66.476 93.759 ;
      RECT MASK 1 72.716 93.699 73.168 93.759 ;
      RECT MASK 1 73.438 93.699 102.144 93.759 ;
      RECT MASK 1 102.414 93.699 102.866 93.759 ;
      RECT MASK 1 25.237 93.871 31.053 94.011 ;
      RECT MASK 1 8.547 94.07 8.607 94.35 ;
      RECT MASK 1 8.879 94.07 8.939 94.35 ;
      RECT MASK 1 9.211 94.07 9.271 94.35 ;
      RECT MASK 1 9.543 94.07 9.603 94.35 ;
      RECT MASK 1 9.875 94.07 9.935 94.35 ;
      RECT MASK 1 10.207 94.07 10.267 94.35 ;
      RECT MASK 1 10.539 94.07 10.599 94.35 ;
      RECT MASK 1 10.871 94.07 10.931 94.35 ;
      RECT MASK 1 11.203 94.07 11.263 94.35 ;
      RECT MASK 1 11.535 94.07 11.595 94.35 ;
      RECT MASK 1 11.867 94.07 11.927 94.35 ;
      RECT MASK 1 12.199 94.07 12.259 94.35 ;
      RECT MASK 1 13.595 94.07 13.655 94.35 ;
      RECT MASK 1 13.927 94.07 13.987 94.35 ;
      RECT MASK 1 14.259 94.07 14.319 94.35 ;
      RECT MASK 1 14.757 94.07 14.817 94.35 ;
      RECT MASK 1 15.089 94.07 15.149 94.35 ;
      RECT MASK 1 15.421 94.07 15.481 94.35 ;
      RECT MASK 1 15.753 94.07 15.813 94.35 ;
      RECT MASK 1 16.085 94.07 16.145 94.35 ;
      RECT MASK 1 16.417 94.07 16.477 94.35 ;
      RECT MASK 1 16.749 94.07 16.809 94.35 ;
      RECT MASK 1 18.145 94.07 18.205 94.35 ;
      RECT MASK 1 18.477 94.07 18.537 94.35 ;
      RECT MASK 1 18.809 94.07 18.869 94.35 ;
      RECT MASK 1 19.141 94.07 19.201 94.35 ;
      RECT MASK 1 19.473 94.07 19.533 94.35 ;
      RECT MASK 1 19.805 94.07 19.865 94.35 ;
      RECT MASK 1 20.137 94.07 20.197 94.35 ;
      RECT MASK 1 20.469 94.07 20.529 94.35 ;
      RECT MASK 1 20.801 94.07 20.861 94.35 ;
      RECT MASK 1 21.133 94.07 21.193 94.35 ;
      RECT MASK 1 21.465 94.07 21.525 94.35 ;
      RECT MASK 1 21.797 94.07 21.857 94.35 ;
      RECT MASK 1 36.326 94.347 66.476 94.407 ;
      RECT MASK 1 72.716 94.347 102.866 94.407 ;
      RECT MASK 1 36.326 94.599 66.476 94.659 ;
      RECT MASK 1 72.716 94.599 102.866 94.659 ;
      RECT MASK 1 34.008 94.625 34.068 95.335 ;
      RECT MASK 1 34.257 94.625 34.317 95.335 ;
      RECT MASK 1 34.506 94.625 34.566 95.335 ;
      RECT MASK 1 34.755 94.625 34.815 95.335 ;
      RECT MASK 1 35.004 94.625 35.064 95.335 ;
      RECT MASK 1 35.253 94.625 35.313 95.335 ;
      RECT MASK 1 67.572 94.625 67.632 95.335 ;
      RECT MASK 1 67.821 94.625 67.881 95.335 ;
      RECT MASK 1 68.07 94.625 68.13 95.335 ;
      RECT MASK 1 68.319 94.625 68.379 95.335 ;
      RECT MASK 1 68.568 94.625 68.628 95.335 ;
      RECT MASK 1 70.398 94.715 70.458 95.425 ;
      RECT MASK 1 70.647 94.715 70.707 95.425 ;
      RECT MASK 1 70.896 94.715 70.956 95.425 ;
      RECT MASK 1 71.145 94.715 71.205 95.425 ;
      RECT MASK 1 71.394 94.715 71.454 95.425 ;
      RECT MASK 1 71.643 94.715 71.703 95.425 ;
      RECT MASK 1 103.879 94.715 103.939 95.425 ;
      RECT MASK 1 104.128 94.715 104.188 95.425 ;
      RECT MASK 1 104.377 94.715 104.437 95.425 ;
      RECT MASK 1 104.626 94.715 104.686 95.425 ;
      RECT MASK 1 104.875 94.715 104.935 95.425 ;
      RECT MASK 1 105.124 94.715 105.184 95.425 ;
      RECT MASK 1 33.51 95.075 33.57 95.335 ;
      RECT MASK 1 33.759 95.075 33.819 95.335 ;
      RECT MASK 1 68.817 95.075 68.877 95.335 ;
      RECT MASK 1 69.066 95.075 69.126 95.335 ;
      RECT MASK 1 36.1535 95.111 66.6485 95.211 ;
      RECT MASK 1 72.5435 95.111 103.0385 95.211 ;
      RECT MASK 1 69.9 95.165 69.96 95.425 ;
      RECT MASK 1 70.149 95.165 70.209 95.425 ;
      RECT MASK 1 105.373 95.165 105.433 95.425 ;
      RECT MASK 1 105.622 95.165 105.682 95.425 ;
      RECT MASK 1 1.454 97.25 1.554 107.66 ;
      RECT MASK 1 44.282 97.25 44.382 107.66 ;
      RECT MASK 1 44.846 97.25 44.946 107.66 ;
      RECT MASK 1 87.674 97.25 87.774 107.67 ;
      RECT MASK 1 88.238 97.25 88.338 107.67 ;
      RECT MASK 1 2.201 97.6 2.261 107.66 ;
      RECT MASK 1 2.475 97.6 2.535 107.61 ;
      RECT MASK 1 2.749 97.6 2.809 107.61 ;
      RECT MASK 1 3.023 97.6 3.083 107.61 ;
      RECT MASK 1 3.297 97.6 3.357 107.61 ;
      RECT MASK 1 3.571 97.6 3.631 107.61 ;
      RECT MASK 1 3.845 97.6 3.905 107.61 ;
      RECT MASK 1 4.119 97.6 4.179 107.61 ;
      RECT MASK 1 4.393 97.6 4.453 107.61 ;
      RECT MASK 1 4.667 97.6 4.727 107.61 ;
      RECT MASK 1 4.941 97.6 5.001 107.61 ;
      RECT MASK 1 5.215 97.6 5.275 107.61 ;
      RECT MASK 1 5.489 97.6 5.549 107.61 ;
      RECT MASK 1 5.763 97.6 5.823 107.61 ;
      RECT MASK 1 6.037 97.6 6.097 107.61 ;
      RECT MASK 1 6.311 97.6 6.371 107.61 ;
      RECT MASK 1 6.585 97.6 6.645 107.61 ;
      RECT MASK 1 6.859 97.6 6.919 107.61 ;
      RECT MASK 1 7.133 97.6 7.193 107.61 ;
      RECT MASK 1 7.407 97.6 7.467 107.61 ;
      RECT MASK 1 7.681 97.6 7.741 107.61 ;
      RECT MASK 1 7.955 97.6 8.015 107.61 ;
      RECT MASK 1 8.229 97.6 8.289 107.61 ;
      RECT MASK 1 8.503 97.6 8.563 107.61 ;
      RECT MASK 1 8.777 97.6 8.837 107.61 ;
      RECT MASK 1 9.051 97.6 9.111 107.61 ;
      RECT MASK 1 9.325 97.6 9.385 107.61 ;
      RECT MASK 1 9.599 97.6 9.659 107.61 ;
      RECT MASK 1 9.873 97.6 9.933 107.61 ;
      RECT MASK 1 10.147 97.6 10.207 107.61 ;
      RECT MASK 1 10.421 97.6 10.481 107.61 ;
      RECT MASK 1 10.695 97.6 10.755 107.61 ;
      RECT MASK 1 10.969 97.6 11.029 107.61 ;
      RECT MASK 1 11.243 97.6 11.303 107.61 ;
      RECT MASK 1 11.517 97.6 11.577 107.61 ;
      RECT MASK 1 11.791 97.6 11.851 107.61 ;
      RECT MASK 1 12.065 97.6 12.125 107.61 ;
      RECT MASK 1 12.339 97.6 12.399 107.61 ;
      RECT MASK 1 12.613 97.6 12.673 107.61 ;
      RECT MASK 1 12.887 97.6 12.947 107.61 ;
      RECT MASK 1 13.161 97.6 13.221 107.61 ;
      RECT MASK 1 13.435 97.6 13.495 107.61 ;
      RECT MASK 1 13.709 97.6 13.769 107.61 ;
      RECT MASK 1 13.983 97.6 14.043 107.61 ;
      RECT MASK 1 14.257 97.6 14.317 107.61 ;
      RECT MASK 1 14.531 97.6 14.591 107.61 ;
      RECT MASK 1 14.805 97.6 14.865 107.61 ;
      RECT MASK 1 15.079 97.6 15.139 107.61 ;
      RECT MASK 1 15.353 97.6 15.413 107.61 ;
      RECT MASK 1 15.627 97.6 15.687 107.61 ;
      RECT MASK 1 15.901 97.6 15.961 107.61 ;
      RECT MASK 1 16.175 97.6 16.235 107.61 ;
      RECT MASK 1 16.449 97.6 16.509 107.61 ;
      RECT MASK 1 16.723 97.6 16.783 107.61 ;
      RECT MASK 1 16.997 97.6 17.057 107.61 ;
      RECT MASK 1 17.271 97.6 17.331 107.61 ;
      RECT MASK 1 17.545 97.6 17.605 107.61 ;
      RECT MASK 1 17.819 97.6 17.879 107.61 ;
      RECT MASK 1 18.093 97.6 18.153 107.61 ;
      RECT MASK 1 18.367 97.6 18.427 107.61 ;
      RECT MASK 1 18.641 97.6 18.701 107.61 ;
      RECT MASK 1 18.915 97.6 18.975 107.61 ;
      RECT MASK 1 19.189 97.6 19.249 107.61 ;
      RECT MASK 1 19.463 97.6 19.523 107.61 ;
      RECT MASK 1 19.737 97.6 19.797 107.61 ;
      RECT MASK 1 20.011 97.6 20.071 107.61 ;
      RECT MASK 1 20.285 97.6 20.345 107.61 ;
      RECT MASK 1 20.559 97.6 20.619 107.61 ;
      RECT MASK 1 20.833 97.6 20.893 107.61 ;
      RECT MASK 1 21.107 97.6 21.167 107.61 ;
      RECT MASK 1 21.381 97.6 21.441 107.61 ;
      RECT MASK 1 21.655 97.6 21.715 107.61 ;
      RECT MASK 1 21.929 97.6 21.989 107.61 ;
      RECT MASK 1 22.203 97.6 22.263 107.61 ;
      RECT MASK 1 22.477 97.6 22.537 107.61 ;
      RECT MASK 1 22.751 97.6 22.811 107.61 ;
      RECT MASK 1 23.025 97.6 23.085 107.61 ;
      RECT MASK 1 23.299 97.6 23.359 107.61 ;
      RECT MASK 1 23.573 97.6 23.633 107.61 ;
      RECT MASK 1 23.847 97.6 23.907 107.61 ;
      RECT MASK 1 24.121 97.6 24.181 107.61 ;
      RECT MASK 1 24.395 97.6 24.455 107.61 ;
      RECT MASK 1 24.669 97.6 24.729 107.61 ;
      RECT MASK 1 24.943 97.6 25.003 107.61 ;
      RECT MASK 1 25.217 97.6 25.277 107.61 ;
      RECT MASK 1 25.491 97.6 25.551 107.61 ;
      RECT MASK 1 25.765 97.6 25.825 107.61 ;
      RECT MASK 1 26.039 97.6 26.099 107.61 ;
      RECT MASK 1 26.313 97.6 26.373 107.61 ;
      RECT MASK 1 26.587 97.6 26.647 107.61 ;
      RECT MASK 1 26.861 97.6 26.921 107.61 ;
      RECT MASK 1 27.135 97.6 27.195 107.61 ;
      RECT MASK 1 27.409 97.6 27.469 107.61 ;
      RECT MASK 1 27.683 97.6 27.743 107.61 ;
      RECT MASK 1 27.957 97.6 28.017 107.61 ;
      RECT MASK 1 28.231 97.6 28.291 107.61 ;
      RECT MASK 1 28.505 97.6 28.565 107.61 ;
      RECT MASK 1 28.779 97.6 28.839 107.61 ;
      RECT MASK 1 29.053 97.6 29.113 107.61 ;
      RECT MASK 1 29.327 97.6 29.387 107.61 ;
      RECT MASK 1 29.601 97.6 29.661 107.61 ;
      RECT MASK 1 29.875 97.6 29.935 107.61 ;
      RECT MASK 1 30.149 97.6 30.209 107.61 ;
      RECT MASK 1 30.423 97.6 30.483 107.61 ;
      RECT MASK 1 30.697 97.6 30.757 107.61 ;
      RECT MASK 1 30.971 97.6 31.031 107.61 ;
      RECT MASK 1 31.245 97.6 31.305 107.61 ;
      RECT MASK 1 31.519 97.6 31.579 107.61 ;
      RECT MASK 1 31.793 97.6 31.853 107.61 ;
      RECT MASK 1 32.067 97.6 32.127 107.61 ;
      RECT MASK 1 32.341 97.6 32.401 107.61 ;
      RECT MASK 1 32.615 97.6 32.675 107.61 ;
      RECT MASK 1 32.889 97.6 32.949 107.61 ;
      RECT MASK 1 33.163 97.6 33.223 107.61 ;
      RECT MASK 1 33.437 97.6 33.497 107.61 ;
      RECT MASK 1 33.711 97.6 33.771 107.61 ;
      RECT MASK 1 33.985 97.6 34.045 107.61 ;
      RECT MASK 1 34.259 97.6 34.319 107.61 ;
      RECT MASK 1 34.533 97.6 34.593 107.61 ;
      RECT MASK 1 34.807 97.6 34.867 107.61 ;
      RECT MASK 1 35.081 97.6 35.141 107.61 ;
      RECT MASK 1 35.355 97.6 35.415 107.61 ;
      RECT MASK 1 35.629 97.6 35.689 107.61 ;
      RECT MASK 1 35.903 97.6 35.963 107.61 ;
      RECT MASK 1 36.177 97.6 36.237 107.61 ;
      RECT MASK 1 36.451 97.6 36.511 107.61 ;
      RECT MASK 1 36.725 97.6 36.785 107.61 ;
      RECT MASK 1 36.999 97.6 37.059 107.61 ;
      RECT MASK 1 37.273 97.6 37.333 107.61 ;
      RECT MASK 1 37.547 97.6 37.607 107.61 ;
      RECT MASK 1 37.821 97.6 37.881 107.61 ;
      RECT MASK 1 38.095 97.6 38.155 107.61 ;
      RECT MASK 1 38.369 97.6 38.429 107.61 ;
      RECT MASK 1 38.643 97.6 38.703 107.61 ;
      RECT MASK 1 38.917 97.6 38.977 107.61 ;
      RECT MASK 1 39.191 97.6 39.251 107.61 ;
      RECT MASK 1 39.465 97.6 39.525 107.61 ;
      RECT MASK 1 39.739 97.6 39.799 107.61 ;
      RECT MASK 1 40.013 97.6 40.073 107.61 ;
      RECT MASK 1 40.287 97.6 40.347 107.61 ;
      RECT MASK 1 40.561 97.6 40.621 107.61 ;
      RECT MASK 1 40.835 97.6 40.895 107.61 ;
      RECT MASK 1 41.109 97.6 41.169 107.61 ;
      RECT MASK 1 41.383 97.6 41.443 107.61 ;
      RECT MASK 1 41.657 97.6 41.717 107.61 ;
      RECT MASK 1 41.931 97.6 41.991 107.61 ;
      RECT MASK 1 42.205 97.6 42.265 107.61 ;
      RECT MASK 1 42.479 97.6 42.539 107.61 ;
      RECT MASK 1 42.753 97.6 42.813 107.61 ;
      RECT MASK 1 43.027 97.6 43.087 107.61 ;
      RECT MASK 1 43.301 97.6 43.361 107.61 ;
      RECT MASK 1 43.575 97.6 43.635 107.66 ;
      RECT MASK 1 45.593 97.6 45.653 107.66 ;
      RECT MASK 1 45.867 97.6 45.927 107.61 ;
      RECT MASK 1 46.141 97.6 46.201 107.61 ;
      RECT MASK 1 46.415 97.6 46.475 107.61 ;
      RECT MASK 1 46.689 97.6 46.749 107.61 ;
      RECT MASK 1 46.963 97.6 47.023 107.61 ;
      RECT MASK 1 47.237 97.6 47.297 107.61 ;
      RECT MASK 1 47.511 97.6 47.571 107.61 ;
      RECT MASK 1 47.785 97.6 47.845 107.61 ;
      RECT MASK 1 48.059 97.6 48.119 107.61 ;
      RECT MASK 1 48.333 97.6 48.393 107.61 ;
      RECT MASK 1 48.607 97.6 48.667 107.61 ;
      RECT MASK 1 48.881 97.6 48.941 107.61 ;
      RECT MASK 1 49.155 97.6 49.215 107.61 ;
      RECT MASK 1 49.429 97.6 49.489 107.61 ;
      RECT MASK 1 49.703 97.6 49.763 107.61 ;
      RECT MASK 1 49.977 97.6 50.037 107.61 ;
      RECT MASK 1 50.251 97.6 50.311 107.61 ;
      RECT MASK 1 50.525 97.6 50.585 107.61 ;
      RECT MASK 1 50.799 97.6 50.859 107.61 ;
      RECT MASK 1 51.073 97.6 51.133 107.61 ;
      RECT MASK 1 51.347 97.6 51.407 107.61 ;
      RECT MASK 1 51.621 97.6 51.681 107.61 ;
      RECT MASK 1 51.895 97.6 51.955 107.61 ;
      RECT MASK 1 52.169 97.6 52.229 107.61 ;
      RECT MASK 1 52.443 97.6 52.503 107.61 ;
      RECT MASK 1 52.717 97.6 52.777 107.61 ;
      RECT MASK 1 52.991 97.6 53.051 107.61 ;
      RECT MASK 1 53.265 97.6 53.325 107.61 ;
      RECT MASK 1 53.539 97.6 53.599 107.61 ;
      RECT MASK 1 53.813 97.6 53.873 107.61 ;
      RECT MASK 1 54.087 97.6 54.147 107.61 ;
      RECT MASK 1 54.361 97.6 54.421 107.61 ;
      RECT MASK 1 54.635 97.6 54.695 107.61 ;
      RECT MASK 1 54.909 97.6 54.969 107.61 ;
      RECT MASK 1 55.183 97.6 55.243 107.61 ;
      RECT MASK 1 55.457 97.6 55.517 107.61 ;
      RECT MASK 1 55.731 97.6 55.791 107.61 ;
      RECT MASK 1 56.005 97.6 56.065 107.61 ;
      RECT MASK 1 56.279 97.6 56.339 107.61 ;
      RECT MASK 1 56.553 97.6 56.613 107.61 ;
      RECT MASK 1 56.827 97.6 56.887 107.61 ;
      RECT MASK 1 57.101 97.6 57.161 107.61 ;
      RECT MASK 1 57.375 97.6 57.435 107.61 ;
      RECT MASK 1 57.649 97.6 57.709 107.61 ;
      RECT MASK 1 57.923 97.6 57.983 107.61 ;
      RECT MASK 1 58.197 97.6 58.257 107.61 ;
      RECT MASK 1 58.471 97.6 58.531 107.61 ;
      RECT MASK 1 58.745 97.6 58.805 107.61 ;
      RECT MASK 1 59.019 97.6 59.079 107.61 ;
      RECT MASK 1 59.293 97.6 59.353 107.61 ;
      RECT MASK 1 59.567 97.6 59.627 107.61 ;
      RECT MASK 1 59.841 97.6 59.901 107.61 ;
      RECT MASK 1 60.115 97.6 60.175 107.61 ;
      RECT MASK 1 60.389 97.6 60.449 107.61 ;
      RECT MASK 1 60.663 97.6 60.723 107.61 ;
      RECT MASK 1 60.937 97.6 60.997 107.61 ;
      RECT MASK 1 61.211 97.6 61.271 107.61 ;
      RECT MASK 1 61.485 97.6 61.545 107.61 ;
      RECT MASK 1 61.759 97.6 61.819 107.61 ;
      RECT MASK 1 62.033 97.6 62.093 107.61 ;
      RECT MASK 1 62.307 97.6 62.367 107.61 ;
      RECT MASK 1 62.581 97.6 62.641 107.61 ;
      RECT MASK 1 62.855 97.6 62.915 107.61 ;
      RECT MASK 1 63.129 97.6 63.189 107.61 ;
      RECT MASK 1 63.403 97.6 63.463 107.61 ;
      RECT MASK 1 63.677 97.6 63.737 107.61 ;
      RECT MASK 1 63.951 97.6 64.011 107.61 ;
      RECT MASK 1 64.225 97.6 64.285 107.61 ;
      RECT MASK 1 64.499 97.6 64.559 107.61 ;
      RECT MASK 1 64.773 97.6 64.833 107.61 ;
      RECT MASK 1 65.047 97.6 65.107 107.61 ;
      RECT MASK 1 65.321 97.6 65.381 107.61 ;
      RECT MASK 1 65.595 97.6 65.655 107.61 ;
      RECT MASK 1 65.869 97.6 65.929 107.61 ;
      RECT MASK 1 66.143 97.6 66.203 107.61 ;
      RECT MASK 1 66.417 97.6 66.477 107.61 ;
      RECT MASK 1 66.691 97.6 66.751 107.61 ;
      RECT MASK 1 66.965 97.6 67.025 107.61 ;
      RECT MASK 1 67.239 97.6 67.299 107.61 ;
      RECT MASK 1 67.513 97.6 67.573 107.61 ;
      RECT MASK 1 67.787 97.6 67.847 107.61 ;
      RECT MASK 1 68.061 97.6 68.121 107.61 ;
      RECT MASK 1 68.335 97.6 68.395 107.61 ;
      RECT MASK 1 68.609 97.6 68.669 107.61 ;
      RECT MASK 1 68.883 97.6 68.943 107.61 ;
      RECT MASK 1 69.157 97.6 69.217 107.61 ;
      RECT MASK 1 69.431 97.6 69.491 107.61 ;
      RECT MASK 1 69.705 97.6 69.765 107.61 ;
      RECT MASK 1 69.979 97.6 70.039 107.61 ;
      RECT MASK 1 70.253 97.6 70.313 107.61 ;
      RECT MASK 1 70.527 97.6 70.587 107.61 ;
      RECT MASK 1 70.801 97.6 70.861 107.61 ;
      RECT MASK 1 71.075 97.6 71.135 107.61 ;
      RECT MASK 1 71.349 97.6 71.409 107.61 ;
      RECT MASK 1 71.623 97.6 71.683 107.61 ;
      RECT MASK 1 71.897 97.6 71.957 107.61 ;
      RECT MASK 1 72.171 97.6 72.231 107.61 ;
      RECT MASK 1 72.445 97.6 72.505 107.61 ;
      RECT MASK 1 72.719 97.6 72.779 107.61 ;
      RECT MASK 1 72.993 97.6 73.053 107.61 ;
      RECT MASK 1 73.267 97.6 73.327 107.61 ;
      RECT MASK 1 73.541 97.6 73.601 107.61 ;
      RECT MASK 1 73.815 97.6 73.875 107.61 ;
      RECT MASK 1 74.089 97.6 74.149 107.61 ;
      RECT MASK 1 74.363 97.6 74.423 107.61 ;
      RECT MASK 1 74.637 97.6 74.697 107.61 ;
      RECT MASK 1 74.911 97.6 74.971 107.61 ;
      RECT MASK 1 75.185 97.6 75.245 107.61 ;
      RECT MASK 1 75.459 97.6 75.519 107.61 ;
      RECT MASK 1 75.733 97.6 75.793 107.61 ;
      RECT MASK 1 76.007 97.6 76.067 107.61 ;
      RECT MASK 1 76.281 97.6 76.341 107.61 ;
      RECT MASK 1 76.555 97.6 76.615 107.61 ;
      RECT MASK 1 76.829 97.6 76.889 107.61 ;
      RECT MASK 1 77.103 97.6 77.163 107.61 ;
      RECT MASK 1 77.377 97.6 77.437 107.61 ;
      RECT MASK 1 77.651 97.6 77.711 107.61 ;
      RECT MASK 1 77.925 97.6 77.985 107.61 ;
      RECT MASK 1 78.199 97.6 78.259 107.61 ;
      RECT MASK 1 78.473 97.6 78.533 107.61 ;
      RECT MASK 1 78.747 97.6 78.807 107.61 ;
      RECT MASK 1 79.021 97.6 79.081 107.61 ;
      RECT MASK 1 79.295 97.6 79.355 107.61 ;
      RECT MASK 1 79.569 97.6 79.629 107.61 ;
      RECT MASK 1 79.843 97.6 79.903 107.61 ;
      RECT MASK 1 80.117 97.6 80.177 107.61 ;
      RECT MASK 1 80.391 97.6 80.451 107.61 ;
      RECT MASK 1 80.665 97.6 80.725 107.61 ;
      RECT MASK 1 80.939 97.6 80.999 107.61 ;
      RECT MASK 1 81.213 97.6 81.273 107.61 ;
      RECT MASK 1 81.487 97.6 81.547 107.61 ;
      RECT MASK 1 81.761 97.6 81.821 107.61 ;
      RECT MASK 1 82.035 97.6 82.095 107.61 ;
      RECT MASK 1 82.309 97.6 82.369 107.61 ;
      RECT MASK 1 82.583 97.6 82.643 107.61 ;
      RECT MASK 1 82.857 97.6 82.917 107.61 ;
      RECT MASK 1 83.131 97.6 83.191 107.61 ;
      RECT MASK 1 83.405 97.6 83.465 107.61 ;
      RECT MASK 1 83.679 97.6 83.739 107.61 ;
      RECT MASK 1 83.953 97.6 84.013 107.61 ;
      RECT MASK 1 84.227 97.6 84.287 107.61 ;
      RECT MASK 1 84.501 97.6 84.561 107.61 ;
      RECT MASK 1 84.775 97.6 84.835 107.61 ;
      RECT MASK 1 85.049 97.6 85.109 107.61 ;
      RECT MASK 1 85.323 97.6 85.383 107.61 ;
      RECT MASK 1 85.597 97.6 85.657 107.61 ;
      RECT MASK 1 85.871 97.6 85.931 107.61 ;
      RECT MASK 1 86.145 97.6 86.205 107.61 ;
      RECT MASK 1 86.419 97.6 86.479 107.61 ;
      RECT MASK 1 86.693 97.6 86.753 107.61 ;
      RECT MASK 1 86.967 97.6 87.027 107.66 ;
      RECT MASK 1 88.952 97.6 89.012 107.66 ;
      RECT MASK 1 89.226 97.6 89.286 107.61 ;
      RECT MASK 1 89.5 97.6 89.56 107.61 ;
      RECT MASK 1 89.774 97.6 89.834 107.61 ;
      RECT MASK 1 90.048 97.6 90.108 107.61 ;
      RECT MASK 1 90.322 97.6 90.382 107.61 ;
      RECT MASK 1 90.596 97.6 90.656 107.61 ;
      RECT MASK 1 90.87 97.6 90.93 107.61 ;
      RECT MASK 1 91.144 97.6 91.204 107.61 ;
      RECT MASK 1 91.418 97.6 91.478 107.61 ;
      RECT MASK 1 91.692 97.6 91.752 107.61 ;
      RECT MASK 1 91.966 97.6 92.026 107.61 ;
      RECT MASK 1 92.24 97.6 92.3 107.61 ;
      RECT MASK 1 92.514 97.6 92.574 107.61 ;
      RECT MASK 1 92.788 97.6 92.848 107.61 ;
      RECT MASK 1 93.062 97.6 93.122 107.61 ;
      RECT MASK 1 93.336 97.6 93.396 107.61 ;
      RECT MASK 1 93.61 97.6 93.67 107.61 ;
      RECT MASK 1 93.884 97.6 93.944 107.61 ;
      RECT MASK 1 94.158 97.6 94.218 107.61 ;
      RECT MASK 1 94.432 97.6 94.492 107.61 ;
      RECT MASK 1 94.706 97.6 94.766 107.61 ;
      RECT MASK 1 94.98 97.6 95.04 107.61 ;
      RECT MASK 1 95.254 97.6 95.314 107.61 ;
      RECT MASK 1 95.528 97.6 95.588 107.61 ;
      RECT MASK 1 95.802 97.6 95.862 107.61 ;
      RECT MASK 1 96.076 97.6 96.136 107.61 ;
      RECT MASK 1 96.35 97.6 96.41 107.61 ;
      RECT MASK 1 96.624 97.6 96.684 107.61 ;
      RECT MASK 1 96.898 97.6 96.958 107.61 ;
      RECT MASK 1 97.172 97.6 97.232 107.61 ;
      RECT MASK 1 97.446 97.6 97.506 107.61 ;
      RECT MASK 1 97.72 97.6 97.78 107.61 ;
      RECT MASK 1 97.994 97.6 98.054 107.61 ;
      RECT MASK 1 98.268 97.6 98.328 107.61 ;
      RECT MASK 1 98.542 97.6 98.602 107.61 ;
      RECT MASK 1 98.816 97.6 98.876 107.61 ;
      RECT MASK 1 99.09 97.6 99.15 107.61 ;
      RECT MASK 1 99.364 97.6 99.424 107.61 ;
      RECT MASK 1 99.638 97.6 99.698 107.61 ;
      RECT MASK 1 99.912 97.6 99.972 107.61 ;
      RECT MASK 1 100.186 97.6 100.246 107.61 ;
      RECT MASK 1 100.46 97.6 100.52 107.61 ;
      RECT MASK 1 100.734 97.6 100.794 107.61 ;
      RECT MASK 1 101.008 97.6 101.068 107.61 ;
      RECT MASK 1 101.282 97.6 101.342 107.61 ;
      RECT MASK 1 101.556 97.6 101.616 107.61 ;
      RECT MASK 1 101.83 97.6 101.89 107.61 ;
      RECT MASK 1 102.104 97.6 102.164 107.61 ;
      RECT MASK 1 102.378 97.6 102.438 107.61 ;
      RECT MASK 1 102.652 97.6 102.712 107.61 ;
      RECT MASK 1 102.926 97.6 102.986 107.61 ;
      RECT MASK 1 103.2 97.6 103.26 107.61 ;
      RECT MASK 1 103.474 97.6 103.534 107.61 ;
      RECT MASK 1 103.748 97.6 103.808 107.61 ;
      RECT MASK 1 104.022 97.6 104.082 107.61 ;
      RECT MASK 1 104.296 97.6 104.356 107.61 ;
      RECT MASK 1 104.57 97.6 104.63 107.61 ;
      RECT MASK 1 104.844 97.6 104.904 107.61 ;
      RECT MASK 1 105.118 97.6 105.178 107.61 ;
      RECT MASK 1 105.392 97.6 105.452 107.61 ;
      RECT MASK 1 105.666 97.6 105.726 107.61 ;
      RECT MASK 1 105.94 97.6 106 107.61 ;
      RECT MASK 1 106.214 97.6 106.274 107.61 ;
      RECT MASK 1 106.488 97.6 106.548 107.61 ;
      RECT MASK 1 106.762 97.6 106.822 107.61 ;
      RECT MASK 1 107.036 97.6 107.096 107.61 ;
      RECT MASK 1 107.31 97.6 107.37 107.61 ;
      RECT MASK 1 107.584 97.6 107.644 107.61 ;
      RECT MASK 1 107.858 97.6 107.918 107.61 ;
      RECT MASK 1 108.132 97.6 108.192 107.61 ;
      RECT MASK 1 108.406 97.6 108.466 107.61 ;
      RECT MASK 1 108.68 97.6 108.74 107.61 ;
      RECT MASK 1 108.954 97.6 109.014 107.61 ;
      RECT MASK 1 109.228 97.6 109.288 107.61 ;
      RECT MASK 1 109.502 97.6 109.562 107.61 ;
      RECT MASK 1 109.776 97.6 109.836 107.61 ;
      RECT MASK 1 110.05 97.6 110.11 107.61 ;
      RECT MASK 1 110.324 97.6 110.384 107.61 ;
      RECT MASK 1 110.598 97.6 110.658 107.61 ;
      RECT MASK 1 110.872 97.6 110.932 107.61 ;
      RECT MASK 1 111.146 97.6 111.206 107.61 ;
      RECT MASK 1 111.42 97.6 111.48 107.61 ;
      RECT MASK 1 111.694 97.6 111.754 107.61 ;
      RECT MASK 1 111.968 97.6 112.028 107.61 ;
      RECT MASK 1 112.242 97.6 112.302 107.61 ;
      RECT MASK 1 112.516 97.6 112.576 107.61 ;
      RECT MASK 1 112.79 97.6 112.85 107.61 ;
      RECT MASK 1 113.064 97.6 113.124 107.61 ;
      RECT MASK 1 113.338 97.6 113.398 107.61 ;
      RECT MASK 1 113.612 97.6 113.672 107.61 ;
      RECT MASK 1 113.886 97.6 113.946 107.61 ;
      RECT MASK 1 114.16 97.6 114.22 107.61 ;
      RECT MASK 1 114.434 97.6 114.494 107.61 ;
      RECT MASK 1 114.708 97.6 114.768 107.61 ;
      RECT MASK 1 114.982 97.6 115.042 107.61 ;
      RECT MASK 1 115.256 97.6 115.316 107.61 ;
      RECT MASK 1 115.53 97.6 115.59 107.61 ;
      RECT MASK 1 115.804 97.6 115.864 107.61 ;
      RECT MASK 1 116.078 97.6 116.138 107.61 ;
      RECT MASK 1 116.352 97.6 116.412 107.61 ;
      RECT MASK 1 116.626 97.6 116.686 107.61 ;
      RECT MASK 1 116.9 97.6 116.96 107.61 ;
      RECT MASK 1 117.174 97.6 117.234 107.61 ;
      RECT MASK 1 117.448 97.6 117.508 107.61 ;
      RECT MASK 1 117.722 97.6 117.782 107.61 ;
      RECT MASK 1 117.996 97.6 118.056 107.61 ;
      RECT MASK 1 118.27 97.6 118.33 107.61 ;
      RECT MASK 1 118.544 97.6 118.604 107.61 ;
      RECT MASK 1 118.818 97.6 118.878 107.61 ;
      RECT MASK 1 119.092 97.6 119.152 107.61 ;
      RECT MASK 1 119.366 97.6 119.426 107.61 ;
      RECT MASK 1 119.64 97.6 119.7 107.61 ;
      RECT MASK 1 119.914 97.6 119.974 107.61 ;
      RECT MASK 1 120.188 97.6 120.248 107.61 ;
      RECT MASK 1 120.462 97.6 120.522 107.61 ;
      RECT MASK 1 120.736 97.6 120.796 107.61 ;
      RECT MASK 1 121.01 97.6 121.07 107.61 ;
      RECT MASK 1 121.284 97.6 121.344 107.61 ;
      RECT MASK 1 121.558 97.6 121.618 107.61 ;
      RECT MASK 1 121.832 97.6 121.892 107.61 ;
      RECT MASK 1 122.106 97.6 122.166 107.61 ;
      RECT MASK 1 122.38 97.6 122.44 107.61 ;
      RECT MASK 1 122.654 97.6 122.714 107.61 ;
      RECT MASK 1 122.928 97.6 122.988 107.61 ;
      RECT MASK 1 123.202 97.6 123.262 107.61 ;
      RECT MASK 1 123.476 97.6 123.536 107.61 ;
      RECT MASK 1 123.75 97.6 123.81 107.61 ;
      RECT MASK 1 124.024 97.6 124.084 107.61 ;
      RECT MASK 1 124.298 97.6 124.358 107.61 ;
      RECT MASK 1 124.572 97.6 124.632 107.61 ;
      RECT MASK 1 124.846 97.6 124.906 107.61 ;
      RECT MASK 1 125.12 97.6 125.18 107.61 ;
      RECT MASK 1 125.394 97.6 125.454 107.61 ;
      RECT MASK 1 125.668 97.6 125.728 107.61 ;
      RECT MASK 1 125.942 97.6 126.002 107.61 ;
      RECT MASK 1 126.216 97.6 126.276 107.61 ;
      RECT MASK 1 126.49 97.6 126.55 107.61 ;
      RECT MASK 1 126.764 97.6 126.824 107.61 ;
      RECT MASK 1 127.038 97.6 127.098 107.61 ;
      RECT MASK 1 127.312 97.6 127.372 107.61 ;
      RECT MASK 1 127.586 97.6 127.646 107.66 ;
    LAYER M2 SPACING 0 ;
      RECT 0 0 130.416 109.44 ;
    LAYER M1 SPACING 0 ;
      RECT MASK 2 48.1405 0.584 48.1805 3.1035 ;
      RECT MASK 2 57.849 0.6 57.909 1.5175 ;
      RECT MASK 2 58.536 0.605 58.596 0.835 ;
      RECT MASK 2 60.597 0.605 60.657 0.835 ;
      RECT MASK 2 61.055 0.605 61.115 0.835 ;
      RECT MASK 2 63.574 0.605 63.634 0.835 ;
      RECT MASK 2 64.032 0.605 64.092 0.835 ;
      RECT MASK 2 47.5405 0.784 47.5805 2.65 ;
      RECT MASK 2 48.3405 0.9265 48.3805 2.4895 ;
      RECT MASK 2 50.2985 1.02 50.3385 1.781 ;
      RECT MASK 2 50.9625 1.02 51.0025 1.781 ;
      RECT MASK 2 51.6265 1.02 51.6665 1.781 ;
      RECT MASK 2 52.2905 1.02 52.3305 1.781 ;
      RECT MASK 2 45.7405 1.084 45.7805 2.3865 ;
      RECT MASK 2 59.452 1.16 59.512 2.315 ;
      RECT MASK 2 64.032 1.16 64.092 2.315 ;
      RECT MASK 2 64.49 1.16 64.55 2.315 ;
      RECT MASK 2 58.994 1.165 59.054 2.315 ;
      RECT MASK 2 64.948 1.165 65.008 2.315 ;
      RECT MASK 2 46.3405 1.1845 46.3805 2.644 ;
      RECT MASK 2 61.055 1.198 61.115 1.535 ;
      RECT MASK 2 61.513 1.198 61.573 1.655 ;
      RECT MASK 2 61.971 1.198 62.031 1.54 ;
      RECT MASK 2 62.429 1.198 62.489 1.66 ;
      RECT MASK 2 62.887 1.198 62.947 1.54 ;
      RECT MASK 2 50.0775 1.429 50.1175 7.495 ;
      RECT MASK 2 50.5195 1.429 50.5595 7.975 ;
      RECT MASK 2 50.7415 1.429 50.7815 7.495 ;
      RECT MASK 2 51.1835 1.429 51.2235 7.975 ;
      RECT MASK 2 51.4055 1.429 51.4455 7.495 ;
      RECT MASK 2 51.8475 1.429 51.8875 7.975 ;
      RECT MASK 2 52.0695 1.429 52.1095 7.495 ;
      RECT MASK 2 52.5115 1.429 52.5515 7.975 ;
      RECT MASK 2 2.2785 1.53 2.3385 2.046 ;
      RECT MASK 2 2.6325 1.53 2.6925 2.308 ;
      RECT MASK 2 10.4185 1.53 10.4785 2.4475 ;
      RECT MASK 2 11.2205 1.53 11.2805 7.89 ;
      RECT MASK 2 12.0325 1.53 12.0925 7.89 ;
      RECT MASK 2 12.8445 1.53 12.9045 7.89 ;
      RECT MASK 2 13.6465 1.53 13.7065 2.4475 ;
      RECT MASK 2 33.2305 1.53 33.2905 2.4475 ;
      RECT MASK 2 34.0325 1.53 34.0925 7.89 ;
      RECT MASK 2 34.8445 1.53 34.9045 7.89 ;
      RECT MASK 2 35.6565 1.53 35.7165 7.89 ;
      RECT MASK 2 36.4585 1.53 36.5185 2.4475 ;
      RECT MASK 2 44.2445 1.53 44.3045 2.308 ;
      RECT MASK 2 44.5985 1.53 44.6585 2.046 ;
      RECT MASK 2 1.7055 1.535 1.7655 2.5075 ;
      RECT MASK 2 45.1715 1.535 45.2315 2.5075 ;
      RECT MASK 2 128.073 1.66 128.133 23.64 ;
      RECT MASK 2 116.291 1.68 116.351 23.64 ;
      RECT MASK 2 116.565 1.68 116.625 23.64 ;
      RECT MASK 2 116.839 1.68 116.899 23.64 ;
      RECT MASK 2 117.113 1.68 117.173 23.64 ;
      RECT MASK 2 117.387 1.68 117.447 23.64 ;
      RECT MASK 2 117.661 1.68 117.721 23.64 ;
      RECT MASK 2 117.935 1.68 117.995 23.64 ;
      RECT MASK 2 118.209 1.68 118.269 23.64 ;
      RECT MASK 2 118.483 1.68 118.543 23.64 ;
      RECT MASK 2 118.757 1.68 118.817 23.64 ;
      RECT MASK 2 119.031 1.68 119.091 23.64 ;
      RECT MASK 2 119.305 1.68 119.365 23.64 ;
      RECT MASK 2 119.579 1.68 119.639 23.64 ;
      RECT MASK 2 119.853 1.68 119.913 23.64 ;
      RECT MASK 2 120.127 1.68 120.187 23.64 ;
      RECT MASK 2 120.401 1.68 120.461 23.64 ;
      RECT MASK 2 120.675 1.68 120.735 23.64 ;
      RECT MASK 2 120.949 1.68 121.009 23.64 ;
      RECT MASK 2 121.223 1.68 121.283 23.64 ;
      RECT MASK 2 121.497 1.68 121.557 23.64 ;
      RECT MASK 2 121.771 1.68 121.831 23.64 ;
      RECT MASK 2 122.045 1.68 122.105 23.64 ;
      RECT MASK 2 122.319 1.68 122.379 23.64 ;
      RECT MASK 2 122.593 1.68 122.653 23.64 ;
      RECT MASK 2 122.867 1.68 122.927 23.64 ;
      RECT MASK 2 123.141 1.68 123.201 23.64 ;
      RECT MASK 2 123.415 1.68 123.475 23.64 ;
      RECT MASK 2 123.689 1.68 123.749 23.64 ;
      RECT MASK 2 123.963 1.68 124.023 23.64 ;
      RECT MASK 2 124.237 1.68 124.297 23.64 ;
      RECT MASK 2 124.511 1.68 124.571 23.64 ;
      RECT MASK 2 124.785 1.68 124.845 23.64 ;
      RECT MASK 2 125.059 1.68 125.119 23.64 ;
      RECT MASK 2 125.333 1.68 125.393 23.64 ;
      RECT MASK 2 125.607 1.68 125.667 23.64 ;
      RECT MASK 2 125.881 1.68 125.941 23.64 ;
      RECT MASK 2 126.155 1.68 126.215 23.64 ;
      RECT MASK 2 126.429 1.68 126.489 23.64 ;
      RECT MASK 2 126.703 1.68 126.763 23.64 ;
      RECT MASK 2 126.977 1.68 127.037 23.64 ;
      RECT MASK 2 127.251 1.68 127.311 23.64 ;
      RECT MASK 2 127.525 1.68 127.585 23.64 ;
      RECT MASK 2 127.799 1.68 127.859 23.64 ;
      RECT MASK 2 22.2385 1.8 22.2985 2.561 ;
      RECT MASK 2 23.2385 1.8 23.2985 2.561 ;
      RECT MASK 2 23.6385 1.8 23.6985 2.561 ;
      RECT MASK 2 24.6385 1.8 24.6985 2.561 ;
      RECT MASK 2 22.4385 1.815 22.4985 2.025 ;
      RECT MASK 2 22.6385 1.815 22.6985 2.414 ;
      RECT MASK 2 22.8385 1.815 22.8985 2.561 ;
      RECT MASK 2 23.0385 1.815 23.0985 2.025 ;
      RECT MASK 2 23.8385 1.815 23.8985 2.025 ;
      RECT MASK 2 24.0385 1.815 24.0985 2.561 ;
      RECT MASK 2 24.2385 1.815 24.2985 2.414 ;
      RECT MASK 2 24.4385 1.815 24.4985 2.025 ;
      RECT MASK 2 50.2985 1.819 50.3385 6.57 ;
      RECT MASK 2 50.9625 1.819 51.0025 6.57 ;
      RECT MASK 2 51.6265 1.819 51.6665 6.57 ;
      RECT MASK 2 52.2905 1.819 52.3305 6.57 ;
      RECT MASK 2 62.429 1.82 62.489 2.282 ;
      RECT MASK 2 61.513 1.825 61.573 2.282 ;
      RECT MASK 2 61.971 1.94 62.031 2.282 ;
      RECT MASK 2 62.887 1.94 62.947 2.282 ;
      RECT MASK 2 61.055 1.945 61.115 2.282 ;
      RECT MASK 2 57.849 1.9625 57.909 3.0775 ;
      RECT MASK 2 65.864 2.0825 65.924 3.138 ;
      RECT MASK 2 10.9705 2.09 11.0305 2.811 ;
      RECT MASK 2 12.4905 2.09 12.5505 2.308 ;
      RECT MASK 2 14.8025 2.09 14.8625 2.308 ;
      RECT MASK 2 15.2605 2.09 15.3205 2.308 ;
      RECT MASK 2 15.7185 2.09 15.7785 2.308 ;
      RECT MASK 2 16.1765 2.09 16.2365 2.308 ;
      RECT MASK 2 16.6345 2.09 16.6945 2.308 ;
      RECT MASK 2 17.0925 2.09 17.1525 2.308 ;
      RECT MASK 2 17.5505 2.09 17.6105 2.308 ;
      RECT MASK 2 18.0085 2.09 18.0685 2.308 ;
      RECT MASK 2 18.4665 2.09 18.5265 2.308 ;
      RECT MASK 2 18.9245 2.09 18.9845 2.308 ;
      RECT MASK 2 19.3825 2.09 19.4425 2.308 ;
      RECT MASK 2 19.8405 2.09 19.9005 2.308 ;
      RECT MASK 2 20.2985 2.09 20.3585 2.308 ;
      RECT MASK 2 20.7565 2.09 20.8165 2.308 ;
      RECT MASK 2 26.1205 2.09 26.1805 2.308 ;
      RECT MASK 2 26.5785 2.09 26.6385 2.308 ;
      RECT MASK 2 27.0365 2.09 27.0965 2.308 ;
      RECT MASK 2 27.4945 2.09 27.5545 2.308 ;
      RECT MASK 2 27.9525 2.09 28.0125 2.308 ;
      RECT MASK 2 28.4105 2.09 28.4705 2.308 ;
      RECT MASK 2 28.8685 2.09 28.9285 2.308 ;
      RECT MASK 2 29.3265 2.09 29.3865 2.308 ;
      RECT MASK 2 29.7845 2.09 29.8445 2.308 ;
      RECT MASK 2 30.2425 2.09 30.3025 2.308 ;
      RECT MASK 2 30.7005 2.09 30.7605 2.308 ;
      RECT MASK 2 31.1585 2.09 31.2185 2.308 ;
      RECT MASK 2 31.6165 2.09 31.6765 2.308 ;
      RECT MASK 2 32.0745 2.09 32.1345 2.308 ;
      RECT MASK 2 34.3865 2.09 34.4465 2.308 ;
      RECT MASK 2 35.9065 2.09 35.9665 2.811 ;
      RECT MASK 2 46.9405 2.09 46.9805 2.65 ;
      RECT MASK 2 47.1405 2.09 47.1805 2.65 ;
      RECT MASK 2 47.3405 2.09 47.3805 2.65 ;
      RECT MASK 2 47.7405 2.09 47.7805 2.65 ;
      RECT MASK 2 47.9405 2.09 47.9805 2.65 ;
      RECT MASK 2 21.2145 2.095 21.2745 2.308 ;
      RECT MASK 2 25.6625 2.095 25.7225 2.308 ;
      RECT MASK 2 11.5745 2.128 11.6345 2.405 ;
      RECT MASK 2 35.3025 2.128 35.3625 2.405 ;
      RECT MASK 2 22.4385 2.21 22.4985 3.175 ;
      RECT MASK 2 23.0385 2.21 23.0985 3.175 ;
      RECT MASK 2 23.8385 2.21 23.8985 3.175 ;
      RECT MASK 2 24.4385 2.21 24.4985 3.175 ;
      RECT MASK 2 3.4235 2.428 3.4835 2.912 ;
      RECT MASK 2 10.1025 2.428 10.1625 2.645 ;
      RECT MASK 2 36.7745 2.428 36.8345 2.645 ;
      RECT MASK 2 43.4535 2.428 43.5135 2.912 ;
      RECT MASK 2 61.284 2.435 61.344 3.6775 ;
      RECT MASK 2 62.658 2.438 62.718 2.938 ;
      RECT MASK 2 63.116 2.438 63.176 2.938 ;
      RECT MASK 2 63.574 2.438 63.634 2.938 ;
      RECT MASK 2 64.032 2.438 64.092 2.938 ;
      RECT MASK 2 64.49 2.438 64.55 2.938 ;
      RECT MASK 2 64.948 2.438 65.008 2.938 ;
      RECT MASK 2 65.406 2.438 65.466 2.938 ;
      RECT MASK 2 5.5145 2.45 5.5745 2.811 ;
      RECT MASK 2 5.7305 2.45 5.7905 2.811 ;
      RECT MASK 2 6.4215 2.45 6.4815 2.811 ;
      RECT MASK 2 6.6335 2.45 6.6935 2.811 ;
      RECT MASK 2 7.3375 2.45 7.3975 2.811 ;
      RECT MASK 2 7.5495 2.45 7.6095 2.811 ;
      RECT MASK 2 8.2495 2.45 8.3095 2.811 ;
      RECT MASK 2 8.4615 2.45 8.5215 2.811 ;
      RECT MASK 2 38.4155 2.45 38.4755 2.811 ;
      RECT MASK 2 38.6275 2.45 38.6875 2.811 ;
      RECT MASK 2 39.3275 2.45 39.3875 2.811 ;
      RECT MASK 2 39.5395 2.45 39.5995 2.811 ;
      RECT MASK 2 40.2435 2.45 40.3035 2.811 ;
      RECT MASK 2 40.4555 2.45 40.5155 2.811 ;
      RECT MASK 2 41.1465 2.45 41.2065 2.811 ;
      RECT MASK 2 41.3625 2.45 41.4225 2.811 ;
      RECT MASK 2 17.894 2.47 17.954 2.65 ;
      RECT MASK 2 19.268 2.47 19.328 2.65 ;
      RECT MASK 2 20.184 2.47 20.244 2.65 ;
      RECT MASK 2 26.693 2.47 26.753 2.65 ;
      RECT MASK 2 27.609 2.47 27.669 2.65 ;
      RECT MASK 2 28.983 2.47 29.043 2.65 ;
      RECT MASK 2 2.6325 2.529 2.6925 2.811 ;
      RECT MASK 2 44.2445 2.529 44.3045 2.811 ;
      RECT MASK 2 22.6385 2.645 22.6985 2.785 ;
      RECT MASK 2 24.2385 2.645 24.2985 2.785 ;
      RECT MASK 2 17.207 2.69 17.267 2.87 ;
      RECT MASK 2 18.581 2.69 18.641 2.87 ;
      RECT MASK 2 28.296 2.69 28.356 2.87 ;
      RECT MASK 2 29.67 2.69 29.73 2.87 ;
      RECT MASK 2 58.765 2.725 58.825 2.938 ;
      RECT MASK 2 59.223 2.725 59.283 2.938 ;
      RECT MASK 2 59.681 2.725 59.741 2.938 ;
      RECT MASK 2 60.139 2.725 60.199 2.938 ;
      RECT MASK 2 22.2385 2.794 22.2985 3.54 ;
      RECT MASK 2 22.8385 2.794 22.8985 3.54 ;
      RECT MASK 2 23.2385 2.794 23.2985 3.54 ;
      RECT MASK 2 23.6385 2.794 23.6985 3.54 ;
      RECT MASK 2 24.0385 2.794 24.0985 3.54 ;
      RECT MASK 2 24.6385 2.794 24.6985 3.54 ;
      RECT MASK 2 46.9405 2.81 46.9805 3.37 ;
      RECT MASK 2 47.1405 2.81 47.1805 3.37 ;
      RECT MASK 2 47.3405 2.81 47.3805 3.37 ;
      RECT MASK 2 47.5405 2.81 47.5805 3.37 ;
      RECT MASK 2 47.7405 2.81 47.7805 3.37 ;
      RECT MASK 2 47.9405 2.81 47.9805 3.37 ;
      RECT MASK 2 12.9915 2.832 13.0515 3.245 ;
      RECT MASK 2 33.8855 2.832 33.9455 3.245 ;
      RECT MASK 2 1.7055 2.8325 1.7655 4.5475 ;
      RECT MASK 2 45.1715 2.8325 45.2315 4.5475 ;
      RECT MASK 2 10.4185 2.8925 10.4785 4.4875 ;
      RECT MASK 2 13.6465 2.8925 13.7065 4.4875 ;
      RECT MASK 2 33.2305 2.8925 33.2905 4.4875 ;
      RECT MASK 2 36.4585 2.8925 36.5185 4.4875 ;
      RECT MASK 2 22.6385 2.941 22.6985 3.54 ;
      RECT MASK 2 24.2385 2.941 24.2985 3.54 ;
      RECT MASK 2 2.6325 3.032 2.6925 4.348 ;
      RECT MASK 2 11.5745 3.032 11.6345 3.25 ;
      RECT MASK 2 12.4905 3.032 12.5505 3.245 ;
      RECT MASK 2 14.8025 3.032 14.8625 3.25 ;
      RECT MASK 2 15.2605 3.032 15.3205 3.25 ;
      RECT MASK 2 15.7185 3.032 15.7785 3.25 ;
      RECT MASK 2 16.1765 3.032 16.2365 3.25 ;
      RECT MASK 2 16.6345 3.032 16.6945 3.25 ;
      RECT MASK 2 17.0925 3.032 17.1525 3.25 ;
      RECT MASK 2 17.5505 3.032 17.6105 3.25 ;
      RECT MASK 2 18.0085 3.032 18.0685 3.25 ;
      RECT MASK 2 18.4665 3.032 18.5265 3.25 ;
      RECT MASK 2 18.9245 3.032 18.9845 3.25 ;
      RECT MASK 2 19.3825 3.032 19.4425 3.25 ;
      RECT MASK 2 19.8405 3.032 19.9005 3.25 ;
      RECT MASK 2 20.2985 3.032 20.3585 3.25 ;
      RECT MASK 2 20.7565 3.032 20.8165 3.25 ;
      RECT MASK 2 21.2145 3.032 21.2745 3.245 ;
      RECT MASK 2 25.6625 3.032 25.7225 3.245 ;
      RECT MASK 2 26.1205 3.032 26.1805 3.25 ;
      RECT MASK 2 26.5785 3.032 26.6385 3.25 ;
      RECT MASK 2 27.0365 3.032 27.0965 3.25 ;
      RECT MASK 2 27.4945 3.032 27.5545 3.25 ;
      RECT MASK 2 27.9525 3.032 28.0125 3.25 ;
      RECT MASK 2 28.4105 3.032 28.4705 3.25 ;
      RECT MASK 2 28.8685 3.032 28.9285 3.25 ;
      RECT MASK 2 29.3265 3.032 29.3865 3.25 ;
      RECT MASK 2 29.7845 3.032 29.8445 3.25 ;
      RECT MASK 2 30.2425 3.032 30.3025 3.25 ;
      RECT MASK 2 30.7005 3.032 30.7605 3.25 ;
      RECT MASK 2 31.1585 3.032 31.2185 3.25 ;
      RECT MASK 2 31.6165 3.032 31.6765 3.25 ;
      RECT MASK 2 32.0745 3.032 32.1345 3.25 ;
      RECT MASK 2 34.3865 3.032 34.4465 3.245 ;
      RECT MASK 2 35.3025 3.032 35.3625 3.25 ;
      RECT MASK 2 44.2445 3.032 44.3045 4.353 ;
      RECT MASK 2 62.658 3.058 62.718 3.542 ;
      RECT MASK 2 65.406 3.085 65.466 3.441 ;
      RECT MASK 2 59.3375 3.159 59.3975 3.4525 ;
      RECT MASK 2 64.719 3.159 64.779 3.4 ;
      RECT MASK 2 64.032 3.205 64.092 3.842 ;
      RECT MASK 2 48.1405 3.235 48.1805 3.993 ;
      RECT MASK 2 2.2785 3.294 2.3385 4.086 ;
      RECT MASK 2 44.5985 3.294 44.6585 4.086 ;
      RECT MASK 2 62.31 3.325 62.37 3.633 ;
      RECT MASK 2 64.948 3.325 65.008 3.842 ;
      RECT MASK 2 22.4385 3.33 22.4985 3.54 ;
      RECT MASK 2 23.0385 3.33 23.0985 3.54 ;
      RECT MASK 2 23.8385 3.33 23.8985 3.54 ;
      RECT MASK 2 24.4385 3.33 24.4985 3.54 ;
      RECT MASK 2 56.4115 3.3435 56.4715 6.179 ;
      RECT MASK 2 58.765 3.361 58.825 4.799 ;
      RECT MASK 2 60.139 3.361 60.199 4.799 ;
      RECT MASK 2 66.7185 3.445 66.7785 9.557 ;
      RECT MASK 2 57.849 3.5225 57.909 4.6375 ;
      RECT MASK 2 46.9405 3.53 46.9805 4.09 ;
      RECT MASK 2 47.1405 3.53 47.1805 4.09 ;
      RECT MASK 2 47.3405 3.53 47.3805 4.09 ;
      RECT MASK 2 47.5405 3.53 47.5805 4.09 ;
      RECT MASK 2 47.7405 3.53 47.7805 4.09 ;
      RECT MASK 2 47.9405 3.53 47.9805 4.09 ;
      RECT MASK 2 76.8795 3.54 76.9795 8.8515 ;
      RECT MASK 2 77.4435 3.54 77.5435 10.5615 ;
      RECT MASK 2 109.1615 3.54 109.2615 10.5615 ;
      RECT MASK 2 109.7255 3.54 109.8255 8.8515 ;
      RECT MASK 2 59.223 3.662 59.283 3.88 ;
      RECT MASK 2 59.681 3.662 59.741 3.88 ;
      RECT MASK 2 62.628 3.662 62.748 4.498 ;
      RECT MASK 2 63.086 3.662 63.206 4.498 ;
      RECT MASK 2 63.544 3.662 63.664 4.498 ;
      RECT MASK 2 64.46 3.662 64.58 4.498 ;
      RECT MASK 2 65.406 3.662 65.466 4.498 ;
      RECT MASK 2 65.864 3.662 65.924 4.498 ;
      RECT MASK 2 83.7935 3.78 83.8935 6.5715 ;
      RECT MASK 2 84.1285 3.78 84.2285 6.603 ;
      RECT MASK 2 91.4325 3.78 91.5325 6.54 ;
      RECT MASK 2 95.1725 3.78 95.2725 6.54 ;
      RECT MASK 2 102.4765 3.78 102.5765 6.603 ;
      RECT MASK 2 102.8115 3.78 102.9115 6.5715 ;
      RECT MASK 2 22.2385 3.84 22.2985 4.586 ;
      RECT MASK 2 22.4385 3.84 22.4985 4.05 ;
      RECT MASK 2 22.6385 3.84 22.6985 4.439 ;
      RECT MASK 2 22.8385 3.84 22.8985 4.586 ;
      RECT MASK 2 23.0385 3.84 23.0985 4.05 ;
      RECT MASK 2 23.2385 3.84 23.2985 4.586 ;
      RECT MASK 2 23.6385 3.84 23.6985 4.586 ;
      RECT MASK 2 23.8385 3.84 23.8985 4.05 ;
      RECT MASK 2 24.0385 3.84 24.0985 4.586 ;
      RECT MASK 2 24.2385 3.84 24.2985 4.439 ;
      RECT MASK 2 24.4385 3.84 24.4985 4.05 ;
      RECT MASK 2 24.6385 3.84 24.6985 4.586 ;
      RECT MASK 2 11.5745 4.13 11.6345 4.348 ;
      RECT MASK 2 14.8025 4.13 14.8625 4.348 ;
      RECT MASK 2 15.2605 4.13 15.3205 4.348 ;
      RECT MASK 2 15.7185 4.13 15.7785 4.348 ;
      RECT MASK 2 16.1765 4.13 16.2365 4.348 ;
      RECT MASK 2 16.6345 4.13 16.6945 4.348 ;
      RECT MASK 2 17.0925 4.13 17.1525 4.348 ;
      RECT MASK 2 17.5505 4.13 17.6105 4.348 ;
      RECT MASK 2 18.0085 4.13 18.0685 4.348 ;
      RECT MASK 2 18.4665 4.13 18.5265 4.348 ;
      RECT MASK 2 18.9245 4.13 18.9845 4.348 ;
      RECT MASK 2 19.3825 4.13 19.4425 4.348 ;
      RECT MASK 2 19.8405 4.13 19.9005 4.348 ;
      RECT MASK 2 20.2985 4.13 20.3585 4.348 ;
      RECT MASK 2 20.7565 4.13 20.8165 4.348 ;
      RECT MASK 2 26.1205 4.13 26.1805 4.348 ;
      RECT MASK 2 26.5785 4.13 26.6385 4.348 ;
      RECT MASK 2 27.0365 4.13 27.0965 4.348 ;
      RECT MASK 2 27.4945 4.13 27.5545 4.348 ;
      RECT MASK 2 27.9525 4.13 28.0125 4.348 ;
      RECT MASK 2 28.4105 4.13 28.4705 4.348 ;
      RECT MASK 2 28.8685 4.13 28.9285 4.348 ;
      RECT MASK 2 29.3265 4.13 29.3865 4.348 ;
      RECT MASK 2 29.7845 4.13 29.8445 4.348 ;
      RECT MASK 2 30.2425 4.13 30.3025 4.348 ;
      RECT MASK 2 30.7005 4.13 30.7605 4.348 ;
      RECT MASK 2 31.1585 4.13 31.2185 4.348 ;
      RECT MASK 2 31.6165 4.13 31.6765 4.348 ;
      RECT MASK 2 32.0745 4.13 32.1345 4.348 ;
      RECT MASK 2 35.3025 4.13 35.3625 4.348 ;
      RECT MASK 2 12.4905 4.135 12.5505 4.348 ;
      RECT MASK 2 12.9915 4.135 13.0515 4.548 ;
      RECT MASK 2 21.2145 4.135 21.2745 4.348 ;
      RECT MASK 2 25.6625 4.135 25.7225 4.348 ;
      RECT MASK 2 33.8855 4.135 33.9455 4.548 ;
      RECT MASK 2 34.3865 4.135 34.4465 4.348 ;
      RECT MASK 2 22.4385 4.205 22.4985 5.17 ;
      RECT MASK 2 23.0385 4.205 23.0985 5.17 ;
      RECT MASK 2 23.8385 4.205 23.8985 5.17 ;
      RECT MASK 2 24.4385 4.205 24.4985 5.17 ;
      RECT MASK 2 59.223 4.28 59.283 4.498 ;
      RECT MASK 2 59.681 4.28 59.741 4.498 ;
      RECT MASK 2 64.032 4.318 64.092 4.955 ;
      RECT MASK 2 64.948 4.318 65.008 4.835 ;
      RECT MASK 2 3.4235 4.468 3.4835 4.952 ;
      RECT MASK 2 43.4535 4.468 43.5135 4.952 ;
      RECT MASK 2 61.284 4.4825 61.344 5.725 ;
      RECT MASK 2 85.1245 4.488 85.2245 5.168 ;
      RECT MASK 2 86.1205 4.488 86.2205 5.168 ;
      RECT MASK 2 87.1165 4.488 87.2165 5.168 ;
      RECT MASK 2 88.7765 4.488 88.8765 5.168 ;
      RECT MASK 2 89.7725 4.488 89.8725 5.168 ;
      RECT MASK 2 90.7685 4.488 90.8685 5.168 ;
      RECT MASK 2 91.7645 4.488 91.8645 5.168 ;
      RECT MASK 2 94.8405 4.488 94.9405 5.168 ;
      RECT MASK 2 95.8365 4.488 95.9365 5.168 ;
      RECT MASK 2 96.8325 4.488 96.9325 5.168 ;
      RECT MASK 2 97.8285 4.488 97.9285 5.168 ;
      RECT MASK 2 99.4885 4.488 99.5885 5.168 ;
      RECT MASK 2 100.4845 4.488 100.5845 5.168 ;
      RECT MASK 2 101.4805 4.488 101.5805 5.168 ;
      RECT MASK 2 17.207 4.51 17.267 4.69 ;
      RECT MASK 2 18.581 4.51 18.641 4.69 ;
      RECT MASK 2 28.296 4.51 28.356 4.69 ;
      RECT MASK 2 29.67 4.51 29.73 4.69 ;
      RECT MASK 2 86.7845 4.557 86.8845 5.889 ;
      RECT MASK 2 87.7805 4.557 87.8805 5.889 ;
      RECT MASK 2 98.8245 4.557 98.9245 5.889 ;
      RECT MASK 2 99.8205 4.557 99.9205 5.889 ;
      RECT MASK 2 2.6325 4.569 2.6925 4.851 ;
      RECT MASK 2 5.5145 4.569 5.5745 4.93 ;
      RECT MASK 2 5.7305 4.569 5.7905 4.93 ;
      RECT MASK 2 6.4215 4.569 6.4815 4.93 ;
      RECT MASK 2 6.6335 4.569 6.6935 4.93 ;
      RECT MASK 2 7.3375 4.569 7.3975 4.93 ;
      RECT MASK 2 7.5495 4.569 7.6095 4.93 ;
      RECT MASK 2 8.2495 4.569 8.3095 4.93 ;
      RECT MASK 2 8.4615 4.569 8.5215 4.93 ;
      RECT MASK 2 10.9705 4.569 11.0305 5.29 ;
      RECT MASK 2 35.9065 4.569 35.9665 5.29 ;
      RECT MASK 2 38.4155 4.569 38.4755 4.93 ;
      RECT MASK 2 38.6275 4.569 38.6875 4.93 ;
      RECT MASK 2 39.3275 4.569 39.3875 4.93 ;
      RECT MASK 2 39.5395 4.569 39.5995 4.93 ;
      RECT MASK 2 40.2435 4.569 40.3035 4.93 ;
      RECT MASK 2 40.4555 4.569 40.5155 4.93 ;
      RECT MASK 2 41.1465 4.569 41.2065 4.93 ;
      RECT MASK 2 41.3625 4.569 41.4225 4.93 ;
      RECT MASK 2 44.2445 4.569 44.3045 4.851 ;
      RECT MASK 2 22.6385 4.595 22.6985 4.735 ;
      RECT MASK 2 24.2385 4.595 24.2985 4.735 ;
      RECT MASK 2 84.7925 4.609 84.8925 6.625 ;
      RECT MASK 2 85.7885 4.609 85.8885 6.625 ;
      RECT MASK 2 89.4405 4.609 89.5405 5.289 ;
      RECT MASK 2 97.1645 4.609 97.2645 5.289 ;
      RECT MASK 2 100.8165 4.609 100.9165 6.625 ;
      RECT MASK 2 101.8125 4.609 101.9125 6.625 ;
      RECT MASK 2 62.658 4.618 62.718 5.102 ;
      RECT MASK 2 56.842 4.645 56.902 7.3035 ;
      RECT MASK 2 59.3375 4.7075 59.3975 5.001 ;
      RECT MASK 2 65.406 4.719 65.466 5.075 ;
      RECT MASK 2 88.4445 4.7235 88.5045 6.54 ;
      RECT MASK 2 98.2005 4.7235 98.2605 6.54 ;
      RECT MASK 2 17.894 4.73 17.954 4.91 ;
      RECT MASK 2 19.268 4.73 19.328 4.91 ;
      RECT MASK 2 20.184 4.73 20.244 4.91 ;
      RECT MASK 2 26.693 4.73 26.753 4.91 ;
      RECT MASK 2 27.609 4.73 27.669 4.91 ;
      RECT MASK 2 28.983 4.73 29.043 4.91 ;
      RECT MASK 2 85.4565 4.73 85.5565 5.41 ;
      RECT MASK 2 86.4525 4.73 86.5525 5.41 ;
      RECT MASK 2 87.4485 4.73 87.5485 5.41 ;
      RECT MASK 2 89.1085 4.73 89.2085 5.41 ;
      RECT MASK 2 90.1045 4.73 90.2045 5.4165 ;
      RECT MASK 2 91.1005 4.73 91.2005 5.4165 ;
      RECT MASK 2 92.0965 4.73 92.1965 5.4165 ;
      RECT MASK 2 94.5085 4.73 94.6085 5.4165 ;
      RECT MASK 2 95.5045 4.73 95.6045 5.4165 ;
      RECT MASK 2 96.5005 4.73 96.6005 5.4165 ;
      RECT MASK 2 97.4965 4.73 97.5965 5.41 ;
      RECT MASK 2 99.1565 4.73 99.2565 5.41 ;
      RECT MASK 2 100.1525 4.73 100.2525 5.41 ;
      RECT MASK 2 101.1485 4.73 101.2485 5.41 ;
      RECT MASK 2 10.1025 4.735 10.1625 4.952 ;
      RECT MASK 2 36.7745 4.735 36.8345 4.952 ;
      RECT MASK 2 64.719 4.76 64.779 5.001 ;
      RECT MASK 2 22.2385 4.819 22.2985 5.58 ;
      RECT MASK 2 22.8385 4.819 22.8985 5.565 ;
      RECT MASK 2 23.2385 4.819 23.2985 5.58 ;
      RECT MASK 2 23.6385 4.819 23.6985 5.58 ;
      RECT MASK 2 24.0385 4.819 24.0985 5.565 ;
      RECT MASK 2 24.6385 4.819 24.6985 5.58 ;
      RECT MASK 2 1.7055 4.8725 1.7655 6.5875 ;
      RECT MASK 2 45.1715 4.8725 45.2315 6.5875 ;
      RECT MASK 2 10.4185 4.9325 10.4785 6.5275 ;
      RECT MASK 2 13.6465 4.9325 13.7065 6.5275 ;
      RECT MASK 2 33.2305 4.9325 33.2905 6.5275 ;
      RECT MASK 2 36.4585 4.9325 36.5185 6.5275 ;
      RECT MASK 2 22.6385 4.966 22.6985 5.565 ;
      RECT MASK 2 24.2385 4.966 24.2985 5.565 ;
      RECT MASK 2 11.5745 4.975 11.6345 5.252 ;
      RECT MASK 2 35.3025 4.975 35.3625 5.252 ;
      RECT MASK 2 65.864 5.022 65.924 6.0775 ;
      RECT MASK 2 2.6325 5.072 2.6925 6.388 ;
      RECT MASK 2 12.4905 5.072 12.5505 5.29 ;
      RECT MASK 2 14.8025 5.072 14.8625 5.29 ;
      RECT MASK 2 15.2605 5.072 15.3205 5.29 ;
      RECT MASK 2 15.7185 5.072 15.7785 5.29 ;
      RECT MASK 2 16.1765 5.072 16.2365 5.29 ;
      RECT MASK 2 16.6345 5.072 16.6945 5.29 ;
      RECT MASK 2 17.0925 5.072 17.1525 5.29 ;
      RECT MASK 2 17.5505 5.072 17.6105 5.29 ;
      RECT MASK 2 18.0085 5.072 18.0685 5.29 ;
      RECT MASK 2 18.4665 5.072 18.5265 5.29 ;
      RECT MASK 2 18.9245 5.072 18.9845 5.29 ;
      RECT MASK 2 19.3825 5.072 19.4425 5.29 ;
      RECT MASK 2 19.8405 5.072 19.9005 5.29 ;
      RECT MASK 2 20.2985 5.072 20.3585 5.29 ;
      RECT MASK 2 20.7565 5.072 20.8165 5.29 ;
      RECT MASK 2 21.2145 5.072 21.2745 5.285 ;
      RECT MASK 2 25.6625 5.072 25.7225 5.285 ;
      RECT MASK 2 26.1205 5.072 26.1805 5.29 ;
      RECT MASK 2 26.5785 5.072 26.6385 5.29 ;
      RECT MASK 2 27.0365 5.072 27.0965 5.29 ;
      RECT MASK 2 27.4945 5.072 27.5545 5.29 ;
      RECT MASK 2 27.9525 5.072 28.0125 5.29 ;
      RECT MASK 2 28.4105 5.072 28.4705 5.29 ;
      RECT MASK 2 28.8685 5.072 28.9285 5.29 ;
      RECT MASK 2 29.3265 5.072 29.3865 5.29 ;
      RECT MASK 2 29.7845 5.072 29.8445 5.29 ;
      RECT MASK 2 30.2425 5.072 30.3025 5.29 ;
      RECT MASK 2 30.7005 5.072 30.7605 5.29 ;
      RECT MASK 2 31.1585 5.072 31.2185 5.29 ;
      RECT MASK 2 31.6165 5.072 31.6765 5.29 ;
      RECT MASK 2 32.0745 5.072 32.1345 5.29 ;
      RECT MASK 2 34.3865 5.072 34.4465 5.29 ;
      RECT MASK 2 44.2445 5.072 44.3045 6.388 ;
      RECT MASK 2 57.849 5.0825 57.909 6.1975 ;
      RECT MASK 2 46.9655 5.135 47.0255 5.606 ;
      RECT MASK 2 47.2975 5.135 47.3575 5.606 ;
      RECT MASK 2 47.6295 5.135 47.6895 5.786 ;
      RECT MASK 2 47.9615 5.135 48.0215 5.781 ;
      RECT MASK 2 48.2935 5.135 48.3535 5.781 ;
      RECT MASK 2 48.6255 5.135 48.6855 5.781 ;
      RECT MASK 2 58.765 5.222 58.825 5.435 ;
      RECT MASK 2 59.223 5.222 59.283 5.435 ;
      RECT MASK 2 59.681 5.222 59.741 5.435 ;
      RECT MASK 2 60.139 5.222 60.199 5.435 ;
      RECT MASK 2 62.658 5.222 62.718 5.722 ;
      RECT MASK 2 63.116 5.222 63.176 5.722 ;
      RECT MASK 2 63.574 5.222 63.634 5.722 ;
      RECT MASK 2 64.032 5.222 64.092 5.722 ;
      RECT MASK 2 64.49 5.222 64.55 5.722 ;
      RECT MASK 2 64.948 5.222 65.008 5.722 ;
      RECT MASK 2 65.406 5.222 65.466 5.722 ;
      RECT MASK 2 54.1785 5.255 54.2385 5.901 ;
      RECT MASK 2 54.5105 5.255 54.5705 5.726 ;
      RECT MASK 2 55.0085 5.255 55.0685 5.901 ;
      RECT MASK 2 55.6725 5.255 55.7325 5.901 ;
      RECT MASK 2 2.2785 5.334 2.3385 6.126 ;
      RECT MASK 2 44.5985 5.334 44.6585 6.126 ;
      RECT MASK 2 22.4385 5.355 22.4985 5.565 ;
      RECT MASK 2 23.0385 5.355 23.0985 5.565 ;
      RECT MASK 2 23.8385 5.355 23.8985 5.565 ;
      RECT MASK 2 24.4385 5.355 24.4985 5.565 ;
      RECT MASK 2 87.1165 5.6585 87.2165 7.891 ;
      RECT MASK 2 99.4885 5.6585 99.5885 7.891 ;
      RECT MASK 2 89.1345 5.673 89.1945 6.54 ;
      RECT MASK 2 89.7045 5.673 89.7645 6.54 ;
      RECT MASK 2 89.9565 5.673 90.0165 6.54 ;
      RECT MASK 2 90.4545 5.673 90.5145 6.54 ;
      RECT MASK 2 96.1905 5.673 96.2505 6.54 ;
      RECT MASK 2 96.6885 5.673 96.7485 6.54 ;
      RECT MASK 2 96.9405 5.673 97.0005 6.54 ;
      RECT MASK 2 97.5105 5.673 97.5705 6.54 ;
      RECT MASK 2 87.4485 5.68 87.5485 6.55 ;
      RECT MASK 2 99.1565 5.68 99.2565 6.55 ;
      RECT MASK 2 88.1925 5.688 88.2525 6.54 ;
      RECT MASK 2 98.4525 5.688 98.5125 6.54 ;
      RECT MASK 2 90.2085 5.7285 90.2685 7.721 ;
      RECT MASK 2 96.4365 5.7285 96.4965 7.721 ;
      RECT MASK 2 88.8935 5.7565 88.9535 7.6 ;
      RECT MASK 2 97.7515 5.7565 97.8115 7.6 ;
      RECT MASK 2 46.9655 5.798 47.0255 6.622 ;
      RECT MASK 2 47.2975 5.798 47.3575 6.622 ;
      RECT MASK 2 90.9645 5.8 91.0245 7.721 ;
      RECT MASK 2 95.6805 5.8 95.7405 9.658 ;
      RECT MASK 2 58.994 5.845 59.054 6.995 ;
      RECT MASK 2 59.452 5.845 59.512 7 ;
      RECT MASK 2 64.032 5.845 64.092 7 ;
      RECT MASK 2 64.49 5.845 64.55 7 ;
      RECT MASK 2 64.948 5.845 65.008 6.995 ;
      RECT MASK 2 90.708 5.8565 90.768 7.6 ;
      RECT MASK 2 95.937 5.8565 95.997 7.6 ;
      RECT MASK 2 61.055 5.878 61.115 6.215 ;
      RECT MASK 2 61.513 5.878 61.573 6.335 ;
      RECT MASK 2 61.971 5.878 62.031 6.22 ;
      RECT MASK 2 62.429 5.878 62.489 6.34 ;
      RECT MASK 2 62.887 5.878 62.947 6.22 ;
      RECT MASK 2 22.2385 5.88 22.2985 6.641 ;
      RECT MASK 2 23.2385 5.88 23.2985 6.641 ;
      RECT MASK 2 23.6385 5.88 23.6985 6.641 ;
      RECT MASK 2 24.6385 5.88 24.6985 6.641 ;
      RECT MASK 2 22.4385 5.895 22.4985 6.105 ;
      RECT MASK 2 22.6385 5.895 22.6985 6.494 ;
      RECT MASK 2 22.8385 5.895 22.8985 6.641 ;
      RECT MASK 2 23.0385 5.895 23.0985 6.105 ;
      RECT MASK 2 23.8385 5.895 23.8985 6.105 ;
      RECT MASK 2 24.0385 5.895 24.0985 6.641 ;
      RECT MASK 2 24.2385 5.895 24.2985 6.494 ;
      RECT MASK 2 24.4385 5.895 24.4985 6.105 ;
      RECT MASK 2 89.3755 5.909 89.4355 7.6 ;
      RECT MASK 2 97.2695 5.909 97.3295 7.6 ;
      RECT MASK 2 54.5105 5.918 54.5705 6.742 ;
      RECT MASK 2 55.3405 5.918 55.4005 6.742 ;
      RECT MASK 2 85.4565 5.93 85.5565 7.6 ;
      RECT MASK 2 86.1205 5.93 86.2205 7.6 ;
      RECT MASK 2 100.4845 5.93 100.5845 7.6 ;
      RECT MASK 2 101.1485 5.93 101.2485 7.6 ;
      RECT MASK 2 55.0085 6.021 55.0685 6.639 ;
      RECT MASK 2 10.9705 6.17 11.0305 6.891 ;
      RECT MASK 2 12.4905 6.17 12.5505 6.388 ;
      RECT MASK 2 14.8025 6.17 14.8625 6.388 ;
      RECT MASK 2 15.2605 6.17 15.3205 6.388 ;
      RECT MASK 2 15.7185 6.17 15.7785 6.388 ;
      RECT MASK 2 16.1765 6.17 16.2365 6.388 ;
      RECT MASK 2 16.6345 6.17 16.6945 6.388 ;
      RECT MASK 2 17.0925 6.17 17.1525 6.388 ;
      RECT MASK 2 17.5505 6.17 17.6105 6.388 ;
      RECT MASK 2 18.0085 6.17 18.0685 6.388 ;
      RECT MASK 2 18.4665 6.17 18.5265 6.388 ;
      RECT MASK 2 18.9245 6.17 18.9845 6.388 ;
      RECT MASK 2 19.3825 6.17 19.4425 6.388 ;
      RECT MASK 2 19.8405 6.17 19.9005 6.388 ;
      RECT MASK 2 20.2985 6.17 20.3585 6.388 ;
      RECT MASK 2 20.7565 6.17 20.8165 6.388 ;
      RECT MASK 2 26.1205 6.17 26.1805 6.388 ;
      RECT MASK 2 26.5785 6.17 26.6385 6.388 ;
      RECT MASK 2 27.0365 6.17 27.0965 6.388 ;
      RECT MASK 2 27.4945 6.17 27.5545 6.388 ;
      RECT MASK 2 27.9525 6.17 28.0125 6.388 ;
      RECT MASK 2 28.4105 6.17 28.4705 6.388 ;
      RECT MASK 2 28.8685 6.17 28.9285 6.388 ;
      RECT MASK 2 29.3265 6.17 29.3865 6.388 ;
      RECT MASK 2 29.7845 6.17 29.8445 6.388 ;
      RECT MASK 2 30.2425 6.17 30.3025 6.388 ;
      RECT MASK 2 30.7005 6.17 30.7605 6.388 ;
      RECT MASK 2 31.1585 6.17 31.2185 6.388 ;
      RECT MASK 2 31.6165 6.17 31.6765 6.388 ;
      RECT MASK 2 32.0745 6.17 32.1345 6.388 ;
      RECT MASK 2 34.3865 6.17 34.4465 6.388 ;
      RECT MASK 2 35.9065 6.17 35.9665 6.891 ;
      RECT MASK 2 21.2145 6.175 21.2745 6.388 ;
      RECT MASK 2 25.6625 6.175 25.7225 6.388 ;
      RECT MASK 2 53.245 6.205 53.305 8.585 ;
      RECT MASK 2 11.5745 6.208 11.6345 6.485 ;
      RECT MASK 2 35.3025 6.208 35.3625 6.485 ;
      RECT MASK 2 22.4385 6.29 22.4985 7.255 ;
      RECT MASK 2 23.0385 6.29 23.0985 7.255 ;
      RECT MASK 2 23.8385 6.29 23.8985 7.255 ;
      RECT MASK 2 24.4385 6.29 24.4985 7.255 ;
      RECT MASK 2 48.8745 6.3725 48.9345 7.4875 ;
      RECT MASK 2 52.913 6.397 52.973 10.253 ;
      RECT MASK 2 53.9295 6.4925 53.9895 7.449 ;
      RECT MASK 2 56.0875 6.4925 56.1475 7.405 ;
      RECT MASK 2 62.429 6.5 62.489 6.962 ;
      RECT MASK 2 61.513 6.505 61.573 6.962 ;
      RECT MASK 2 3.4235 6.508 3.4835 6.992 ;
      RECT MASK 2 10.1025 6.508 10.1625 6.725 ;
      RECT MASK 2 36.7745 6.508 36.8345 6.725 ;
      RECT MASK 2 43.4535 6.508 43.5135 6.992 ;
      RECT MASK 2 5.5145 6.53 5.5745 6.891 ;
      RECT MASK 2 5.7305 6.53 5.7905 6.891 ;
      RECT MASK 2 6.4215 6.53 6.4815 6.891 ;
      RECT MASK 2 6.6335 6.53 6.6935 6.891 ;
      RECT MASK 2 7.3375 6.53 7.3975 6.891 ;
      RECT MASK 2 7.5495 6.53 7.6095 6.891 ;
      RECT MASK 2 8.2495 6.53 8.3095 6.891 ;
      RECT MASK 2 8.4615 6.53 8.5215 6.891 ;
      RECT MASK 2 38.4155 6.53 38.4755 6.891 ;
      RECT MASK 2 38.6275 6.53 38.6875 6.891 ;
      RECT MASK 2 39.3275 6.53 39.3875 6.891 ;
      RECT MASK 2 39.5395 6.53 39.5995 6.891 ;
      RECT MASK 2 40.2435 6.53 40.3035 6.891 ;
      RECT MASK 2 40.4555 6.53 40.5155 6.891 ;
      RECT MASK 2 41.1465 6.53 41.2065 6.891 ;
      RECT MASK 2 41.3625 6.53 41.4225 6.891 ;
      RECT MASK 2 17.894 6.55 17.954 6.73 ;
      RECT MASK 2 19.268 6.55 19.328 6.73 ;
      RECT MASK 2 20.184 6.55 20.244 6.73 ;
      RECT MASK 2 26.693 6.55 26.753 6.73 ;
      RECT MASK 2 27.609 6.55 27.669 6.73 ;
      RECT MASK 2 28.983 6.55 29.043 6.73 ;
      RECT MASK 2 2.6325 6.609 2.6925 6.891 ;
      RECT MASK 2 44.2445 6.609 44.3045 6.891 ;
      RECT MASK 2 61.971 6.62 62.031 6.962 ;
      RECT MASK 2 62.887 6.62 62.947 6.962 ;
      RECT MASK 2 61.055 6.625 61.115 6.962 ;
      RECT MASK 2 48.1275 6.639 48.1875 7.221 ;
      RECT MASK 2 57.849 6.6425 57.909 7.7575 ;
      RECT MASK 2 22.6385 6.725 22.6985 6.865 ;
      RECT MASK 2 24.2385 6.725 24.2985 6.865 ;
      RECT MASK 2 55.0085 6.759 55.0685 7.405 ;
      RECT MASK 2 55.6725 6.759 55.7325 7.405 ;
      RECT MASK 2 17.207 6.77 17.267 6.95 ;
      RECT MASK 2 18.581 6.77 18.641 6.95 ;
      RECT MASK 2 28.296 6.77 28.356 6.95 ;
      RECT MASK 2 29.67 6.77 29.73 6.95 ;
      RECT MASK 2 46.9655 6.814 47.0255 7.046 ;
      RECT MASK 2 47.2975 6.814 47.3575 7.046 ;
      RECT MASK 2 47.6295 6.814 47.6895 7.046 ;
      RECT MASK 2 22.2385 6.874 22.2985 7.62 ;
      RECT MASK 2 22.8385 6.874 22.8985 7.62 ;
      RECT MASK 2 23.2385 6.874 23.2985 7.62 ;
      RECT MASK 2 23.6385 6.874 23.6985 7.62 ;
      RECT MASK 2 24.0385 6.874 24.0985 7.62 ;
      RECT MASK 2 24.6385 6.874 24.6985 7.62 ;
      RECT MASK 2 12.9915 6.912 13.0515 7.325 ;
      RECT MASK 2 33.8855 6.912 33.9455 7.325 ;
      RECT MASK 2 1.7055 6.9125 1.7655 7.885 ;
      RECT MASK 2 45.1715 6.9125 45.2315 7.885 ;
      RECT MASK 2 91.5785 6.9305 91.6785 8.46 ;
      RECT MASK 2 95.0265 6.9305 95.1265 8.46 ;
      RECT MASK 2 54.5105 6.934 54.5705 7.405 ;
      RECT MASK 2 83.7925 6.96 83.8925 8.46 ;
      RECT MASK 2 84.1285 6.96 84.2285 8.46 ;
      RECT MASK 2 86.7845 6.96 86.8845 8.46 ;
      RECT MASK 2 87.7805 6.96 87.8805 8.46 ;
      RECT MASK 2 88.1125 6.96 88.2125 8.46 ;
      RECT MASK 2 98.4925 6.96 98.5925 8.46 ;
      RECT MASK 2 98.8245 6.96 98.9245 8.46 ;
      RECT MASK 2 99.8205 6.96 99.9205 8.46 ;
      RECT MASK 2 102.4765 6.96 102.5765 8.46 ;
      RECT MASK 2 102.8125 6.96 102.9125 8.46 ;
      RECT MASK 2 88.4445 6.965 88.5045 8.46 ;
      RECT MASK 2 89.1345 6.965 89.1945 8.46 ;
      RECT MASK 2 89.7005 6.965 89.7605 8.46 ;
      RECT MASK 2 89.9565 6.965 90.0165 8.46 ;
      RECT MASK 2 90.4545 6.965 90.5145 8.46 ;
      RECT MASK 2 91.2165 6.965 91.2765 8.46 ;
      RECT MASK 2 95.4285 6.965 95.4885 8.46 ;
      RECT MASK 2 96.1905 6.965 96.2505 8.46 ;
      RECT MASK 2 96.6885 6.965 96.7485 8.46 ;
      RECT MASK 2 96.9445 6.965 97.0045 8.46 ;
      RECT MASK 2 97.5105 6.965 97.5705 8.46 ;
      RECT MASK 2 98.2005 6.965 98.2605 8.46 ;
      RECT MASK 2 10.4185 6.9725 10.4785 7.89 ;
      RECT MASK 2 13.6465 6.9725 13.7065 7.89 ;
      RECT MASK 2 33.2305 6.9725 33.2905 7.89 ;
      RECT MASK 2 36.4585 6.9725 36.5185 7.89 ;
      RECT MASK 2 22.6385 7.021 22.6985 7.62 ;
      RECT MASK 2 24.2385 7.021 24.2985 7.62 ;
      RECT MASK 2 2.6325 7.112 2.6925 7.89 ;
      RECT MASK 2 11.5745 7.112 11.6345 7.33 ;
      RECT MASK 2 12.4905 7.112 12.5505 7.325 ;
      RECT MASK 2 14.8025 7.112 14.8625 7.33 ;
      RECT MASK 2 15.2605 7.112 15.3205 7.33 ;
      RECT MASK 2 15.7185 7.112 15.7785 7.33 ;
      RECT MASK 2 16.1765 7.112 16.2365 7.33 ;
      RECT MASK 2 16.6345 7.112 16.6945 7.33 ;
      RECT MASK 2 17.0925 7.112 17.1525 7.33 ;
      RECT MASK 2 17.5505 7.112 17.6105 7.33 ;
      RECT MASK 2 18.0085 7.112 18.0685 7.33 ;
      RECT MASK 2 18.4665 7.112 18.5265 7.33 ;
      RECT MASK 2 18.9245 7.112 18.9845 7.33 ;
      RECT MASK 2 19.3825 7.112 19.4425 7.33 ;
      RECT MASK 2 19.8405 7.112 19.9005 7.33 ;
      RECT MASK 2 20.2985 7.112 20.3585 7.33 ;
      RECT MASK 2 20.7565 7.112 20.8165 7.33 ;
      RECT MASK 2 21.2145 7.112 21.2745 7.325 ;
      RECT MASK 2 25.6625 7.112 25.7225 7.325 ;
      RECT MASK 2 26.1205 7.112 26.1805 7.33 ;
      RECT MASK 2 26.5785 7.112 26.6385 7.33 ;
      RECT MASK 2 27.0365 7.112 27.0965 7.33 ;
      RECT MASK 2 27.4945 7.112 27.5545 7.33 ;
      RECT MASK 2 27.9525 7.112 28.0125 7.33 ;
      RECT MASK 2 28.4105 7.112 28.4705 7.33 ;
      RECT MASK 2 28.8685 7.112 28.9285 7.33 ;
      RECT MASK 2 29.3265 7.112 29.3865 7.33 ;
      RECT MASK 2 29.7845 7.112 29.8445 7.33 ;
      RECT MASK 2 30.2425 7.112 30.3025 7.33 ;
      RECT MASK 2 30.7005 7.112 30.7605 7.33 ;
      RECT MASK 2 31.1585 7.112 31.2185 7.33 ;
      RECT MASK 2 31.6165 7.112 31.6765 7.33 ;
      RECT MASK 2 32.0745 7.112 32.1345 7.33 ;
      RECT MASK 2 34.3865 7.112 34.4465 7.325 ;
      RECT MASK 2 35.3025 7.112 35.3625 7.33 ;
      RECT MASK 2 44.2445 7.112 44.3045 7.89 ;
      RECT MASK 2 54.1825 7.2335 54.2425 9.587 ;
      RECT MASK 2 46.9655 7.238 47.0255 8.062 ;
      RECT MASK 2 47.2975 7.238 47.3575 8.062 ;
      RECT MASK 2 47.6295 7.238 47.6895 8.062 ;
      RECT MASK 2 84.7925 7.315 84.8925 7.721 ;
      RECT MASK 2 85.1245 7.315 85.2245 7.721 ;
      RECT MASK 2 85.7885 7.315 85.8885 7.721 ;
      RECT MASK 2 86.4525 7.315 86.5525 7.721 ;
      RECT MASK 2 100.1525 7.315 100.2525 7.721 ;
      RECT MASK 2 100.8165 7.315 100.9165 7.721 ;
      RECT MASK 2 101.4805 7.315 101.5805 7.721 ;
      RECT MASK 2 101.8125 7.315 101.9125 7.721 ;
      RECT MASK 2 48.1275 7.341 48.1875 7.959 ;
      RECT MASK 2 2.2785 7.374 2.3385 7.89 ;
      RECT MASK 2 44.5985 7.374 44.6585 7.89 ;
      RECT MASK 2 50.2985 7.385 50.3385 7.61 ;
      RECT MASK 2 50.9625 7.385 51.0025 7.61 ;
      RECT MASK 2 51.6265 7.385 51.6665 7.61 ;
      RECT MASK 2 52.2905 7.385 52.3305 7.61 ;
      RECT MASK 2 59.452 7.4 59.512 8.555 ;
      RECT MASK 2 64.032 7.4 64.092 8.555 ;
      RECT MASK 2 64.49 7.4 64.55 8.555 ;
      RECT MASK 2 58.994 7.405 59.054 8.555 ;
      RECT MASK 2 64.948 7.405 65.008 8.555 ;
      RECT MASK 2 22.4385 7.41 22.4985 7.62 ;
      RECT MASK 2 23.0385 7.41 23.0985 7.62 ;
      RECT MASK 2 23.8385 7.41 23.8985 7.62 ;
      RECT MASK 2 24.4385 7.41 24.4985 7.62 ;
      RECT MASK 2 61.055 7.438 61.115 7.775 ;
      RECT MASK 2 61.513 7.438 61.573 7.895 ;
      RECT MASK 2 61.971 7.438 62.031 7.78 ;
      RECT MASK 2 62.429 7.438 62.489 7.9 ;
      RECT MASK 2 62.887 7.438 62.947 7.78 ;
      RECT MASK 2 87.4485 7.5595 87.5485 7.891 ;
      RECT MASK 2 99.1565 7.5595 99.2565 7.891 ;
      RECT MASK 2 49.5105 7.6475 49.5705 8.8845 ;
      RECT MASK 2 50.2985 7.865 50.3385 8.09 ;
      RECT MASK 2 50.9625 7.865 51.0025 8.09 ;
      RECT MASK 2 51.6265 7.865 51.6665 8.09 ;
      RECT MASK 2 52.2905 7.865 52.3305 8.09 ;
      RECT MASK 2 49.1785 7.8665 49.2385 9.1765 ;
      RECT MASK 2 62.429 8.06 62.489 8.522 ;
      RECT MASK 2 61.513 8.065 61.573 8.522 ;
      RECT MASK 2 2.2785 8.07 2.3385 8.586 ;
      RECT MASK 2 2.6325 8.07 2.6925 8.848 ;
      RECT MASK 2 10.4185 8.07 10.4785 8.9875 ;
      RECT MASK 2 11.2205 8.07 11.2805 10.35 ;
      RECT MASK 2 12.0325 8.07 12.0925 10.35 ;
      RECT MASK 2 12.8445 8.07 12.9045 10.35 ;
      RECT MASK 2 13.6465 8.07 13.7065 8.9875 ;
      RECT MASK 2 1.7055 8.075 1.7655 9.0475 ;
      RECT MASK 2 48.1275 8.079 48.1875 8.486 ;
      RECT MASK 2 48.4595 8.079 48.5195 8.661 ;
      RECT MASK 2 61.971 8.18 62.031 8.522 ;
      RECT MASK 2 62.887 8.18 62.947 8.522 ;
      RECT MASK 2 61.055 8.185 61.115 8.522 ;
      RECT MASK 2 57.849 8.2025 57.909 9.3175 ;
      RECT MASK 2 46.9655 8.254 47.0255 8.486 ;
      RECT MASK 2 47.2975 8.254 47.3575 8.486 ;
      RECT MASK 2 65.864 8.3225 65.924 9.378 ;
      RECT MASK 2 22.2385 8.34 22.2985 9.086 ;
      RECT MASK 2 22.4385 8.34 22.4985 8.55 ;
      RECT MASK 2 22.6385 8.34 22.6985 8.939 ;
      RECT MASK 2 22.8385 8.34 22.8985 9.086 ;
      RECT MASK 2 23.0385 8.34 23.0985 8.55 ;
      RECT MASK 2 23.2385 8.34 23.2985 9.086 ;
      RECT MASK 2 50.2985 8.465 50.3385 10.015 ;
      RECT MASK 2 50.9625 8.465 51.0025 10.015 ;
      RECT MASK 2 51.6265 8.465 51.6665 10.015 ;
      RECT MASK 2 52.2905 8.465 52.3305 10.015 ;
      RECT MASK 2 47.7955 8.47 47.8555 8.661 ;
      RECT MASK 2 68.117 8.495 68.177 8.966 ;
      RECT MASK 2 70.178 8.495 70.238 8.966 ;
      RECT MASK 2 32.246 8.501 32.306 9.171 ;
      RECT MASK 2 32.9395 8.501 32.9995 9.171 ;
      RECT MASK 2 33.162 8.501 33.222 9.171 ;
      RECT MASK 2 33.8555 8.501 33.9155 9.171 ;
      RECT MASK 2 34.078 8.501 34.138 9.171 ;
      RECT MASK 2 34.7715 8.501 34.8315 9.171 ;
      RECT MASK 2 34.994 8.501 35.054 9.171 ;
      RECT MASK 2 35.6875 8.501 35.7475 9.171 ;
      RECT MASK 2 35.91 8.501 35.97 9.171 ;
      RECT MASK 2 36.6035 8.501 36.6635 9.171 ;
      RECT MASK 2 36.826 8.501 36.886 9.171 ;
      RECT MASK 2 37.5195 8.501 37.5795 9.171 ;
      RECT MASK 2 37.742 8.501 37.802 9.171 ;
      RECT MASK 2 38.4355 8.501 38.4955 9.171 ;
      RECT MASK 2 11.5745 8.63 11.6345 8.848 ;
      RECT MASK 2 14.8025 8.63 14.8625 8.848 ;
      RECT MASK 2 15.2605 8.63 15.3205 8.848 ;
      RECT MASK 2 15.7185 8.63 15.7785 8.848 ;
      RECT MASK 2 16.1765 8.63 16.2365 8.848 ;
      RECT MASK 2 16.6345 8.63 16.6945 8.848 ;
      RECT MASK 2 17.0925 8.63 17.1525 8.848 ;
      RECT MASK 2 17.5505 8.63 17.6105 8.848 ;
      RECT MASK 2 18.0085 8.63 18.0685 8.848 ;
      RECT MASK 2 18.4665 8.63 18.5265 8.848 ;
      RECT MASK 2 18.9245 8.63 18.9845 8.848 ;
      RECT MASK 2 19.3825 8.63 19.4425 8.848 ;
      RECT MASK 2 19.8405 8.63 19.9005 8.848 ;
      RECT MASK 2 20.2985 8.63 20.3585 8.848 ;
      RECT MASK 2 20.7565 8.63 20.8165 8.848 ;
      RECT MASK 2 12.4905 8.635 12.5505 8.848 ;
      RECT MASK 2 12.9915 8.635 13.0515 9.048 ;
      RECT MASK 2 21.2145 8.635 21.2745 8.848 ;
      RECT MASK 2 61.284 8.675 61.344 9.9175 ;
      RECT MASK 2 46.9655 8.678 47.0255 9.502 ;
      RECT MASK 2 47.2975 8.678 47.3575 9.502 ;
      RECT MASK 2 48.1275 8.678 48.1875 9.502 ;
      RECT MASK 2 62.658 8.678 62.718 9.178 ;
      RECT MASK 2 63.116 8.678 63.176 9.178 ;
      RECT MASK 2 63.574 8.678 63.634 9.178 ;
      RECT MASK 2 64.032 8.678 64.092 9.178 ;
      RECT MASK 2 64.49 8.678 64.55 9.178 ;
      RECT MASK 2 64.948 8.678 65.008 9.178 ;
      RECT MASK 2 65.406 8.678 65.466 9.178 ;
      RECT MASK 2 22.4385 8.705 22.4985 9.67 ;
      RECT MASK 2 23.0385 8.705 23.0985 9.67 ;
      RECT MASK 2 47.7955 8.781 47.8555 9.399 ;
      RECT MASK 2 58.765 8.965 58.825 9.178 ;
      RECT MASK 2 59.223 8.965 59.283 9.178 ;
      RECT MASK 2 59.681 8.965 59.741 9.178 ;
      RECT MASK 2 60.139 8.965 60.199 9.178 ;
      RECT MASK 2 3.4235 8.968 3.4835 9.452 ;
      RECT MASK 2 32.488 8.98 32.548 9.171 ;
      RECT MASK 2 33.404 8.98 33.464 9.171 ;
      RECT MASK 2 34.32 8.98 34.38 9.171 ;
      RECT MASK 2 35.236 8.98 35.296 9.171 ;
      RECT MASK 2 36.152 8.98 36.212 9.171 ;
      RECT MASK 2 37.068 8.98 37.128 9.171 ;
      RECT MASK 2 37.984 8.98 38.044 9.171 ;
      RECT MASK 2 17.207 9.01 17.267 9.19 ;
      RECT MASK 2 18.581 9.01 18.641 9.19 ;
      RECT MASK 2 2.6325 9.069 2.6925 9.351 ;
      RECT MASK 2 5.5145 9.069 5.5745 9.43 ;
      RECT MASK 2 5.7305 9.069 5.7905 9.43 ;
      RECT MASK 2 6.4215 9.069 6.4815 9.43 ;
      RECT MASK 2 6.6335 9.069 6.6935 9.43 ;
      RECT MASK 2 7.3375 9.069 7.3975 9.43 ;
      RECT MASK 2 7.5495 9.069 7.6095 9.43 ;
      RECT MASK 2 8.2495 9.069 8.3095 9.43 ;
      RECT MASK 2 8.4615 9.069 8.5215 9.43 ;
      RECT MASK 2 10.9705 9.069 11.0305 9.79 ;
      RECT MASK 2 22.6385 9.095 22.6985 9.235 ;
      RECT MASK 2 80.1445 9.202 80.4645 9.926 ;
      RECT MASK 2 106.2405 9.202 106.5605 9.926 ;
      RECT MASK 2 17.894 9.23 17.954 9.41 ;
      RECT MASK 2 19.268 9.23 19.328 9.41 ;
      RECT MASK 2 20.184 9.23 20.244 9.41 ;
      RECT MASK 2 42.9555 9.231 43.0155 11.037 ;
      RECT MASK 2 10.1025 9.235 10.1625 9.452 ;
      RECT MASK 2 48.8745 9.2525 48.9345 10.165 ;
      RECT MASK 2 32.596 9.291 32.656 9.909 ;
      RECT MASK 2 33.512 9.291 33.572 9.909 ;
      RECT MASK 2 34.428 9.291 34.488 9.909 ;
      RECT MASK 2 35.344 9.291 35.404 9.909 ;
      RECT MASK 2 36.26 9.291 36.32 9.909 ;
      RECT MASK 2 37.176 9.291 37.236 9.909 ;
      RECT MASK 2 38.092 9.291 38.152 9.909 ;
      RECT MASK 2 62.658 9.298 62.718 9.782 ;
      RECT MASK 2 22.2385 9.319 22.2985 10.08 ;
      RECT MASK 2 22.8385 9.319 22.8985 10.065 ;
      RECT MASK 2 23.2385 9.319 23.2985 10.08 ;
      RECT MASK 2 65.406 9.325 65.466 9.681 ;
      RECT MASK 2 43.2975 9.327 43.3575 10.253 ;
      RECT MASK 2 1.7055 9.3725 1.7655 10.345 ;
      RECT MASK 2 59.3375 9.399 59.3975 9.6925 ;
      RECT MASK 2 64.719 9.399 64.779 9.64 ;
      RECT MASK 2 68.454 9.417 68.514 9.723 ;
      RECT MASK 2 68.696 9.417 68.756 9.723 ;
      RECT MASK 2 68.912 9.417 68.972 9.723 ;
      RECT MASK 2 69.154 9.417 69.214 9.723 ;
      RECT MASK 2 69.599 9.417 69.659 9.723 ;
      RECT MASK 2 69.841 9.417 69.901 9.723 ;
      RECT MASK 2 10.4185 9.4325 10.4785 10.35 ;
      RECT MASK 2 13.6465 9.4325 13.7065 10.35 ;
      RECT MASK 2 64.032 9.445 64.092 10.082 ;
      RECT MASK 2 54.5865 9.447 54.6465 9.753 ;
      RECT MASK 2 54.8285 9.447 54.8885 9.753 ;
      RECT MASK 2 55.0445 9.447 55.1045 9.753 ;
      RECT MASK 2 55.2865 9.447 55.3465 9.753 ;
      RECT MASK 2 22.6385 9.466 22.6985 10.065 ;
      RECT MASK 2 11.5745 9.475 11.6345 9.752 ;
      RECT MASK 2 47.7955 9.519 47.8555 10.165 ;
      RECT MASK 2 48.4595 9.519 48.5195 10.165 ;
      RECT MASK 2 57.266 9.5615 57.326 10.353 ;
      RECT MASK 2 64.948 9.565 65.008 10.082 ;
      RECT MASK 2 2.6325 9.572 2.6925 10.35 ;
      RECT MASK 2 12.4905 9.572 12.5505 9.79 ;
      RECT MASK 2 14.8025 9.572 14.8625 9.79 ;
      RECT MASK 2 15.2605 9.572 15.3205 9.79 ;
      RECT MASK 2 15.7185 9.572 15.7785 9.79 ;
      RECT MASK 2 16.1765 9.572 16.2365 9.79 ;
      RECT MASK 2 16.6345 9.572 16.6945 9.79 ;
      RECT MASK 2 17.0925 9.572 17.1525 9.79 ;
      RECT MASK 2 17.5505 9.572 17.6105 9.79 ;
      RECT MASK 2 18.0085 9.572 18.0685 9.79 ;
      RECT MASK 2 18.4665 9.572 18.5265 9.79 ;
      RECT MASK 2 18.9245 9.572 18.9845 9.79 ;
      RECT MASK 2 19.3825 9.572 19.4425 9.79 ;
      RECT MASK 2 19.8405 9.572 19.9005 9.79 ;
      RECT MASK 2 20.2985 9.572 20.3585 9.79 ;
      RECT MASK 2 20.7565 9.572 20.8165 9.79 ;
      RECT MASK 2 21.2145 9.572 21.2745 9.785 ;
      RECT MASK 2 58.765 9.601 58.825 10.68 ;
      RECT MASK 2 60.139 9.601 60.199 10.68 ;
      RECT MASK 2 46.9655 9.694 47.0255 10.165 ;
      RECT MASK 2 47.2975 9.694 47.3575 10.165 ;
      RECT MASK 2 67.659 9.7325 67.719 10.645 ;
      RECT MASK 2 70.636 9.7325 70.696 10.645 ;
      RECT MASK 2 31.5655 9.7625 31.6255 10.218 ;
      RECT MASK 2 39.1225 9.7625 39.1825 10.218 ;
      RECT MASK 2 53.7915 9.7625 53.8515 10.675 ;
      RECT MASK 2 56.0815 9.7625 56.1415 10.675 ;
      RECT MASK 2 57.849 9.7625 57.909 10.68 ;
      RECT MASK 2 2.2785 9.834 2.3385 10.35 ;
      RECT MASK 2 22.4385 9.855 22.4985 10.065 ;
      RECT MASK 2 23.0385 9.855 23.0985 10.065 ;
      RECT MASK 2 66.7185 9.876 66.7785 10.545 ;
      RECT MASK 2 59.223 9.902 59.283 10.12 ;
      RECT MASK 2 59.681 9.902 59.741 10.12 ;
      RECT MASK 2 62.658 9.902 62.718 10.68 ;
      RECT MASK 2 63.116 9.902 63.176 10.68 ;
      RECT MASK 2 63.574 9.902 63.634 10.68 ;
      RECT MASK 2 64.49 9.902 64.55 10.68 ;
      RECT MASK 2 65.406 9.902 65.466 10.68 ;
      RECT MASK 2 65.864 9.902 65.924 10.68 ;
      RECT MASK 2 32.246 10.029 32.306 10.699 ;
      RECT MASK 2 32.9395 10.029 32.9995 10.699 ;
      RECT MASK 2 33.162 10.029 33.222 10.699 ;
      RECT MASK 2 33.8555 10.029 33.9155 10.699 ;
      RECT MASK 2 34.078 10.029 34.138 10.699 ;
      RECT MASK 2 34.7715 10.029 34.8315 10.699 ;
      RECT MASK 2 34.994 10.029 35.054 10.699 ;
      RECT MASK 2 35.6875 10.029 35.7475 10.699 ;
      RECT MASK 2 35.91 10.029 35.97 10.699 ;
      RECT MASK 2 36.6035 10.029 36.6635 10.699 ;
      RECT MASK 2 36.826 10.029 36.886 10.699 ;
      RECT MASK 2 37.5195 10.029 37.5795 10.699 ;
      RECT MASK 2 37.742 10.029 37.802 10.699 ;
      RECT MASK 2 38.4355 10.029 38.4955 10.699 ;
      RECT MASK 2 68.117 10.174 68.177 10.645 ;
      RECT MASK 2 58.307 10.445 58.367 10.675 ;
      RECT MASK 2 62.2 10.445 62.26 10.675 ;
      RECT MASK 2 39.6455 11.639 39.7055 12.731 ;
      RECT MASK 2 4.377 11.76 4.457 12.7 ;
      RECT MASK 2 8.527 11.76 8.607 12.416 ;
      RECT MASK 2 8.776 11.76 8.856 12.241 ;
      RECT MASK 2 9.108 11.76 9.188 12.241 ;
      RECT MASK 2 9.357 11.76 9.437 12.416 ;
      RECT MASK 2 10.187 11.76 10.267 12.416 ;
      RECT MASK 2 10.436 11.76 10.516 12.241 ;
      RECT MASK 2 10.768 11.76 10.848 12.241 ;
      RECT MASK 2 11.017 11.76 11.097 12.416 ;
      RECT MASK 2 22.637 11.76 22.717 12.416 ;
      RECT MASK 2 23.467 11.76 23.547 12.416 ;
      RECT MASK 2 24.297 11.76 24.377 12.416 ;
      RECT MASK 2 25.127 11.76 25.207 12.416 ;
      RECT MASK 2 25.957 11.76 26.037 12.416 ;
      RECT MASK 2 26.787 11.76 26.867 12.416 ;
      RECT MASK 2 28.447 11.76 28.527 12.416 ;
      RECT MASK 2 29.277 11.76 29.357 12.416 ;
      RECT MASK 2 30.937 11.76 31.017 12.416 ;
      RECT MASK 2 31.767 11.76 31.847 12.416 ;
      RECT MASK 2 32.597 11.76 32.677 12.416 ;
      RECT MASK 2 33.427 11.76 33.507 12.416 ;
      RECT MASK 2 34.257 11.76 34.337 12.416 ;
      RECT MASK 2 35.087 11.76 35.167 12.416 ;
      RECT MASK 2 35.917 11.76 35.997 12.416 ;
      RECT MASK 2 36.747 11.76 36.827 12.416 ;
      RECT MASK 2 37.577 11.76 37.657 12.416 ;
      RECT MASK 2 38.407 11.76 38.487 12.416 ;
      RECT MASK 2 39.237 11.76 39.317 12.416 ;
      RECT MASK 2 40.067 11.76 40.147 12.416 ;
      RECT MASK 2 42.557 11.76 42.637 12.416 ;
      RECT MASK 2 43.387 11.76 43.467 12.416 ;
      RECT MASK 2 44.217 11.76 44.297 12.416 ;
      RECT MASK 2 45.047 11.76 45.127 12.416 ;
      RECT MASK 2 45.462 11.76 45.542 12.552 ;
      RECT MASK 2 45.877 11.76 45.957 12.416 ;
      RECT MASK 2 46.292 11.76 46.372 12.5595 ;
      RECT MASK 2 46.707 11.76 46.787 12.416 ;
      RECT MASK 2 47.537 11.76 47.617 12.416 ;
      RECT MASK 2 48.367 11.76 48.447 12.416 ;
      RECT MASK 2 49.197 11.76 49.277 12.416 ;
      RECT MASK 2 50.027 11.76 50.107 12.416 ;
      RECT MASK 2 50.857 11.76 50.937 12.416 ;
      RECT MASK 2 51.687 11.76 51.767 12.416 ;
      RECT MASK 2 52.517 11.76 52.597 12.416 ;
      RECT MASK 2 53.347 11.76 53.427 12.416 ;
      RECT MASK 2 54.177 11.76 54.257 12.416 ;
      RECT MASK 2 55.007 11.76 55.087 12.416 ;
      RECT MASK 2 56.823 11.76 56.923 12.416 ;
      RECT MASK 2 57.653 11.76 57.753 12.416 ;
      RECT MASK 2 58.483 11.76 58.583 12.416 ;
      RECT MASK 2 59.313 11.76 59.413 12.416 ;
      RECT MASK 2 60.973 11.76 61.073 12.416 ;
      RECT MASK 2 61.803 11.76 61.903 12.416 ;
      RECT MASK 2 63.473 11.76 63.553 12.416 ;
      RECT MASK 2 64.303 11.76 64.383 12.416 ;
      RECT MASK 2 65.133 11.76 65.213 12.416 ;
      RECT MASK 2 65.963 11.76 66.043 12.416 ;
      RECT MASK 2 66.793 11.76 66.873 12.416 ;
      RECT MASK 2 67.623 11.76 67.703 12.416 ;
      RECT MASK 2 68.443 11.76 68.543 12.416 ;
      RECT MASK 2 69.273 11.76 69.373 12.416 ;
      RECT MASK 2 70.113 11.76 70.193 12.416 ;
      RECT MASK 2 70.943 11.76 71.023 12.416 ;
      RECT MASK 2 71.773 11.76 71.853 12.416 ;
      RECT MASK 2 72.603 11.76 72.683 12.416 ;
      RECT MASK 2 77.583 11.76 77.663 12.416 ;
      RECT MASK 2 78.413 11.76 78.493 12.416 ;
      RECT MASK 2 79.243 11.76 79.323 12.416 ;
      RECT MASK 2 80.073 11.76 80.153 12.416 ;
      RECT MASK 2 83.393 11.76 83.473 12.416 ;
      RECT MASK 2 84.223 11.76 84.303 12.416 ;
      RECT MASK 2 89.203 11.76 89.283 12.416 ;
      RECT MASK 2 90.033 11.76 90.113 12.416 ;
      RECT MASK 2 90.863 11.76 90.943 12.416 ;
      RECT MASK 2 91.693 11.76 91.773 12.416 ;
      RECT MASK 2 101.653 11.76 101.733 12.416 ;
      RECT MASK 2 102.483 11.76 102.563 12.416 ;
      RECT MASK 2 103.313 11.76 103.393 12.416 ;
      RECT MASK 2 104.143 11.76 104.223 12.416 ;
      RECT MASK 2 111.613 11.76 111.693 12.683 ;
      RECT MASK 2 73.36 12.38 73.42 13.1425 ;
      RECT MASK 2 69.708 12.383 69.768 13.019 ;
      RECT MASK 2 68.048 12.4045 68.108 13.017 ;
      RECT MASK 2 8.786 12.428 8.846 13.252 ;
      RECT MASK 2 9.118 12.428 9.178 13.252 ;
      RECT MASK 2 10.446 12.428 10.506 13.252 ;
      RECT MASK 2 10.778 12.428 10.838 13.252 ;
      RECT MASK 2 22.398 12.428 22.458 13.252 ;
      RECT MASK 2 23.726 12.428 23.786 13.252 ;
      RECT MASK 2 24.058 12.428 24.118 13.252 ;
      RECT MASK 2 25.386 12.428 25.446 13.252 ;
      RECT MASK 2 25.718 12.428 25.778 13.264 ;
      RECT MASK 2 27.046 12.428 27.106 13.264 ;
      RECT MASK 2 27.544 12.428 27.604 13.252 ;
      RECT MASK 2 28.706 12.428 28.766 13.264 ;
      RECT MASK 2 29.038 12.428 29.098 13.264 ;
      RECT MASK 2 30.034 12.428 30.094 13.252 ;
      RECT MASK 2 30.698 12.428 30.758 13.264 ;
      RECT MASK 2 32.026 12.428 32.086 13.264 ;
      RECT MASK 2 32.358 12.428 32.418 13.264 ;
      RECT MASK 2 33.686 12.428 33.746 13.264 ;
      RECT MASK 2 34.516 12.428 34.576 13.252 ;
      RECT MASK 2 34.848 12.428 34.908 13.252 ;
      RECT MASK 2 35.678 12.428 35.738 13.252 ;
      RECT MASK 2 37.006 12.428 37.066 13.252 ;
      RECT MASK 2 37.338 12.428 37.398 13.264 ;
      RECT MASK 2 38.666 12.428 38.726 13.264 ;
      RECT MASK 2 38.998 12.428 39.058 13.264 ;
      RECT MASK 2 40.326 12.428 40.386 13.264 ;
      RECT MASK 2 40.824 12.428 40.884 13.252 ;
      RECT MASK 2 41.654 12.428 41.714 13.252 ;
      RECT MASK 2 42.318 12.428 42.378 13.264 ;
      RECT MASK 2 43.646 12.428 43.706 13.264 ;
      RECT MASK 2 43.978 12.428 44.038 13.252 ;
      RECT MASK 2 45.306 12.428 45.366 13.252 ;
      RECT MASK 2 46.136 12.428 46.196 13.252 ;
      RECT MASK 2 46.966 12.428 47.026 13.252 ;
      RECT MASK 2 47.298 12.428 47.358 13.264 ;
      RECT MASK 2 48.626 12.428 48.686 13.264 ;
      RECT MASK 2 48.958 12.428 49.018 13.252 ;
      RECT MASK 2 50.286 12.428 50.346 13.252 ;
      RECT MASK 2 50.618 12.428 50.678 13.252 ;
      RECT MASK 2 51.946 12.428 52.006 13.252 ;
      RECT MASK 2 52.278 12.428 52.338 13.252 ;
      RECT MASK 2 53.606 12.428 53.666 13.252 ;
      RECT MASK 2 53.938 12.428 53.998 13.264 ;
      RECT MASK 2 55.266 12.428 55.326 13.264 ;
      RECT MASK 2 55.598 12.428 55.658 13.252 ;
      RECT MASK 2 57.092 12.428 57.152 13.264 ;
      RECT MASK 2 57.424 12.428 57.484 13.264 ;
      RECT MASK 2 58.752 12.428 58.812 13.252 ;
      RECT MASK 2 59.084 12.428 59.144 13.252 ;
      RECT MASK 2 60.08 12.428 60.14 13.252 ;
      RECT MASK 2 60.744 12.428 60.804 13.252 ;
      RECT MASK 2 62.072 12.428 62.132 13.252 ;
      RECT MASK 2 62.57 12.428 62.63 13.252 ;
      RECT MASK 2 63.732 12.428 63.792 13.264 ;
      RECT MASK 2 64.064 12.428 64.124 13.264 ;
      RECT MASK 2 65.392 12.428 65.452 13.252 ;
      RECT MASK 2 65.724 12.428 65.784 13.252 ;
      RECT MASK 2 67.052 12.428 67.112 13.252 ;
      RECT MASK 2 67.384 12.428 67.444 13.252 ;
      RECT MASK 2 68.712 12.428 68.772 13.252 ;
      RECT MASK 2 69.044 12.428 69.104 13.252 ;
      RECT MASK 2 70.372 12.428 70.432 13.252 ;
      RECT MASK 2 70.704 12.428 70.764 13.252 ;
      RECT MASK 2 72.032 12.428 72.092 13.252 ;
      RECT MASK 2 72.364 12.428 72.424 13.252 ;
      RECT MASK 2 77.344 12.428 77.404 13.252 ;
      RECT MASK 2 78.672 12.428 78.732 13.252 ;
      RECT MASK 2 79.004 12.428 79.064 13.252 ;
      RECT MASK 2 80.332 12.428 80.392 13.252 ;
      RECT MASK 2 83.652 12.428 83.712 13.264 ;
      RECT MASK 2 83.984 12.428 84.044 13.264 ;
      RECT MASK 2 88.964 12.428 89.024 13.252 ;
      RECT MASK 2 90.292 12.428 90.352 13.252 ;
      RECT MASK 2 90.624 12.428 90.684 13.252 ;
      RECT MASK 2 91.952 12.428 92.012 13.252 ;
      RECT MASK 2 101.912 12.428 101.972 13.252 ;
      RECT MASK 2 102.244 12.428 102.304 13.252 ;
      RECT MASK 2 103.572 12.428 103.632 13.252 ;
      RECT MASK 2 103.904 12.428 103.964 13.252 ;
      RECT MASK 2 45.4725 13.043 45.5325 14.459 ;
      RECT MASK 2 5.217 13.264 5.277 14.336 ;
      RECT MASK 2 6.047 13.264 6.107 14.336 ;
      RECT MASK 2 6.877 13.264 6.937 14.336 ;
      RECT MASK 2 7.707 13.264 7.767 14.336 ;
      RECT MASK 2 8.537 13.264 8.597 14.336 ;
      RECT MASK 2 9.367 13.264 9.427 14.336 ;
      RECT MASK 2 10.197 13.264 10.257 14.336 ;
      RECT MASK 2 11.027 13.264 11.087 14.336 ;
      RECT MASK 2 11.857 13.264 11.917 14.336 ;
      RECT MASK 2 12.687 13.264 12.747 14.336 ;
      RECT MASK 2 13.517 13.264 13.577 14.336 ;
      RECT MASK 2 14.347 13.264 14.407 14.336 ;
      RECT MASK 2 15.177 13.264 15.237 14.336 ;
      RECT MASK 2 16.007 13.264 16.067 14.336 ;
      RECT MASK 2 16.837 13.264 16.897 14.336 ;
      RECT MASK 2 17.667 13.264 17.727 14.336 ;
      RECT MASK 2 18.497 13.264 18.557 14.336 ;
      RECT MASK 2 19.327 13.264 19.387 14.336 ;
      RECT MASK 2 20.157 13.264 20.217 14.336 ;
      RECT MASK 2 20.987 13.264 21.047 14.336 ;
      RECT MASK 2 21.817 13.264 21.877 14.336 ;
      RECT MASK 2 22.647 13.264 22.707 14.336 ;
      RECT MASK 2 23.477 13.264 23.537 14.336 ;
      RECT MASK 2 24.307 13.264 24.367 14.336 ;
      RECT MASK 2 25.137 13.264 25.197 14.336 ;
      RECT MASK 2 25.967 13.264 26.027 14.336 ;
      RECT MASK 2 26.797 13.264 26.857 14.336 ;
      RECT MASK 2 28.457 13.264 28.517 14.336 ;
      RECT MASK 2 29.287 13.264 29.347 14.336 ;
      RECT MASK 2 30.947 13.264 31.007 14.336 ;
      RECT MASK 2 31.777 13.264 31.837 14.336 ;
      RECT MASK 2 32.607 13.264 32.667 14.336 ;
      RECT MASK 2 33.437 13.264 33.497 14.336 ;
      RECT MASK 2 34.267 13.264 34.327 13.458 ;
      RECT MASK 2 35.097 13.264 35.157 13.458 ;
      RECT MASK 2 35.927 13.264 35.987 14.336 ;
      RECT MASK 2 36.757 13.264 36.817 14.336 ;
      RECT MASK 2 37.587 13.264 37.647 14.336 ;
      RECT MASK 2 38.417 13.264 38.477 14.336 ;
      RECT MASK 2 39.247 13.264 39.307 14.336 ;
      RECT MASK 2 40.077 13.264 40.137 14.336 ;
      RECT MASK 2 42.567 13.264 42.627 14.336 ;
      RECT MASK 2 43.397 13.264 43.457 14.336 ;
      RECT MASK 2 44.227 13.264 44.287 14.336 ;
      RECT MASK 2 45.057 13.264 45.117 14.336 ;
      RECT MASK 2 45.887 13.264 45.947 13.458 ;
      RECT MASK 2 46.717 13.264 46.777 14.336 ;
      RECT MASK 2 47.547 13.264 47.607 14.336 ;
      RECT MASK 2 48.377 13.264 48.437 14.336 ;
      RECT MASK 2 49.207 13.264 49.267 14.336 ;
      RECT MASK 2 50.037 13.264 50.097 14.336 ;
      RECT MASK 2 50.867 13.264 50.927 14.336 ;
      RECT MASK 2 51.697 13.264 51.757 14.336 ;
      RECT MASK 2 52.527 13.264 52.587 14.336 ;
      RECT MASK 2 53.357 13.264 53.417 14.336 ;
      RECT MASK 2 54.187 13.264 54.247 14.336 ;
      RECT MASK 2 55.017 13.264 55.077 14.336 ;
      RECT MASK 2 56.843 13.264 56.903 14.336 ;
      RECT MASK 2 57.673 13.264 57.733 14.336 ;
      RECT MASK 2 58.503 13.264 58.563 14.336 ;
      RECT MASK 2 59.333 13.264 59.393 14.336 ;
      RECT MASK 2 60.993 13.264 61.053 14.336 ;
      RECT MASK 2 61.823 13.264 61.883 14.336 ;
      RECT MASK 2 63.483 13.264 63.543 14.336 ;
      RECT MASK 2 64.313 13.264 64.373 14.336 ;
      RECT MASK 2 65.143 13.264 65.203 14.336 ;
      RECT MASK 2 65.973 13.264 66.033 14.336 ;
      RECT MASK 2 66.803 13.264 66.863 14.336 ;
      RECT MASK 2 67.633 13.264 67.693 14.336 ;
      RECT MASK 2 68.463 13.264 68.523 14.336 ;
      RECT MASK 2 69.293 13.264 69.353 14.336 ;
      RECT MASK 2 70.123 13.264 70.183 14.336 ;
      RECT MASK 2 70.953 13.264 71.013 14.336 ;
      RECT MASK 2 71.783 13.264 71.843 14.336 ;
      RECT MASK 2 72.613 13.264 72.673 14.336 ;
      RECT MASK 2 73.443 13.264 73.503 14.336 ;
      RECT MASK 2 74.273 13.264 74.333 14.336 ;
      RECT MASK 2 75.103 13.264 75.163 14.336 ;
      RECT MASK 2 75.933 13.264 75.993 14.336 ;
      RECT MASK 2 76.763 13.264 76.823 14.336 ;
      RECT MASK 2 77.593 13.264 77.653 14.336 ;
      RECT MASK 2 78.423 13.264 78.483 14.336 ;
      RECT MASK 2 79.253 13.264 79.313 14.336 ;
      RECT MASK 2 80.083 13.264 80.143 14.336 ;
      RECT MASK 2 80.913 13.264 80.973 14.336 ;
      RECT MASK 2 81.743 13.264 81.803 14.336 ;
      RECT MASK 2 82.573 13.264 82.633 14.336 ;
      RECT MASK 2 83.403 13.264 83.463 14.336 ;
      RECT MASK 2 84.233 13.264 84.293 14.336 ;
      RECT MASK 2 85.063 13.264 85.123 14.336 ;
      RECT MASK 2 85.893 13.264 85.953 14.336 ;
      RECT MASK 2 86.723 13.264 86.783 14.336 ;
      RECT MASK 2 87.553 13.264 87.613 14.336 ;
      RECT MASK 2 88.383 13.264 88.443 14.336 ;
      RECT MASK 2 89.213 13.264 89.273 14.336 ;
      RECT MASK 2 90.043 13.264 90.103 14.336 ;
      RECT MASK 2 90.873 13.264 90.933 14.336 ;
      RECT MASK 2 91.703 13.264 91.763 14.336 ;
      RECT MASK 2 92.533 13.264 92.593 14.336 ;
      RECT MASK 2 93.363 13.264 93.423 14.336 ;
      RECT MASK 2 94.193 13.264 94.253 14.336 ;
      RECT MASK 2 95.023 13.264 95.083 14.336 ;
      RECT MASK 2 95.853 13.264 95.913 14.336 ;
      RECT MASK 2 96.683 13.264 96.743 14.336 ;
      RECT MASK 2 97.513 13.264 97.573 14.336 ;
      RECT MASK 2 98.343 13.264 98.403 14.336 ;
      RECT MASK 2 99.173 13.264 99.233 14.336 ;
      RECT MASK 2 100.003 13.264 100.063 14.336 ;
      RECT MASK 2 100.833 13.264 100.893 14.336 ;
      RECT MASK 2 101.663 13.264 101.723 14.336 ;
      RECT MASK 2 102.493 13.264 102.553 14.336 ;
      RECT MASK 2 103.323 13.264 103.383 14.336 ;
      RECT MASK 2 104.153 13.264 104.213 14.336 ;
      RECT MASK 2 104.983 13.264 105.043 14.336 ;
      RECT MASK 2 105.813 13.264 105.873 14.336 ;
      RECT MASK 2 106.643 13.264 106.703 14.336 ;
      RECT MASK 2 107.473 13.264 107.533 14.336 ;
      RECT MASK 2 108.303 13.264 108.363 14.336 ;
      RECT MASK 2 109.133 13.264 109.193 14.336 ;
      RECT MASK 2 109.963 13.264 110.023 14.336 ;
      RECT MASK 2 110.793 13.264 110.853 14.336 ;
      RECT MASK 2 27.627 13.439 27.687 14.336 ;
      RECT MASK 2 40.907 13.439 40.967 14.336 ;
      RECT MASK 2 41.737 13.439 41.797 14.336 ;
      RECT MASK 2 62.653 13.439 62.713 14.336 ;
      RECT MASK 2 55.847 13.678 55.907 14.336 ;
      RECT MASK 2 30.117 14.14 30.177 14.336 ;
      RECT MASK 2 34.267 14.14 34.327 14.336 ;
      RECT MASK 2 35.097 14.14 35.157 14.336 ;
      RECT MASK 2 45.887 14.14 45.947 14.336 ;
      RECT MASK 2 60.163 14.14 60.223 14.336 ;
      RECT MASK 2 5.466 14.336 5.526 15.172 ;
      RECT MASK 2 5.798 14.336 5.858 15.172 ;
      RECT MASK 2 7.126 14.336 7.186 15.172 ;
      RECT MASK 2 7.458 14.336 7.518 15.172 ;
      RECT MASK 2 8.786 14.336 8.846 15.172 ;
      RECT MASK 2 9.118 14.336 9.178 15.172 ;
      RECT MASK 2 10.446 14.336 10.506 15.172 ;
      RECT MASK 2 10.778 14.336 10.838 15.172 ;
      RECT MASK 2 12.106 14.336 12.166 15.172 ;
      RECT MASK 2 12.438 14.336 12.498 15.172 ;
      RECT MASK 2 13.766 14.336 13.826 15.172 ;
      RECT MASK 2 14.098 14.336 14.158 15.172 ;
      RECT MASK 2 15.426 14.336 15.486 15.172 ;
      RECT MASK 2 15.758 14.336 15.818 15.172 ;
      RECT MASK 2 17.086 14.336 17.146 15.172 ;
      RECT MASK 2 17.418 14.336 17.478 15.172 ;
      RECT MASK 2 18.746 14.336 18.806 15.172 ;
      RECT MASK 2 19.078 14.336 19.138 15.172 ;
      RECT MASK 2 20.406 14.336 20.466 15.172 ;
      RECT MASK 2 20.738 14.336 20.798 15.172 ;
      RECT MASK 2 22.066 14.336 22.126 15.172 ;
      RECT MASK 2 22.398 14.336 22.458 15.172 ;
      RECT MASK 2 23.726 14.336 23.786 15.172 ;
      RECT MASK 2 24.058 14.336 24.118 15.172 ;
      RECT MASK 2 25.386 14.336 25.446 15.172 ;
      RECT MASK 2 25.718 14.336 25.778 15.172 ;
      RECT MASK 2 27.046 14.336 27.106 15.172 ;
      RECT MASK 2 27.378 14.336 27.438 15.172 ;
      RECT MASK 2 28.706 14.336 28.766 15.172 ;
      RECT MASK 2 29.038 14.336 29.098 15.172 ;
      RECT MASK 2 30.366 14.336 30.426 15.172 ;
      RECT MASK 2 30.698 14.336 30.758 15.172 ;
      RECT MASK 2 32.026 14.336 32.086 15.172 ;
      RECT MASK 2 32.358 14.336 32.418 15.172 ;
      RECT MASK 2 33.686 14.336 33.746 15.172 ;
      RECT MASK 2 34.018 14.336 34.078 15.172 ;
      RECT MASK 2 35.346 14.336 35.406 15.172 ;
      RECT MASK 2 35.678 14.336 35.738 15.172 ;
      RECT MASK 2 37.006 14.336 37.066 15.172 ;
      RECT MASK 2 37.338 14.336 37.398 15.172 ;
      RECT MASK 2 38.666 14.336 38.726 15.172 ;
      RECT MASK 2 38.998 14.336 39.058 15.172 ;
      RECT MASK 2 40.326 14.336 40.386 15.172 ;
      RECT MASK 2 40.658 14.336 40.718 15.172 ;
      RECT MASK 2 41.986 14.336 42.046 15.172 ;
      RECT MASK 2 42.318 14.336 42.378 15.172 ;
      RECT MASK 2 43.646 14.336 43.706 15.172 ;
      RECT MASK 2 43.978 14.336 44.038 15.172 ;
      RECT MASK 2 45.306 14.336 45.366 15.172 ;
      RECT MASK 2 45.638 14.336 45.698 15.172 ;
      RECT MASK 2 46.966 14.336 47.026 15.172 ;
      RECT MASK 2 47.298 14.336 47.358 15.172 ;
      RECT MASK 2 48.626 14.336 48.686 15.172 ;
      RECT MASK 2 48.958 14.336 49.018 15.172 ;
      RECT MASK 2 50.286 14.336 50.346 15.172 ;
      RECT MASK 2 50.618 14.336 50.678 15.172 ;
      RECT MASK 2 51.946 14.336 52.006 15.172 ;
      RECT MASK 2 52.278 14.336 52.338 15.172 ;
      RECT MASK 2 53.606 14.336 53.666 15.172 ;
      RECT MASK 2 53.938 14.336 53.998 15.172 ;
      RECT MASK 2 55.266 14.336 55.326 15.172 ;
      RECT MASK 2 55.598 14.336 55.658 15.172 ;
      RECT MASK 2 57.092 14.336 57.152 15.172 ;
      RECT MASK 2 57.424 14.336 57.484 15.172 ;
      RECT MASK 2 58.752 14.336 58.812 15.172 ;
      RECT MASK 2 59.084 14.336 59.144 15.172 ;
      RECT MASK 2 60.412 14.336 60.472 15.172 ;
      RECT MASK 2 60.744 14.336 60.804 15.172 ;
      RECT MASK 2 62.072 14.336 62.132 15.172 ;
      RECT MASK 2 62.404 14.336 62.464 15.172 ;
      RECT MASK 2 63.732 14.336 63.792 15.172 ;
      RECT MASK 2 64.064 14.336 64.124 15.172 ;
      RECT MASK 2 65.392 14.336 65.452 15.172 ;
      RECT MASK 2 65.724 14.336 65.784 15.172 ;
      RECT MASK 2 67.052 14.336 67.112 15.172 ;
      RECT MASK 2 67.384 14.336 67.444 15.172 ;
      RECT MASK 2 68.712 14.336 68.772 15.172 ;
      RECT MASK 2 69.044 14.336 69.104 15.172 ;
      RECT MASK 2 70.372 14.336 70.432 15.172 ;
      RECT MASK 2 70.704 14.336 70.764 15.172 ;
      RECT MASK 2 72.032 14.336 72.092 15.172 ;
      RECT MASK 2 72.364 14.336 72.424 15.172 ;
      RECT MASK 2 73.692 14.336 73.752 15.172 ;
      RECT MASK 2 74.024 14.336 74.084 15.172 ;
      RECT MASK 2 75.352 14.336 75.412 15.172 ;
      RECT MASK 2 75.684 14.336 75.744 15.172 ;
      RECT MASK 2 77.012 14.336 77.072 15.172 ;
      RECT MASK 2 77.344 14.336 77.404 15.172 ;
      RECT MASK 2 78.672 14.336 78.732 15.172 ;
      RECT MASK 2 79.004 14.336 79.064 15.172 ;
      RECT MASK 2 80.332 14.336 80.392 15.172 ;
      RECT MASK 2 80.664 14.336 80.724 15.172 ;
      RECT MASK 2 81.992 14.336 82.052 15.172 ;
      RECT MASK 2 82.324 14.336 82.384 15.172 ;
      RECT MASK 2 83.652 14.336 83.712 15.172 ;
      RECT MASK 2 83.984 14.336 84.044 15.172 ;
      RECT MASK 2 85.312 14.336 85.372 15.172 ;
      RECT MASK 2 85.644 14.336 85.704 15.172 ;
      RECT MASK 2 86.972 14.336 87.032 15.172 ;
      RECT MASK 2 87.304 14.336 87.364 15.172 ;
      RECT MASK 2 88.632 14.336 88.692 15.172 ;
      RECT MASK 2 88.964 14.336 89.024 15.172 ;
      RECT MASK 2 90.292 14.336 90.352 15.172 ;
      RECT MASK 2 90.624 14.336 90.684 15.172 ;
      RECT MASK 2 91.952 14.336 92.012 15.172 ;
      RECT MASK 2 92.284 14.336 92.344 15.172 ;
      RECT MASK 2 93.612 14.336 93.672 15.172 ;
      RECT MASK 2 93.944 14.336 94.004 15.172 ;
      RECT MASK 2 95.272 14.336 95.332 15.172 ;
      RECT MASK 2 95.604 14.336 95.664 15.172 ;
      RECT MASK 2 96.932 14.336 96.992 15.172 ;
      RECT MASK 2 97.264 14.336 97.324 15.172 ;
      RECT MASK 2 98.592 14.336 98.652 15.172 ;
      RECT MASK 2 98.924 14.336 98.984 15.172 ;
      RECT MASK 2 100.252 14.336 100.312 15.172 ;
      RECT MASK 2 100.584 14.336 100.644 15.172 ;
      RECT MASK 2 101.912 14.336 101.972 15.172 ;
      RECT MASK 2 102.244 14.336 102.304 15.172 ;
      RECT MASK 2 103.572 14.336 103.632 15.172 ;
      RECT MASK 2 103.904 14.336 103.964 15.172 ;
      RECT MASK 2 105.232 14.336 105.292 15.172 ;
      RECT MASK 2 105.564 14.336 105.624 15.172 ;
      RECT MASK 2 106.892 14.336 106.952 15.172 ;
      RECT MASK 2 107.224 14.336 107.284 15.172 ;
      RECT MASK 2 108.552 14.336 108.612 15.172 ;
      RECT MASK 2 108.884 14.336 108.944 15.172 ;
      RECT MASK 2 110.212 14.336 110.272 15.172 ;
      RECT MASK 2 110.544 14.336 110.604 15.172 ;
      RECT MASK 2 4.387 14.9225 4.447 16.5175 ;
      RECT MASK 2 111.623 14.9225 111.683 16.5175 ;
      RECT MASK 2 58.088 15.055 58.148 17.429 ;
      RECT MASK 2 5.217 15.184 5.277 16.256 ;
      RECT MASK 2 6.047 15.184 6.107 16.256 ;
      RECT MASK 2 6.877 15.184 6.937 16.256 ;
      RECT MASK 2 7.707 15.184 7.767 16.256 ;
      RECT MASK 2 8.537 15.184 8.597 16.256 ;
      RECT MASK 2 9.367 15.184 9.427 16.256 ;
      RECT MASK 2 10.197 15.184 10.257 16.256 ;
      RECT MASK 2 11.027 15.184 11.087 16.256 ;
      RECT MASK 2 11.857 15.184 11.917 16.256 ;
      RECT MASK 2 12.687 15.184 12.747 16.256 ;
      RECT MASK 2 13.517 15.184 13.577 16.256 ;
      RECT MASK 2 14.347 15.184 14.407 16.256 ;
      RECT MASK 2 15.177 15.184 15.237 16.256 ;
      RECT MASK 2 16.007 15.184 16.067 16.256 ;
      RECT MASK 2 16.837 15.184 16.897 16.256 ;
      RECT MASK 2 17.667 15.184 17.727 16.256 ;
      RECT MASK 2 18.497 15.184 18.557 16.256 ;
      RECT MASK 2 19.327 15.184 19.387 16.256 ;
      RECT MASK 2 20.157 15.184 20.217 16.256 ;
      RECT MASK 2 20.987 15.184 21.047 16.256 ;
      RECT MASK 2 21.817 15.184 21.877 16.256 ;
      RECT MASK 2 22.647 15.184 22.707 16.256 ;
      RECT MASK 2 23.477 15.184 23.537 16.256 ;
      RECT MASK 2 24.307 15.184 24.367 16.256 ;
      RECT MASK 2 25.137 15.184 25.197 16.256 ;
      RECT MASK 2 25.967 15.184 26.027 16.256 ;
      RECT MASK 2 26.797 15.184 26.857 16.256 ;
      RECT MASK 2 27.627 15.184 27.687 16.256 ;
      RECT MASK 2 28.457 15.184 28.517 16.256 ;
      RECT MASK 2 29.287 15.184 29.347 16.256 ;
      RECT MASK 2 30.117 15.184 30.177 16.256 ;
      RECT MASK 2 30.947 15.184 31.007 16.256 ;
      RECT MASK 2 31.777 15.184 31.837 16.256 ;
      RECT MASK 2 32.607 15.184 32.667 16.256 ;
      RECT MASK 2 33.437 15.184 33.497 16.256 ;
      RECT MASK 2 34.267 15.184 34.327 16.256 ;
      RECT MASK 2 35.097 15.184 35.157 16.256 ;
      RECT MASK 2 35.927 15.184 35.987 16.256 ;
      RECT MASK 2 36.757 15.184 36.817 16.256 ;
      RECT MASK 2 37.587 15.184 37.647 16.256 ;
      RECT MASK 2 38.417 15.184 38.477 16.256 ;
      RECT MASK 2 39.247 15.184 39.307 16.256 ;
      RECT MASK 2 40.077 15.184 40.137 16.256 ;
      RECT MASK 2 40.907 15.184 40.967 16.256 ;
      RECT MASK 2 41.737 15.184 41.797 16.256 ;
      RECT MASK 2 42.567 15.184 42.627 16.256 ;
      RECT MASK 2 43.397 15.184 43.457 16.256 ;
      RECT MASK 2 44.227 15.184 44.287 16.256 ;
      RECT MASK 2 45.057 15.184 45.117 16.256 ;
      RECT MASK 2 45.887 15.184 45.947 16.256 ;
      RECT MASK 2 46.717 15.184 46.777 16.256 ;
      RECT MASK 2 47.547 15.184 47.607 16.256 ;
      RECT MASK 2 48.377 15.184 48.437 16.256 ;
      RECT MASK 2 49.207 15.184 49.267 16.256 ;
      RECT MASK 2 50.037 15.184 50.097 16.256 ;
      RECT MASK 2 50.867 15.184 50.927 16.256 ;
      RECT MASK 2 51.697 15.184 51.757 16.256 ;
      RECT MASK 2 52.527 15.184 52.587 16.256 ;
      RECT MASK 2 53.357 15.184 53.417 16.256 ;
      RECT MASK 2 54.187 15.184 54.247 16.256 ;
      RECT MASK 2 55.017 15.184 55.077 16.256 ;
      RECT MASK 2 55.847 15.184 55.907 16.256 ;
      RECT MASK 2 56.823 15.184 56.923 16.256 ;
      RECT MASK 2 57.653 15.184 57.753 16.256 ;
      RECT MASK 2 58.483 15.184 58.583 16.256 ;
      RECT MASK 2 59.313 15.184 59.413 16.256 ;
      RECT MASK 2 60.143 15.184 60.243 16.256 ;
      RECT MASK 2 60.973 15.184 61.073 16.256 ;
      RECT MASK 2 61.823 15.184 61.883 16.256 ;
      RECT MASK 2 62.653 15.184 62.713 16.256 ;
      RECT MASK 2 63.483 15.184 63.543 16.256 ;
      RECT MASK 2 64.313 15.184 64.373 16.256 ;
      RECT MASK 2 65.143 15.184 65.203 16.256 ;
      RECT MASK 2 65.973 15.184 66.033 16.256 ;
      RECT MASK 2 66.803 15.184 66.863 16.256 ;
      RECT MASK 2 67.633 15.184 67.693 16.256 ;
      RECT MASK 2 68.463 15.184 68.523 16.256 ;
      RECT MASK 2 69.293 15.184 69.353 16.256 ;
      RECT MASK 2 70.123 15.184 70.183 16.256 ;
      RECT MASK 2 70.953 15.184 71.013 16.256 ;
      RECT MASK 2 71.783 15.184 71.843 16.256 ;
      RECT MASK 2 72.613 15.184 72.673 16.256 ;
      RECT MASK 2 73.443 15.184 73.503 16.256 ;
      RECT MASK 2 74.273 15.184 74.333 16.256 ;
      RECT MASK 2 75.103 15.184 75.163 16.256 ;
      RECT MASK 2 75.933 15.184 75.993 16.256 ;
      RECT MASK 2 76.763 15.184 76.823 16.256 ;
      RECT MASK 2 77.593 15.184 77.653 16.256 ;
      RECT MASK 2 78.423 15.184 78.483 16.256 ;
      RECT MASK 2 79.253 15.184 79.313 16.256 ;
      RECT MASK 2 80.083 15.184 80.143 16.256 ;
      RECT MASK 2 80.913 15.184 80.973 16.256 ;
      RECT MASK 2 81.743 15.184 81.803 16.256 ;
      RECT MASK 2 82.573 15.184 82.633 16.256 ;
      RECT MASK 2 83.403 15.184 83.463 16.256 ;
      RECT MASK 2 84.233 15.184 84.293 16.256 ;
      RECT MASK 2 85.063 15.184 85.123 16.256 ;
      RECT MASK 2 85.893 15.184 85.953 16.256 ;
      RECT MASK 2 86.723 15.184 86.783 16.256 ;
      RECT MASK 2 87.553 15.184 87.613 16.256 ;
      RECT MASK 2 88.383 15.184 88.443 16.256 ;
      RECT MASK 2 89.213 15.184 89.273 16.256 ;
      RECT MASK 2 90.043 15.184 90.103 16.256 ;
      RECT MASK 2 90.873 15.184 90.933 16.256 ;
      RECT MASK 2 91.703 15.184 91.763 16.256 ;
      RECT MASK 2 92.533 15.184 92.593 16.256 ;
      RECT MASK 2 93.363 15.184 93.423 16.256 ;
      RECT MASK 2 94.193 15.184 94.253 16.256 ;
      RECT MASK 2 95.023 15.184 95.083 16.256 ;
      RECT MASK 2 95.853 15.184 95.913 16.256 ;
      RECT MASK 2 96.683 15.184 96.743 16.256 ;
      RECT MASK 2 97.513 15.184 97.573 16.256 ;
      RECT MASK 2 98.343 15.184 98.403 16.256 ;
      RECT MASK 2 99.173 15.184 99.233 16.256 ;
      RECT MASK 2 100.003 15.184 100.063 16.256 ;
      RECT MASK 2 100.833 15.184 100.893 16.256 ;
      RECT MASK 2 101.663 15.184 101.723 16.256 ;
      RECT MASK 2 102.493 15.184 102.553 16.256 ;
      RECT MASK 2 103.323 15.184 103.383 16.256 ;
      RECT MASK 2 104.153 15.184 104.213 16.256 ;
      RECT MASK 2 104.983 15.184 105.043 16.256 ;
      RECT MASK 2 105.813 15.184 105.873 16.256 ;
      RECT MASK 2 106.643 15.184 106.703 16.256 ;
      RECT MASK 2 107.473 15.184 107.533 16.256 ;
      RECT MASK 2 108.303 15.184 108.363 16.256 ;
      RECT MASK 2 109.133 15.184 109.193 16.256 ;
      RECT MASK 2 109.963 15.184 110.023 16.256 ;
      RECT MASK 2 110.793 15.184 110.853 16.256 ;
      RECT MASK 2 5.466 16.268 5.526 17.104 ;
      RECT MASK 2 5.798 16.268 5.858 17.104 ;
      RECT MASK 2 7.126 16.268 7.186 17.104 ;
      RECT MASK 2 7.458 16.268 7.518 17.104 ;
      RECT MASK 2 8.786 16.268 8.846 17.104 ;
      RECT MASK 2 9.118 16.268 9.178 17.104 ;
      RECT MASK 2 10.446 16.268 10.506 17.104 ;
      RECT MASK 2 10.778 16.268 10.838 17.104 ;
      RECT MASK 2 12.106 16.268 12.166 17.104 ;
      RECT MASK 2 12.438 16.268 12.498 17.104 ;
      RECT MASK 2 13.766 16.268 13.826 17.104 ;
      RECT MASK 2 14.098 16.268 14.158 17.104 ;
      RECT MASK 2 15.426 16.268 15.486 17.104 ;
      RECT MASK 2 15.758 16.268 15.818 17.104 ;
      RECT MASK 2 17.086 16.268 17.146 17.104 ;
      RECT MASK 2 17.418 16.268 17.478 17.104 ;
      RECT MASK 2 18.746 16.268 18.806 17.104 ;
      RECT MASK 2 19.078 16.268 19.138 17.104 ;
      RECT MASK 2 20.406 16.268 20.466 17.104 ;
      RECT MASK 2 20.738 16.268 20.798 17.104 ;
      RECT MASK 2 22.066 16.268 22.126 17.104 ;
      RECT MASK 2 22.398 16.268 22.458 17.104 ;
      RECT MASK 2 23.726 16.268 23.786 17.104 ;
      RECT MASK 2 24.058 16.268 24.118 17.104 ;
      RECT MASK 2 25.386 16.268 25.446 17.104 ;
      RECT MASK 2 25.718 16.268 25.778 17.104 ;
      RECT MASK 2 27.046 16.268 27.106 17.104 ;
      RECT MASK 2 27.378 16.268 27.438 17.104 ;
      RECT MASK 2 28.706 16.268 28.766 17.104 ;
      RECT MASK 2 29.038 16.268 29.098 17.104 ;
      RECT MASK 2 30.366 16.268 30.426 17.104 ;
      RECT MASK 2 30.698 16.268 30.758 17.104 ;
      RECT MASK 2 32.026 16.268 32.086 17.104 ;
      RECT MASK 2 32.358 16.268 32.418 17.104 ;
      RECT MASK 2 33.686 16.268 33.746 17.104 ;
      RECT MASK 2 34.018 16.268 34.078 17.104 ;
      RECT MASK 2 35.346 16.268 35.406 17.104 ;
      RECT MASK 2 35.678 16.268 35.738 17.104 ;
      RECT MASK 2 37.006 16.268 37.066 17.104 ;
      RECT MASK 2 37.338 16.268 37.398 17.104 ;
      RECT MASK 2 38.666 16.268 38.726 17.104 ;
      RECT MASK 2 38.998 16.268 39.058 17.104 ;
      RECT MASK 2 40.326 16.268 40.386 17.104 ;
      RECT MASK 2 40.658 16.268 40.718 17.104 ;
      RECT MASK 2 41.986 16.268 42.046 17.104 ;
      RECT MASK 2 42.318 16.268 42.378 17.104 ;
      RECT MASK 2 43.646 16.268 43.706 17.104 ;
      RECT MASK 2 43.978 16.268 44.038 17.104 ;
      RECT MASK 2 45.306 16.268 45.366 17.104 ;
      RECT MASK 2 45.638 16.268 45.698 17.104 ;
      RECT MASK 2 46.966 16.268 47.026 17.104 ;
      RECT MASK 2 47.298 16.268 47.358 17.104 ;
      RECT MASK 2 48.626 16.268 48.686 17.104 ;
      RECT MASK 2 48.958 16.268 49.018 17.104 ;
      RECT MASK 2 50.286 16.268 50.346 17.104 ;
      RECT MASK 2 50.618 16.268 50.678 17.104 ;
      RECT MASK 2 51.946 16.268 52.006 17.104 ;
      RECT MASK 2 52.278 16.268 52.338 17.104 ;
      RECT MASK 2 53.606 16.268 53.666 17.104 ;
      RECT MASK 2 53.938 16.268 53.998 17.104 ;
      RECT MASK 2 55.266 16.268 55.326 17.104 ;
      RECT MASK 2 55.598 16.268 55.658 17.104 ;
      RECT MASK 2 57.092 16.268 57.152 17.104 ;
      RECT MASK 2 57.424 16.268 57.484 17.104 ;
      RECT MASK 2 58.752 16.268 58.812 17.104 ;
      RECT MASK 2 59.084 16.268 59.144 17.104 ;
      RECT MASK 2 60.412 16.268 60.472 17.104 ;
      RECT MASK 2 60.744 16.268 60.804 17.104 ;
      RECT MASK 2 62.072 16.268 62.132 17.104 ;
      RECT MASK 2 62.404 16.268 62.464 17.104 ;
      RECT MASK 2 63.732 16.268 63.792 17.104 ;
      RECT MASK 2 64.064 16.268 64.124 17.104 ;
      RECT MASK 2 65.392 16.268 65.452 17.104 ;
      RECT MASK 2 65.724 16.268 65.784 17.104 ;
      RECT MASK 2 67.052 16.268 67.112 17.104 ;
      RECT MASK 2 67.384 16.268 67.444 17.104 ;
      RECT MASK 2 68.712 16.268 68.772 17.104 ;
      RECT MASK 2 69.044 16.268 69.104 17.104 ;
      RECT MASK 2 70.372 16.268 70.432 17.104 ;
      RECT MASK 2 70.704 16.268 70.764 17.104 ;
      RECT MASK 2 72.032 16.268 72.092 17.104 ;
      RECT MASK 2 72.364 16.268 72.424 17.104 ;
      RECT MASK 2 73.692 16.268 73.752 17.104 ;
      RECT MASK 2 74.024 16.268 74.084 17.104 ;
      RECT MASK 2 75.352 16.268 75.412 17.104 ;
      RECT MASK 2 75.684 16.268 75.744 17.104 ;
      RECT MASK 2 77.012 16.268 77.072 17.104 ;
      RECT MASK 2 77.344 16.268 77.404 17.104 ;
      RECT MASK 2 78.672 16.268 78.732 17.104 ;
      RECT MASK 2 79.004 16.268 79.064 17.104 ;
      RECT MASK 2 80.332 16.268 80.392 17.104 ;
      RECT MASK 2 80.664 16.268 80.724 17.104 ;
      RECT MASK 2 81.992 16.268 82.052 17.104 ;
      RECT MASK 2 82.324 16.268 82.384 17.104 ;
      RECT MASK 2 83.652 16.268 83.712 17.104 ;
      RECT MASK 2 83.984 16.268 84.044 17.104 ;
      RECT MASK 2 85.312 16.268 85.372 17.104 ;
      RECT MASK 2 85.644 16.268 85.704 17.104 ;
      RECT MASK 2 86.972 16.268 87.032 17.104 ;
      RECT MASK 2 87.304 16.268 87.364 17.104 ;
      RECT MASK 2 88.632 16.268 88.692 17.104 ;
      RECT MASK 2 88.964 16.268 89.024 17.104 ;
      RECT MASK 2 90.292 16.268 90.352 17.104 ;
      RECT MASK 2 90.624 16.268 90.684 17.104 ;
      RECT MASK 2 91.952 16.268 92.012 17.104 ;
      RECT MASK 2 92.284 16.268 92.344 17.104 ;
      RECT MASK 2 93.612 16.268 93.672 17.104 ;
      RECT MASK 2 93.944 16.268 94.004 17.104 ;
      RECT MASK 2 95.272 16.268 95.332 17.104 ;
      RECT MASK 2 95.604 16.268 95.664 17.104 ;
      RECT MASK 2 96.932 16.268 96.992 17.104 ;
      RECT MASK 2 97.264 16.268 97.324 17.104 ;
      RECT MASK 2 98.592 16.268 98.652 17.104 ;
      RECT MASK 2 98.924 16.268 98.984 17.104 ;
      RECT MASK 2 100.252 16.268 100.312 17.104 ;
      RECT MASK 2 100.584 16.268 100.644 17.104 ;
      RECT MASK 2 101.912 16.268 101.972 17.104 ;
      RECT MASK 2 102.244 16.268 102.304 17.104 ;
      RECT MASK 2 103.572 16.268 103.632 17.104 ;
      RECT MASK 2 103.904 16.268 103.964 17.104 ;
      RECT MASK 2 105.232 16.268 105.292 17.104 ;
      RECT MASK 2 105.564 16.268 105.624 17.104 ;
      RECT MASK 2 106.892 16.268 106.952 17.104 ;
      RECT MASK 2 107.224 16.268 107.284 17.104 ;
      RECT MASK 2 108.552 16.268 108.612 17.104 ;
      RECT MASK 2 108.884 16.268 108.944 17.104 ;
      RECT MASK 2 110.212 16.268 110.272 17.104 ;
      RECT MASK 2 110.544 16.268 110.604 17.104 ;
      RECT MASK 2 23.8885 16.981 23.9485 17.429 ;
      RECT MASK 2 5.217 17.104 5.277 17.76 ;
      RECT MASK 2 6.047 17.104 6.107 17.76 ;
      RECT MASK 2 6.877 17.104 6.937 17.76 ;
      RECT MASK 2 7.707 17.104 7.767 17.76 ;
      RECT MASK 2 8.537 17.104 8.597 17.76 ;
      RECT MASK 2 9.367 17.104 9.427 17.76 ;
      RECT MASK 2 10.197 17.104 10.257 17.76 ;
      RECT MASK 2 11.027 17.104 11.087 17.76 ;
      RECT MASK 2 11.857 17.104 11.917 17.76 ;
      RECT MASK 2 12.687 17.104 12.747 17.76 ;
      RECT MASK 2 13.517 17.104 13.577 17.76 ;
      RECT MASK 2 14.347 17.104 14.407 17.76 ;
      RECT MASK 2 15.177 17.104 15.237 17.76 ;
      RECT MASK 2 16.007 17.104 16.067 17.76 ;
      RECT MASK 2 16.837 17.104 16.897 17.76 ;
      RECT MASK 2 17.667 17.104 17.727 17.76 ;
      RECT MASK 2 18.497 17.104 18.557 17.76 ;
      RECT MASK 2 19.327 17.104 19.387 17.76 ;
      RECT MASK 2 20.157 17.104 20.217 17.76 ;
      RECT MASK 2 20.987 17.104 21.047 17.76 ;
      RECT MASK 2 21.817 17.104 21.877 17.76 ;
      RECT MASK 2 22.647 17.104 22.707 17.76 ;
      RECT MASK 2 23.477 17.104 23.537 17.76 ;
      RECT MASK 2 24.307 17.104 24.367 17.76 ;
      RECT MASK 2 25.137 17.104 25.197 17.76 ;
      RECT MASK 2 25.967 17.104 26.027 17.76 ;
      RECT MASK 2 26.797 17.104 26.857 17.76 ;
      RECT MASK 2 27.627 17.104 27.687 17.76 ;
      RECT MASK 2 28.457 17.104 28.517 17.76 ;
      RECT MASK 2 29.287 17.104 29.347 17.76 ;
      RECT MASK 2 30.117 17.104 30.177 17.76 ;
      RECT MASK 2 30.947 17.104 31.007 17.76 ;
      RECT MASK 2 31.777 17.104 31.837 17.76 ;
      RECT MASK 2 32.607 17.104 32.667 17.76 ;
      RECT MASK 2 33.437 17.104 33.497 17.76 ;
      RECT MASK 2 34.267 17.104 34.327 17.76 ;
      RECT MASK 2 35.097 17.104 35.157 17.76 ;
      RECT MASK 2 35.927 17.104 35.987 17.76 ;
      RECT MASK 2 36.757 17.104 36.817 17.76 ;
      RECT MASK 2 37.587 17.104 37.647 17.76 ;
      RECT MASK 2 38.417 17.104 38.477 17.76 ;
      RECT MASK 2 39.247 17.104 39.307 17.76 ;
      RECT MASK 2 40.077 17.104 40.137 17.76 ;
      RECT MASK 2 40.907 17.104 40.967 17.76 ;
      RECT MASK 2 41.737 17.104 41.797 17.76 ;
      RECT MASK 2 42.567 17.104 42.627 17.76 ;
      RECT MASK 2 43.397 17.104 43.457 17.76 ;
      RECT MASK 2 44.227 17.104 44.287 17.76 ;
      RECT MASK 2 45.057 17.104 45.117 17.76 ;
      RECT MASK 2 45.887 17.104 45.947 17.76 ;
      RECT MASK 2 46.717 17.104 46.777 17.76 ;
      RECT MASK 2 47.547 17.104 47.607 17.76 ;
      RECT MASK 2 48.377 17.104 48.437 17.76 ;
      RECT MASK 2 49.207 17.104 49.267 17.76 ;
      RECT MASK 2 50.037 17.104 50.097 17.76 ;
      RECT MASK 2 50.867 17.104 50.927 17.76 ;
      RECT MASK 2 51.697 17.104 51.757 17.76 ;
      RECT MASK 2 52.527 17.104 52.587 17.76 ;
      RECT MASK 2 53.357 17.104 53.417 17.76 ;
      RECT MASK 2 54.187 17.104 54.247 17.76 ;
      RECT MASK 2 55.017 17.104 55.077 17.76 ;
      RECT MASK 2 55.847 17.104 55.907 17.76 ;
      RECT MASK 2 56.843 17.104 56.903 17.76 ;
      RECT MASK 2 57.673 17.104 57.733 17.76 ;
      RECT MASK 2 58.503 17.104 58.563 17.76 ;
      RECT MASK 2 59.333 17.104 59.393 17.76 ;
      RECT MASK 2 60.163 17.104 60.223 17.76 ;
      RECT MASK 2 60.993 17.104 61.053 17.76 ;
      RECT MASK 2 61.823 17.104 61.883 17.76 ;
      RECT MASK 2 62.653 17.104 62.713 17.76 ;
      RECT MASK 2 63.483 17.104 63.543 17.76 ;
      RECT MASK 2 64.313 17.104 64.373 17.76 ;
      RECT MASK 2 65.143 17.104 65.203 17.76 ;
      RECT MASK 2 65.963 17.104 66.043 17.76 ;
      RECT MASK 2 66.793 17.104 66.873 17.76 ;
      RECT MASK 2 67.633 17.104 67.693 17.76 ;
      RECT MASK 2 68.463 17.104 68.523 17.76 ;
      RECT MASK 2 69.293 17.104 69.353 17.76 ;
      RECT MASK 2 70.123 17.104 70.183 17.76 ;
      RECT MASK 2 70.953 17.104 71.013 17.76 ;
      RECT MASK 2 71.783 17.104 71.843 17.76 ;
      RECT MASK 2 72.613 17.104 72.673 17.76 ;
      RECT MASK 2 73.443 17.104 73.503 17.76 ;
      RECT MASK 2 74.273 17.104 74.333 17.76 ;
      RECT MASK 2 75.103 17.104 75.163 17.76 ;
      RECT MASK 2 75.933 17.104 75.993 17.76 ;
      RECT MASK 2 76.763 17.104 76.823 17.76 ;
      RECT MASK 2 77.593 17.104 77.653 17.76 ;
      RECT MASK 2 78.423 17.104 78.483 17.76 ;
      RECT MASK 2 79.253 17.104 79.313 17.76 ;
      RECT MASK 2 80.083 17.104 80.143 17.76 ;
      RECT MASK 2 80.913 17.104 80.973 17.76 ;
      RECT MASK 2 81.743 17.104 81.803 17.76 ;
      RECT MASK 2 82.573 17.104 82.633 17.76 ;
      RECT MASK 2 83.403 17.104 83.463 17.76 ;
      RECT MASK 2 84.233 17.104 84.293 17.76 ;
      RECT MASK 2 85.063 17.104 85.123 17.76 ;
      RECT MASK 2 85.893 17.104 85.953 17.76 ;
      RECT MASK 2 86.723 17.104 86.783 17.76 ;
      RECT MASK 2 87.553 17.104 87.613 17.76 ;
      RECT MASK 2 88.383 17.104 88.443 17.76 ;
      RECT MASK 2 89.213 17.104 89.273 17.76 ;
      RECT MASK 2 90.043 17.104 90.103 17.76 ;
      RECT MASK 2 90.873 17.104 90.933 17.76 ;
      RECT MASK 2 91.703 17.104 91.763 17.76 ;
      RECT MASK 2 92.533 17.104 92.593 17.76 ;
      RECT MASK 2 93.363 17.104 93.423 17.76 ;
      RECT MASK 2 94.193 17.104 94.253 17.76 ;
      RECT MASK 2 95.023 17.104 95.083 17.76 ;
      RECT MASK 2 95.853 17.104 95.913 17.76 ;
      RECT MASK 2 96.683 17.104 96.743 17.76 ;
      RECT MASK 2 97.513 17.104 97.573 17.76 ;
      RECT MASK 2 98.343 17.104 98.403 17.76 ;
      RECT MASK 2 99.173 17.104 99.233 17.76 ;
      RECT MASK 2 100.003 17.104 100.063 17.76 ;
      RECT MASK 2 100.833 17.104 100.893 17.76 ;
      RECT MASK 2 101.663 17.104 101.723 17.76 ;
      RECT MASK 2 102.493 17.104 102.553 17.76 ;
      RECT MASK 2 103.323 17.104 103.383 17.76 ;
      RECT MASK 2 104.153 17.104 104.213 17.76 ;
      RECT MASK 2 104.983 17.104 105.043 17.76 ;
      RECT MASK 2 105.813 17.104 105.873 17.76 ;
      RECT MASK 2 106.643 17.104 106.703 17.76 ;
      RECT MASK 2 107.473 17.104 107.533 17.76 ;
      RECT MASK 2 108.303 17.104 108.363 17.76 ;
      RECT MASK 2 109.133 17.104 109.193 17.76 ;
      RECT MASK 2 109.963 17.104 110.023 17.76 ;
      RECT MASK 2 110.793 17.104 110.853 17.76 ;
      RECT MASK 2 103.943 18.376 104.003 24.334 ;
      RECT MASK 2 5.914 18.739 5.974 21.9395 ;
      RECT MASK 2 6.246 18.739 6.306 21.738 ;
      RECT MASK 2 7.076 18.739 7.136 21.9395 ;
      RECT MASK 2 7.408 18.739 7.468 21.738 ;
      RECT MASK 2 8.238 18.739 8.298 21.9395 ;
      RECT MASK 2 8.57 18.739 8.63 21.738 ;
      RECT MASK 2 9.4 18.739 9.46 21.9395 ;
      RECT MASK 2 9.732 18.739 9.792 21.738 ;
      RECT MASK 2 12.532 18.739 12.592 21.9395 ;
      RECT MASK 2 12.864 18.739 12.924 21.738 ;
      RECT MASK 2 13.694 18.739 13.754 21.9395 ;
      RECT MASK 2 14.026 18.739 14.086 21.738 ;
      RECT MASK 2 14.856 18.739 14.916 21.9395 ;
      RECT MASK 2 15.188 18.739 15.248 21.738 ;
      RECT MASK 2 16.018 18.739 16.078 21.9395 ;
      RECT MASK 2 16.35 18.739 16.41 21.738 ;
      RECT MASK 2 19.15 18.739 19.21 21.9395 ;
      RECT MASK 2 19.482 18.739 19.542 21.738 ;
      RECT MASK 2 20.312 18.739 20.372 21.9395 ;
      RECT MASK 2 20.644 18.739 20.704 21.738 ;
      RECT MASK 2 21.474 18.739 21.534 21.9395 ;
      RECT MASK 2 21.806 18.739 21.866 21.738 ;
      RECT MASK 2 22.636 18.739 22.696 21.9395 ;
      RECT MASK 2 22.968 18.739 23.028 21.738 ;
      RECT MASK 2 25.768 18.739 25.828 21.9395 ;
      RECT MASK 2 26.1 18.739 26.16 21.738 ;
      RECT MASK 2 26.93 18.739 26.99 21.9395 ;
      RECT MASK 2 27.262 18.739 27.322 21.738 ;
      RECT MASK 2 28.092 18.739 28.152 21.9395 ;
      RECT MASK 2 28.424 18.739 28.484 21.738 ;
      RECT MASK 2 29.254 18.739 29.314 21.9395 ;
      RECT MASK 2 29.586 18.739 29.646 21.738 ;
      RECT MASK 2 32.386 18.739 32.446 21.9395 ;
      RECT MASK 2 32.718 18.739 32.778 21.738 ;
      RECT MASK 2 33.548 18.739 33.608 21.9395 ;
      RECT MASK 2 33.88 18.739 33.94 21.738 ;
      RECT MASK 2 34.71 18.739 34.77 21.9395 ;
      RECT MASK 2 35.042 18.739 35.102 21.738 ;
      RECT MASK 2 35.872 18.739 35.932 21.9395 ;
      RECT MASK 2 36.204 18.739 36.264 21.738 ;
      RECT MASK 2 39.004 18.739 39.064 21.9395 ;
      RECT MASK 2 39.336 18.739 39.396 21.738 ;
      RECT MASK 2 40.166 18.739 40.226 21.9395 ;
      RECT MASK 2 40.498 18.739 40.558 21.738 ;
      RECT MASK 2 41.328 18.739 41.388 21.9395 ;
      RECT MASK 2 41.66 18.739 41.72 21.738 ;
      RECT MASK 2 42.49 18.739 42.55 21.9395 ;
      RECT MASK 2 42.822 18.739 42.882 21.738 ;
      RECT MASK 2 45.622 18.739 45.682 21.9395 ;
      RECT MASK 2 45.954 18.739 46.014 21.738 ;
      RECT MASK 2 46.784 18.739 46.844 21.9395 ;
      RECT MASK 2 47.116 18.739 47.176 21.738 ;
      RECT MASK 2 47.946 18.739 48.006 21.9395 ;
      RECT MASK 2 48.278 18.739 48.338 21.738 ;
      RECT MASK 2 49.108 18.739 49.168 21.9395 ;
      RECT MASK 2 49.44 18.739 49.5 21.738 ;
      RECT MASK 2 52.24 18.739 52.3 21.9395 ;
      RECT MASK 2 52.572 18.739 52.632 21.738 ;
      RECT MASK 2 53.402 18.739 53.462 21.9395 ;
      RECT MASK 2 53.734 18.739 53.794 21.738 ;
      RECT MASK 2 54.564 18.739 54.624 21.9395 ;
      RECT MASK 2 54.896 18.739 54.956 21.738 ;
      RECT MASK 2 55.726 18.739 55.786 21.9395 ;
      RECT MASK 2 56.058 18.739 56.118 21.738 ;
      RECT MASK 2 58.858 18.739 58.918 21.9395 ;
      RECT MASK 2 59.19 18.739 59.25 21.738 ;
      RECT MASK 2 60.02 18.739 60.08 21.9395 ;
      RECT MASK 2 60.352 18.739 60.412 21.738 ;
      RECT MASK 2 61.182 18.739 61.242 21.9395 ;
      RECT MASK 2 61.514 18.739 61.574 21.738 ;
      RECT MASK 2 62.344 18.739 62.404 21.9395 ;
      RECT MASK 2 62.676 18.739 62.736 21.738 ;
      RECT MASK 2 65.476 18.739 65.536 21.9395 ;
      RECT MASK 2 65.808 18.739 65.868 21.738 ;
      RECT MASK 2 66.638 18.739 66.698 21.9395 ;
      RECT MASK 2 66.97 18.739 67.03 21.738 ;
      RECT MASK 2 67.8 18.739 67.86 21.9395 ;
      RECT MASK 2 68.132 18.739 68.192 21.738 ;
      RECT MASK 2 68.962 18.739 69.022 21.9395 ;
      RECT MASK 2 69.294 18.739 69.354 21.738 ;
      RECT MASK 2 72.094 18.739 72.154 21.9395 ;
      RECT MASK 2 72.426 18.739 72.486 21.738 ;
      RECT MASK 2 73.256 18.739 73.316 21.9395 ;
      RECT MASK 2 73.588 18.739 73.648 21.738 ;
      RECT MASK 2 74.418 18.739 74.478 21.9395 ;
      RECT MASK 2 74.75 18.739 74.81 21.738 ;
      RECT MASK 2 75.58 18.739 75.64 21.9395 ;
      RECT MASK 2 75.912 18.739 75.972 21.738 ;
      RECT MASK 2 78.712 18.739 78.772 21.9395 ;
      RECT MASK 2 79.044 18.739 79.104 21.738 ;
      RECT MASK 2 79.874 18.739 79.934 21.9395 ;
      RECT MASK 2 80.206 18.739 80.266 21.738 ;
      RECT MASK 2 81.036 18.739 81.096 21.9395 ;
      RECT MASK 2 81.368 18.739 81.428 21.738 ;
      RECT MASK 2 82.198 18.739 82.258 21.9395 ;
      RECT MASK 2 82.53 18.739 82.59 21.738 ;
      RECT MASK 2 85.33 18.739 85.39 21.9395 ;
      RECT MASK 2 85.662 18.739 85.722 21.738 ;
      RECT MASK 2 86.492 18.739 86.552 21.9395 ;
      RECT MASK 2 86.824 18.739 86.884 21.738 ;
      RECT MASK 2 87.654 18.739 87.714 21.9395 ;
      RECT MASK 2 87.986 18.739 88.046 21.738 ;
      RECT MASK 2 88.816 18.739 88.876 21.9395 ;
      RECT MASK 2 89.148 18.739 89.208 21.738 ;
      RECT MASK 2 91.948 18.739 92.008 21.9395 ;
      RECT MASK 2 92.28 18.739 92.34 21.738 ;
      RECT MASK 2 93.11 18.739 93.17 21.9395 ;
      RECT MASK 2 93.442 18.739 93.502 21.738 ;
      RECT MASK 2 94.272 18.739 94.332 21.9395 ;
      RECT MASK 2 94.604 18.739 94.664 21.738 ;
      RECT MASK 2 95.434 18.739 95.494 21.9395 ;
      RECT MASK 2 95.766 18.739 95.826 21.738 ;
      RECT MASK 2 98.566 18.739 98.626 21.9395 ;
      RECT MASK 2 98.898 18.739 98.958 21.738 ;
      RECT MASK 2 99.728 18.739 99.788 21.9395 ;
      RECT MASK 2 100.06 18.739 100.12 21.738 ;
      RECT MASK 2 100.89 18.739 100.95 21.9395 ;
      RECT MASK 2 101.222 18.739 101.282 21.738 ;
      RECT MASK 2 102.052 18.739 102.112 21.9395 ;
      RECT MASK 2 102.384 18.739 102.444 21.738 ;
      RECT MASK 2 105.184 18.739 105.244 21.9395 ;
      RECT MASK 2 105.516 18.739 105.576 21.738 ;
      RECT MASK 2 106.346 18.739 106.406 21.9395 ;
      RECT MASK 2 106.678 18.739 106.738 21.738 ;
      RECT MASK 2 107.508 18.739 107.568 21.9395 ;
      RECT MASK 2 107.84 18.739 107.9 21.738 ;
      RECT MASK 2 108.67 18.739 108.73 21.9395 ;
      RECT MASK 2 109.002 18.739 109.062 21.738 ;
      RECT MASK 2 2.362 19.56 2.422 24.53 ;
      RECT MASK 2 2.636 19.56 2.696 24.53 ;
      RECT MASK 2 2.91 19.56 2.97 24.53 ;
      RECT MASK 2 3.184 19.56 3.244 24.53 ;
      RECT MASK 2 3.458 19.56 3.518 24.53 ;
      RECT MASK 2 3.732 19.56 3.792 24.53 ;
      RECT MASK 2 5.499 19.818 5.559 21.6 ;
      RECT MASK 2 57.059 20.387 57.119 21.9635 ;
      RECT MASK 2 57.391 20.387 57.451 21.9635 ;
      RECT MASK 2 57.723 20.387 57.783 21.9635 ;
      RECT MASK 2 59.605 20.791 59.665 21.6 ;
      RECT MASK 2 58.443 20.8655 58.503 21.9635 ;
      RECT MASK 2 6.661 21.33 6.721 21.6 ;
      RECT MASK 2 7.823 21.33 7.883 21.6 ;
      RECT MASK 2 8.985 21.33 9.045 21.6 ;
      RECT MASK 2 10.147 21.33 10.207 21.6 ;
      RECT MASK 2 12.117 21.33 12.177 21.6 ;
      RECT MASK 2 13.279 21.33 13.339 21.6 ;
      RECT MASK 2 14.441 21.33 14.501 21.6 ;
      RECT MASK 2 15.603 21.33 15.663 21.6 ;
      RECT MASK 2 16.765 21.33 16.825 21.6 ;
      RECT MASK 2 18.735 21.33 18.795 21.6 ;
      RECT MASK 2 19.897 21.33 19.957 21.6 ;
      RECT MASK 2 21.059 21.33 21.119 21.6 ;
      RECT MASK 2 22.221 21.33 22.281 21.6 ;
      RECT MASK 2 23.383 21.33 23.443 21.6 ;
      RECT MASK 2 25.353 21.33 25.413 21.6 ;
      RECT MASK 2 26.515 21.33 26.575 21.6 ;
      RECT MASK 2 27.677 21.33 27.737 21.6 ;
      RECT MASK 2 28.839 21.33 28.899 21.6 ;
      RECT MASK 2 30.001 21.33 30.061 21.6 ;
      RECT MASK 2 31.971 21.33 32.031 21.6 ;
      RECT MASK 2 33.133 21.33 33.193 21.6 ;
      RECT MASK 2 34.295 21.33 34.355 21.6 ;
      RECT MASK 2 35.457 21.33 35.517 21.6 ;
      RECT MASK 2 36.619 21.33 36.679 21.6 ;
      RECT MASK 2 38.589 21.33 38.649 21.6 ;
      RECT MASK 2 39.751 21.33 39.811 21.6 ;
      RECT MASK 2 40.913 21.33 40.973 21.6 ;
      RECT MASK 2 42.075 21.33 42.135 21.6 ;
      RECT MASK 2 43.237 21.33 43.297 21.6 ;
      RECT MASK 2 45.207 21.33 45.267 21.6 ;
      RECT MASK 2 46.369 21.33 46.429 21.6 ;
      RECT MASK 2 47.531 21.33 47.591 21.6 ;
      RECT MASK 2 48.693 21.33 48.753 21.6 ;
      RECT MASK 2 49.855 21.33 49.915 21.6 ;
      RECT MASK 2 51.825 21.33 51.885 21.6 ;
      RECT MASK 2 52.987 21.33 53.047 21.6 ;
      RECT MASK 2 54.149 21.33 54.209 21.6 ;
      RECT MASK 2 55.311 21.33 55.371 21.6 ;
      RECT MASK 2 56.473 21.33 56.533 21.6 ;
      RECT MASK 2 60.767 21.33 60.827 21.6 ;
      RECT MASK 2 61.929 21.33 61.989 21.6 ;
      RECT MASK 2 63.091 21.33 63.151 21.6 ;
      RECT MASK 2 65.061 21.33 65.121 21.6 ;
      RECT MASK 2 66.223 21.33 66.283 21.6 ;
      RECT MASK 2 67.385 21.33 67.445 21.6 ;
      RECT MASK 2 68.547 21.33 68.607 21.6 ;
      RECT MASK 2 69.709 21.33 69.769 21.6 ;
      RECT MASK 2 71.679 21.33 71.739 21.6 ;
      RECT MASK 2 72.841 21.33 72.901 21.6 ;
      RECT MASK 2 74.003 21.33 74.063 21.6 ;
      RECT MASK 2 75.165 21.33 75.225 21.6 ;
      RECT MASK 2 76.327 21.33 76.387 21.6 ;
      RECT MASK 2 78.297 21.33 78.357 21.6 ;
      RECT MASK 2 79.459 21.33 79.519 21.6 ;
      RECT MASK 2 80.621 21.33 80.681 21.6 ;
      RECT MASK 2 81.783 21.33 81.843 21.6 ;
      RECT MASK 2 82.945 21.33 83.005 21.6 ;
      RECT MASK 2 84.915 21.33 84.975 21.6 ;
      RECT MASK 2 86.077 21.33 86.137 21.6 ;
      RECT MASK 2 87.239 21.33 87.299 21.6 ;
      RECT MASK 2 88.401 21.33 88.461 21.6 ;
      RECT MASK 2 89.563 21.33 89.623 21.6 ;
      RECT MASK 2 91.533 21.33 91.593 21.6 ;
      RECT MASK 2 92.695 21.33 92.755 21.6 ;
      RECT MASK 2 93.857 21.33 93.917 21.6 ;
      RECT MASK 2 95.019 21.33 95.079 21.6 ;
      RECT MASK 2 96.181 21.33 96.241 21.6 ;
      RECT MASK 2 98.151 21.33 98.211 21.6 ;
      RECT MASK 2 99.313 21.33 99.373 21.6 ;
      RECT MASK 2 100.475 21.33 100.535 21.6 ;
      RECT MASK 2 101.637 21.33 101.697 21.6 ;
      RECT MASK 2 102.799 21.33 102.859 21.6 ;
      RECT MASK 2 104.769 21.33 104.829 21.6 ;
      RECT MASK 2 105.931 21.33 105.991 21.6 ;
      RECT MASK 2 107.093 21.33 107.153 21.6 ;
      RECT MASK 2 108.255 21.33 108.315 21.6 ;
      RECT MASK 2 109.417 21.33 109.477 21.6 ;
      RECT MASK 2 17.097 21.335 17.157 23.545 ;
      RECT MASK 2 18.403 21.335 18.463 23.545 ;
      RECT MASK 2 5.655 22.0915 5.735 25.394 ;
      RECT MASK 2 5.987 22.0915 6.067 25.394 ;
      RECT MASK 2 6.319 22.0915 6.399 25.394 ;
      RECT MASK 2 6.817 22.0915 6.897 25.394 ;
      RECT MASK 2 7.149 22.0915 7.229 25.394 ;
      RECT MASK 2 7.481 22.0915 7.561 25.394 ;
      RECT MASK 2 7.979 22.0915 8.059 25.394 ;
      RECT MASK 2 8.311 22.0915 8.391 25.394 ;
      RECT MASK 2 8.643 22.0915 8.723 25.394 ;
      RECT MASK 2 9.141 22.0915 9.221 25.394 ;
      RECT MASK 2 9.473 22.0915 9.553 25.394 ;
      RECT MASK 2 9.805 22.0915 9.885 25.394 ;
      RECT MASK 2 12.273 22.0915 12.353 25.394 ;
      RECT MASK 2 12.605 22.0915 12.685 25.394 ;
      RECT MASK 2 12.937 22.0915 13.017 25.394 ;
      RECT MASK 2 13.435 22.0915 13.515 25.394 ;
      RECT MASK 2 13.767 22.0915 13.847 25.394 ;
      RECT MASK 2 14.099 22.0915 14.179 25.394 ;
      RECT MASK 2 14.597 22.0915 14.677 25.394 ;
      RECT MASK 2 14.929 22.0915 15.009 25.394 ;
      RECT MASK 2 15.261 22.0915 15.341 25.394 ;
      RECT MASK 2 15.759 22.0915 15.839 25.394 ;
      RECT MASK 2 16.091 22.0915 16.171 25.394 ;
      RECT MASK 2 16.423 22.0915 16.503 25.394 ;
      RECT MASK 2 18.891 22.0915 18.971 25.394 ;
      RECT MASK 2 19.223 22.0915 19.303 25.394 ;
      RECT MASK 2 19.555 22.0915 19.635 25.394 ;
      RECT MASK 2 20.053 22.0915 20.133 25.394 ;
      RECT MASK 2 20.385 22.0915 20.465 25.394 ;
      RECT MASK 2 20.717 22.0915 20.797 25.394 ;
      RECT MASK 2 21.215 22.0915 21.295 25.394 ;
      RECT MASK 2 21.547 22.0915 21.627 25.394 ;
      RECT MASK 2 21.879 22.0915 21.959 25.394 ;
      RECT MASK 2 22.377 22.0915 22.457 25.394 ;
      RECT MASK 2 22.709 22.0915 22.789 25.394 ;
      RECT MASK 2 23.041 22.0915 23.121 25.394 ;
      RECT MASK 2 25.509 22.0915 25.589 25.394 ;
      RECT MASK 2 25.841 22.0915 25.921 25.394 ;
      RECT MASK 2 26.173 22.0915 26.253 25.394 ;
      RECT MASK 2 26.671 22.0915 26.751 25.394 ;
      RECT MASK 2 27.003 22.0915 27.083 25.394 ;
      RECT MASK 2 27.335 22.0915 27.415 25.394 ;
      RECT MASK 2 27.833 22.0915 27.913 25.394 ;
      RECT MASK 2 28.165 22.0915 28.245 25.394 ;
      RECT MASK 2 28.497 22.0915 28.577 25.394 ;
      RECT MASK 2 28.995 22.0915 29.075 25.394 ;
      RECT MASK 2 29.327 22.0915 29.407 25.394 ;
      RECT MASK 2 29.659 22.0915 29.739 25.394 ;
      RECT MASK 2 32.127 22.0915 32.207 25.394 ;
      RECT MASK 2 32.459 22.0915 32.539 25.394 ;
      RECT MASK 2 32.791 22.0915 32.871 25.394 ;
      RECT MASK 2 33.289 22.0915 33.369 25.394 ;
      RECT MASK 2 33.621 22.0915 33.701 25.394 ;
      RECT MASK 2 33.953 22.0915 34.033 25.394 ;
      RECT MASK 2 34.451 22.0915 34.531 25.394 ;
      RECT MASK 2 34.783 22.0915 34.863 25.394 ;
      RECT MASK 2 35.115 22.0915 35.195 25.394 ;
      RECT MASK 2 35.613 22.0915 35.693 25.394 ;
      RECT MASK 2 35.945 22.0915 36.025 25.394 ;
      RECT MASK 2 36.277 22.0915 36.357 25.394 ;
      RECT MASK 2 38.745 22.0915 38.825 25.394 ;
      RECT MASK 2 39.077 22.0915 39.157 25.394 ;
      RECT MASK 2 39.409 22.0915 39.489 25.394 ;
      RECT MASK 2 39.907 22.0915 39.987 25.394 ;
      RECT MASK 2 40.239 22.0915 40.319 25.394 ;
      RECT MASK 2 40.571 22.0915 40.651 25.394 ;
      RECT MASK 2 41.069 22.0915 41.149 25.394 ;
      RECT MASK 2 41.401 22.0915 41.481 25.394 ;
      RECT MASK 2 41.733 22.0915 41.813 25.394 ;
      RECT MASK 2 42.231 22.0915 42.311 25.394 ;
      RECT MASK 2 42.563 22.0915 42.643 25.394 ;
      RECT MASK 2 42.895 22.0915 42.975 25.394 ;
      RECT MASK 2 45.363 22.0915 45.443 25.394 ;
      RECT MASK 2 45.695 22.0915 45.775 25.394 ;
      RECT MASK 2 46.027 22.0915 46.107 25.394 ;
      RECT MASK 2 46.525 22.0915 46.605 25.394 ;
      RECT MASK 2 46.857 22.0915 46.937 25.394 ;
      RECT MASK 2 47.189 22.0915 47.269 25.394 ;
      RECT MASK 2 47.687 22.0915 47.767 25.394 ;
      RECT MASK 2 48.019 22.0915 48.099 25.394 ;
      RECT MASK 2 48.351 22.0915 48.431 25.394 ;
      RECT MASK 2 48.849 22.0915 48.929 25.394 ;
      RECT MASK 2 49.181 22.0915 49.261 25.394 ;
      RECT MASK 2 49.513 22.0915 49.593 25.394 ;
      RECT MASK 2 51.981 22.0915 52.061 25.394 ;
      RECT MASK 2 52.313 22.0915 52.393 25.394 ;
      RECT MASK 2 52.645 22.0915 52.725 25.394 ;
      RECT MASK 2 53.143 22.0915 53.223 25.394 ;
      RECT MASK 2 53.475 22.0915 53.555 25.394 ;
      RECT MASK 2 53.807 22.0915 53.887 25.394 ;
      RECT MASK 2 54.305 22.0915 54.385 25.394 ;
      RECT MASK 2 54.637 22.0915 54.717 25.394 ;
      RECT MASK 2 54.969 22.0915 55.049 25.394 ;
      RECT MASK 2 55.467 22.0915 55.547 25.394 ;
      RECT MASK 2 55.799 22.0915 55.879 25.394 ;
      RECT MASK 2 56.131 22.0915 56.211 25.394 ;
      RECT MASK 2 58.599 22.0915 58.679 25.394 ;
      RECT MASK 2 58.931 22.0915 59.011 25.394 ;
      RECT MASK 2 59.263 22.0915 59.343 25.394 ;
      RECT MASK 2 59.761 22.0915 59.841 25.394 ;
      RECT MASK 2 60.093 22.0915 60.173 25.394 ;
      RECT MASK 2 60.425 22.0915 60.505 25.394 ;
      RECT MASK 2 60.923 22.0915 61.003 25.394 ;
      RECT MASK 2 61.255 22.0915 61.335 25.394 ;
      RECT MASK 2 61.587 22.0915 61.667 25.394 ;
      RECT MASK 2 62.085 22.0915 62.165 25.394 ;
      RECT MASK 2 62.417 22.0915 62.497 25.394 ;
      RECT MASK 2 62.749 22.0915 62.829 25.394 ;
      RECT MASK 2 65.217 22.0915 65.297 25.394 ;
      RECT MASK 2 65.549 22.0915 65.629 25.394 ;
      RECT MASK 2 65.881 22.0915 65.961 25.394 ;
      RECT MASK 2 66.379 22.0915 66.459 25.394 ;
      RECT MASK 2 66.711 22.0915 66.791 25.394 ;
      RECT MASK 2 67.043 22.0915 67.123 25.394 ;
      RECT MASK 2 67.541 22.0915 67.621 25.394 ;
      RECT MASK 2 67.873 22.0915 67.953 25.394 ;
      RECT MASK 2 68.205 22.0915 68.285 25.394 ;
      RECT MASK 2 68.703 22.0915 68.783 25.394 ;
      RECT MASK 2 69.035 22.0915 69.115 25.394 ;
      RECT MASK 2 69.367 22.0915 69.447 25.394 ;
      RECT MASK 2 71.835 22.0915 71.915 25.394 ;
      RECT MASK 2 72.167 22.0915 72.247 25.394 ;
      RECT MASK 2 72.499 22.0915 72.579 25.394 ;
      RECT MASK 2 72.997 22.0915 73.077 25.394 ;
      RECT MASK 2 73.329 22.0915 73.409 25.394 ;
      RECT MASK 2 73.661 22.0915 73.741 25.394 ;
      RECT MASK 2 74.159 22.0915 74.239 25.394 ;
      RECT MASK 2 74.491 22.0915 74.571 25.394 ;
      RECT MASK 2 74.823 22.0915 74.903 25.394 ;
      RECT MASK 2 75.321 22.0915 75.401 25.394 ;
      RECT MASK 2 75.653 22.0915 75.733 25.394 ;
      RECT MASK 2 75.985 22.0915 76.065 25.394 ;
      RECT MASK 2 78.453 22.0915 78.533 25.394 ;
      RECT MASK 2 78.785 22.0915 78.865 25.394 ;
      RECT MASK 2 79.117 22.0915 79.197 25.394 ;
      RECT MASK 2 79.615 22.0915 79.695 25.394 ;
      RECT MASK 2 79.947 22.0915 80.027 25.394 ;
      RECT MASK 2 80.279 22.0915 80.359 25.394 ;
      RECT MASK 2 80.777 22.0915 80.857 25.394 ;
      RECT MASK 2 81.109 22.0915 81.189 25.394 ;
      RECT MASK 2 81.441 22.0915 81.521 25.394 ;
      RECT MASK 2 81.939 22.0915 82.019 25.394 ;
      RECT MASK 2 82.271 22.0915 82.351 25.394 ;
      RECT MASK 2 82.603 22.0915 82.683 25.394 ;
      RECT MASK 2 85.071 22.0915 85.151 25.394 ;
      RECT MASK 2 85.403 22.0915 85.483 25.394 ;
      RECT MASK 2 85.735 22.0915 85.815 25.394 ;
      RECT MASK 2 86.233 22.0915 86.313 25.394 ;
      RECT MASK 2 86.565 22.0915 86.645 25.394 ;
      RECT MASK 2 86.897 22.0915 86.977 25.394 ;
      RECT MASK 2 87.395 22.0915 87.475 25.394 ;
      RECT MASK 2 87.727 22.0915 87.807 25.394 ;
      RECT MASK 2 88.059 22.0915 88.139 25.394 ;
      RECT MASK 2 88.557 22.0915 88.637 25.394 ;
      RECT MASK 2 88.889 22.0915 88.969 25.394 ;
      RECT MASK 2 89.221 22.0915 89.301 25.394 ;
      RECT MASK 2 91.689 22.0915 91.769 25.394 ;
      RECT MASK 2 92.021 22.0915 92.101 25.394 ;
      RECT MASK 2 92.353 22.0915 92.433 25.394 ;
      RECT MASK 2 92.851 22.0915 92.931 25.394 ;
      RECT MASK 2 93.183 22.0915 93.263 25.394 ;
      RECT MASK 2 93.515 22.0915 93.595 25.394 ;
      RECT MASK 2 94.013 22.0915 94.093 25.394 ;
      RECT MASK 2 94.345 22.0915 94.425 25.394 ;
      RECT MASK 2 94.677 22.0915 94.757 25.394 ;
      RECT MASK 2 95.175 22.0915 95.255 25.394 ;
      RECT MASK 2 95.507 22.0915 95.587 25.394 ;
      RECT MASK 2 95.839 22.0915 95.919 25.394 ;
      RECT MASK 2 98.307 22.0915 98.387 25.394 ;
      RECT MASK 2 98.639 22.0915 98.719 25.394 ;
      RECT MASK 2 98.971 22.0915 99.051 25.394 ;
      RECT MASK 2 99.469 22.0915 99.549 25.394 ;
      RECT MASK 2 99.801 22.0915 99.881 25.394 ;
      RECT MASK 2 100.133 22.0915 100.213 25.394 ;
      RECT MASK 2 100.631 22.0915 100.711 25.394 ;
      RECT MASK 2 100.963 22.0915 101.043 25.394 ;
      RECT MASK 2 101.295 22.0915 101.375 25.394 ;
      RECT MASK 2 101.793 22.0915 101.873 25.394 ;
      RECT MASK 2 102.125 22.0915 102.205 25.394 ;
      RECT MASK 2 102.457 22.0915 102.537 25.394 ;
      RECT MASK 2 104.925 22.0915 105.005 25.394 ;
      RECT MASK 2 105.257 22.0915 105.337 25.394 ;
      RECT MASK 2 105.589 22.0915 105.669 25.394 ;
      RECT MASK 2 106.087 22.0915 106.167 25.394 ;
      RECT MASK 2 106.419 22.0915 106.499 25.394 ;
      RECT MASK 2 106.751 22.0915 106.831 25.394 ;
      RECT MASK 2 107.249 22.0915 107.329 25.394 ;
      RECT MASK 2 107.581 22.0915 107.661 25.394 ;
      RECT MASK 2 107.913 22.0915 107.993 25.394 ;
      RECT MASK 2 108.411 22.0915 108.491 25.394 ;
      RECT MASK 2 108.743 22.0915 108.823 25.394 ;
      RECT MASK 2 109.075 22.0915 109.155 25.394 ;
      RECT MASK 2 5.499 23.28 5.559 23.55 ;
      RECT MASK 2 6.661 23.28 6.721 23.55 ;
      RECT MASK 2 7.823 23.28 7.883 23.55 ;
      RECT MASK 2 8.985 23.28 9.045 23.55 ;
      RECT MASK 2 10.147 23.28 10.207 23.55 ;
      RECT MASK 2 12.117 23.28 12.177 23.55 ;
      RECT MASK 2 13.279 23.28 13.339 23.55 ;
      RECT MASK 2 14.441 23.28 14.501 23.55 ;
      RECT MASK 2 15.603 23.28 15.663 23.55 ;
      RECT MASK 2 16.765 23.28 16.825 23.55 ;
      RECT MASK 2 18.735 23.28 18.795 23.55 ;
      RECT MASK 2 19.897 23.28 19.957 23.55 ;
      RECT MASK 2 21.059 23.28 21.119 23.55 ;
      RECT MASK 2 22.221 23.28 22.281 23.55 ;
      RECT MASK 2 23.383 23.28 23.443 23.55 ;
      RECT MASK 2 25.353 23.28 25.413 23.55 ;
      RECT MASK 2 26.515 23.28 26.575 23.55 ;
      RECT MASK 2 27.677 23.28 27.737 23.55 ;
      RECT MASK 2 28.839 23.28 28.899 23.55 ;
      RECT MASK 2 30.001 23.28 30.061 23.55 ;
      RECT MASK 2 31.971 23.28 32.031 23.55 ;
      RECT MASK 2 33.133 23.28 33.193 23.55 ;
      RECT MASK 2 34.295 23.28 34.355 23.55 ;
      RECT MASK 2 35.457 23.28 35.517 23.55 ;
      RECT MASK 2 36.619 23.28 36.679 23.55 ;
      RECT MASK 2 38.589 23.28 38.649 23.55 ;
      RECT MASK 2 39.751 23.28 39.811 23.55 ;
      RECT MASK 2 40.913 23.28 40.973 23.55 ;
      RECT MASK 2 42.075 23.28 42.135 23.55 ;
      RECT MASK 2 43.237 23.28 43.297 23.55 ;
      RECT MASK 2 45.207 23.28 45.267 23.55 ;
      RECT MASK 2 46.369 23.28 46.429 23.55 ;
      RECT MASK 2 47.531 23.28 47.591 23.55 ;
      RECT MASK 2 48.693 23.28 48.753 23.55 ;
      RECT MASK 2 49.855 23.28 49.915 23.55 ;
      RECT MASK 2 51.825 23.28 51.885 23.55 ;
      RECT MASK 2 52.987 23.28 53.047 23.55 ;
      RECT MASK 2 54.149 23.28 54.209 23.55 ;
      RECT MASK 2 55.311 23.28 55.371 23.55 ;
      RECT MASK 2 56.473 23.28 56.533 23.55 ;
      RECT MASK 2 58.443 23.28 58.503 23.55 ;
      RECT MASK 2 59.605 23.28 59.665 23.55 ;
      RECT MASK 2 60.767 23.28 60.827 23.55 ;
      RECT MASK 2 61.929 23.28 61.989 23.55 ;
      RECT MASK 2 63.091 23.28 63.151 23.55 ;
      RECT MASK 2 65.061 23.28 65.121 23.55 ;
      RECT MASK 2 66.223 23.28 66.283 23.55 ;
      RECT MASK 2 67.385 23.28 67.445 23.55 ;
      RECT MASK 2 68.547 23.28 68.607 23.55 ;
      RECT MASK 2 69.709 23.28 69.769 23.55 ;
      RECT MASK 2 71.679 23.28 71.739 23.55 ;
      RECT MASK 2 72.841 23.28 72.901 23.55 ;
      RECT MASK 2 74.003 23.28 74.063 23.55 ;
      RECT MASK 2 75.165 23.28 75.225 23.55 ;
      RECT MASK 2 76.327 23.28 76.387 23.55 ;
      RECT MASK 2 78.297 23.28 78.357 23.55 ;
      RECT MASK 2 79.459 23.28 79.519 23.55 ;
      RECT MASK 2 80.621 23.28 80.681 23.55 ;
      RECT MASK 2 81.783 23.28 81.843 23.55 ;
      RECT MASK 2 82.945 23.28 83.005 23.55 ;
      RECT MASK 2 84.915 23.28 84.975 23.55 ;
      RECT MASK 2 86.077 23.28 86.137 23.55 ;
      RECT MASK 2 87.239 23.28 87.299 23.55 ;
      RECT MASK 2 88.401 23.28 88.461 23.55 ;
      RECT MASK 2 89.563 23.28 89.623 23.55 ;
      RECT MASK 2 91.533 23.28 91.593 23.55 ;
      RECT MASK 2 92.695 23.28 92.755 23.55 ;
      RECT MASK 2 93.857 23.28 93.917 23.55 ;
      RECT MASK 2 95.019 23.28 95.079 23.55 ;
      RECT MASK 2 96.181 23.28 96.241 23.55 ;
      RECT MASK 2 98.151 23.28 98.211 23.55 ;
      RECT MASK 2 99.313 23.28 99.373 23.55 ;
      RECT MASK 2 100.475 23.28 100.535 23.55 ;
      RECT MASK 2 101.637 23.28 101.697 23.55 ;
      RECT MASK 2 102.799 23.28 102.859 23.55 ;
      RECT MASK 2 104.769 23.28 104.829 23.55 ;
      RECT MASK 2 105.931 23.28 105.991 23.55 ;
      RECT MASK 2 107.093 23.28 107.153 23.55 ;
      RECT MASK 2 108.255 23.28 108.315 23.55 ;
      RECT MASK 2 109.417 23.28 109.477 23.55 ;
      RECT MASK 2 5.499 23.73 5.559 24 ;
      RECT MASK 2 6.661 23.73 6.721 24 ;
      RECT MASK 2 7.823 23.73 7.883 24 ;
      RECT MASK 2 8.985 23.73 9.045 24 ;
      RECT MASK 2 10.147 23.73 10.207 24 ;
      RECT MASK 2 12.117 23.73 12.177 24 ;
      RECT MASK 2 13.279 23.73 13.339 24 ;
      RECT MASK 2 14.441 23.73 14.501 24 ;
      RECT MASK 2 15.603 23.73 15.663 24 ;
      RECT MASK 2 16.765 23.73 16.825 24 ;
      RECT MASK 2 18.735 23.73 18.795 24 ;
      RECT MASK 2 19.897 23.73 19.957 24 ;
      RECT MASK 2 21.059 23.73 21.119 24 ;
      RECT MASK 2 22.221 23.73 22.281 24 ;
      RECT MASK 2 23.383 23.73 23.443 24 ;
      RECT MASK 2 25.353 23.73 25.413 24 ;
      RECT MASK 2 26.515 23.73 26.575 24 ;
      RECT MASK 2 27.677 23.73 27.737 24 ;
      RECT MASK 2 28.839 23.73 28.899 24 ;
      RECT MASK 2 30.001 23.73 30.061 24 ;
      RECT MASK 2 31.971 23.73 32.031 24 ;
      RECT MASK 2 33.133 23.73 33.193 24 ;
      RECT MASK 2 34.295 23.73 34.355 24 ;
      RECT MASK 2 35.457 23.73 35.517 24 ;
      RECT MASK 2 36.619 23.73 36.679 24 ;
      RECT MASK 2 38.589 23.73 38.649 24 ;
      RECT MASK 2 39.751 23.73 39.811 24 ;
      RECT MASK 2 40.913 23.73 40.973 24 ;
      RECT MASK 2 42.075 23.73 42.135 24 ;
      RECT MASK 2 43.237 23.73 43.297 24 ;
      RECT MASK 2 45.207 23.73 45.267 24 ;
      RECT MASK 2 46.369 23.73 46.429 24 ;
      RECT MASK 2 47.531 23.73 47.591 24 ;
      RECT MASK 2 48.693 23.73 48.753 24 ;
      RECT MASK 2 49.855 23.73 49.915 24 ;
      RECT MASK 2 51.825 23.73 51.885 24 ;
      RECT MASK 2 52.987 23.73 53.047 24 ;
      RECT MASK 2 54.149 23.73 54.209 24 ;
      RECT MASK 2 55.311 23.73 55.371 24 ;
      RECT MASK 2 56.473 23.73 56.533 24 ;
      RECT MASK 2 58.443 23.73 58.503 24 ;
      RECT MASK 2 59.605 23.73 59.665 24 ;
      RECT MASK 2 60.767 23.73 60.827 24 ;
      RECT MASK 2 61.929 23.73 61.989 24 ;
      RECT MASK 2 63.091 23.73 63.151 24 ;
      RECT MASK 2 65.061 23.73 65.121 24 ;
      RECT MASK 2 66.223 23.73 66.283 24 ;
      RECT MASK 2 67.385 23.73 67.445 24 ;
      RECT MASK 2 68.547 23.73 68.607 24 ;
      RECT MASK 2 69.709 23.73 69.769 24 ;
      RECT MASK 2 71.679 23.73 71.739 24 ;
      RECT MASK 2 72.841 23.73 72.901 24 ;
      RECT MASK 2 74.003 23.73 74.063 24 ;
      RECT MASK 2 75.165 23.73 75.225 24 ;
      RECT MASK 2 76.327 23.73 76.387 24 ;
      RECT MASK 2 78.297 23.73 78.357 24 ;
      RECT MASK 2 79.459 23.73 79.519 24 ;
      RECT MASK 2 80.621 23.73 80.681 24 ;
      RECT MASK 2 81.783 23.73 81.843 24 ;
      RECT MASK 2 82.945 23.73 83.005 24 ;
      RECT MASK 2 84.915 23.73 84.975 24 ;
      RECT MASK 2 86.077 23.73 86.137 24 ;
      RECT MASK 2 87.239 23.73 87.299 24 ;
      RECT MASK 2 88.401 23.73 88.461 24 ;
      RECT MASK 2 89.563 23.73 89.623 24 ;
      RECT MASK 2 91.533 23.73 91.593 24 ;
      RECT MASK 2 92.695 23.73 92.755 24 ;
      RECT MASK 2 93.857 23.73 93.917 24 ;
      RECT MASK 2 95.019 23.73 95.079 24 ;
      RECT MASK 2 96.181 23.73 96.241 24 ;
      RECT MASK 2 98.151 23.73 98.211 24 ;
      RECT MASK 2 99.313 23.73 99.373 24 ;
      RECT MASK 2 100.475 23.73 100.535 24 ;
      RECT MASK 2 101.637 23.73 101.697 24 ;
      RECT MASK 2 102.799 23.73 102.859 24 ;
      RECT MASK 2 104.769 23.73 104.829 24 ;
      RECT MASK 2 105.931 23.73 105.991 24 ;
      RECT MASK 2 107.093 23.73 107.153 24 ;
      RECT MASK 2 108.255 23.73 108.315 24 ;
      RECT MASK 2 109.417 23.73 109.477 24 ;
      RECT MASK 2 5.499 25.68 5.559 25.95 ;
      RECT MASK 2 5.997 25.68 6.057 25.95 ;
      RECT MASK 2 6.329 25.68 6.389 25.95 ;
      RECT MASK 2 6.661 25.68 6.721 25.95 ;
      RECT MASK 2 7.159 25.68 7.219 25.95 ;
      RECT MASK 2 7.491 25.68 7.551 25.95 ;
      RECT MASK 2 7.823 25.68 7.883 25.95 ;
      RECT MASK 2 8.321 25.68 8.381 25.95 ;
      RECT MASK 2 8.653 25.68 8.713 25.95 ;
      RECT MASK 2 8.985 25.68 9.045 25.95 ;
      RECT MASK 2 9.483 25.68 9.543 25.95 ;
      RECT MASK 2 9.815 25.68 9.875 25.95 ;
      RECT MASK 2 10.147 25.68 10.207 25.95 ;
      RECT MASK 2 12.117 25.68 12.177 25.95 ;
      RECT MASK 2 12.615 25.68 12.675 25.95 ;
      RECT MASK 2 12.947 25.68 13.007 25.95 ;
      RECT MASK 2 13.279 25.68 13.339 25.95 ;
      RECT MASK 2 13.777 25.68 13.837 25.95 ;
      RECT MASK 2 14.109 25.68 14.169 25.95 ;
      RECT MASK 2 14.441 25.68 14.501 25.95 ;
      RECT MASK 2 14.939 25.68 14.999 25.95 ;
      RECT MASK 2 15.271 25.68 15.331 25.95 ;
      RECT MASK 2 15.603 25.68 15.663 25.95 ;
      RECT MASK 2 16.101 25.68 16.161 25.95 ;
      RECT MASK 2 16.433 25.68 16.493 25.95 ;
      RECT MASK 2 16.765 25.68 16.825 25.95 ;
      RECT MASK 2 18.735 25.68 18.795 25.95 ;
      RECT MASK 2 19.233 25.68 19.293 25.95 ;
      RECT MASK 2 19.565 25.68 19.625 25.95 ;
      RECT MASK 2 19.897 25.68 19.957 25.95 ;
      RECT MASK 2 20.395 25.68 20.455 25.95 ;
      RECT MASK 2 20.727 25.68 20.787 25.95 ;
      RECT MASK 2 21.059 25.68 21.119 25.95 ;
      RECT MASK 2 21.557 25.68 21.617 25.95 ;
      RECT MASK 2 21.889 25.68 21.949 25.95 ;
      RECT MASK 2 22.221 25.68 22.281 25.95 ;
      RECT MASK 2 22.719 25.68 22.779 25.95 ;
      RECT MASK 2 23.051 25.68 23.111 25.95 ;
      RECT MASK 2 23.383 25.68 23.443 25.95 ;
      RECT MASK 2 25.353 25.68 25.413 25.95 ;
      RECT MASK 2 25.851 25.68 25.911 25.95 ;
      RECT MASK 2 26.183 25.68 26.243 25.95 ;
      RECT MASK 2 26.515 25.68 26.575 25.95 ;
      RECT MASK 2 27.013 25.68 27.073 25.95 ;
      RECT MASK 2 27.345 25.68 27.405 25.95 ;
      RECT MASK 2 27.677 25.68 27.737 25.95 ;
      RECT MASK 2 28.175 25.68 28.235 25.95 ;
      RECT MASK 2 28.507 25.68 28.567 25.95 ;
      RECT MASK 2 28.839 25.68 28.899 25.95 ;
      RECT MASK 2 29.337 25.68 29.397 25.95 ;
      RECT MASK 2 29.669 25.68 29.729 25.95 ;
      RECT MASK 2 30.001 25.68 30.061 25.95 ;
      RECT MASK 2 31.971 25.68 32.031 25.95 ;
      RECT MASK 2 32.469 25.68 32.529 25.95 ;
      RECT MASK 2 32.801 25.68 32.861 25.95 ;
      RECT MASK 2 33.133 25.68 33.193 25.95 ;
      RECT MASK 2 33.631 25.68 33.691 25.95 ;
      RECT MASK 2 33.963 25.68 34.023 25.95 ;
      RECT MASK 2 34.295 25.68 34.355 25.95 ;
      RECT MASK 2 34.793 25.68 34.853 25.95 ;
      RECT MASK 2 35.125 25.68 35.185 25.95 ;
      RECT MASK 2 35.457 25.68 35.517 25.95 ;
      RECT MASK 2 35.955 25.68 36.015 25.95 ;
      RECT MASK 2 36.287 25.68 36.347 25.95 ;
      RECT MASK 2 36.619 25.68 36.679 25.95 ;
      RECT MASK 2 38.589 25.68 38.649 25.95 ;
      RECT MASK 2 39.087 25.68 39.147 25.95 ;
      RECT MASK 2 39.419 25.68 39.479 25.95 ;
      RECT MASK 2 39.751 25.68 39.811 25.95 ;
      RECT MASK 2 40.249 25.68 40.309 25.95 ;
      RECT MASK 2 40.581 25.68 40.641 25.95 ;
      RECT MASK 2 40.913 25.68 40.973 25.95 ;
      RECT MASK 2 41.411 25.68 41.471 25.95 ;
      RECT MASK 2 41.743 25.68 41.803 25.95 ;
      RECT MASK 2 42.075 25.68 42.135 25.95 ;
      RECT MASK 2 42.573 25.68 42.633 25.95 ;
      RECT MASK 2 42.905 25.68 42.965 25.95 ;
      RECT MASK 2 43.237 25.68 43.297 25.95 ;
      RECT MASK 2 45.207 25.68 45.267 25.95 ;
      RECT MASK 2 45.705 25.68 45.765 25.95 ;
      RECT MASK 2 46.037 25.68 46.097 25.95 ;
      RECT MASK 2 46.369 25.68 46.429 25.95 ;
      RECT MASK 2 46.867 25.68 46.927 25.95 ;
      RECT MASK 2 47.199 25.68 47.259 25.95 ;
      RECT MASK 2 47.531 25.68 47.591 25.95 ;
      RECT MASK 2 48.029 25.68 48.089 25.95 ;
      RECT MASK 2 48.361 25.68 48.421 25.95 ;
      RECT MASK 2 48.693 25.68 48.753 25.95 ;
      RECT MASK 2 49.191 25.68 49.251 25.95 ;
      RECT MASK 2 49.523 25.68 49.583 25.95 ;
      RECT MASK 2 49.855 25.68 49.915 25.95 ;
      RECT MASK 2 51.825 25.68 51.885 25.95 ;
      RECT MASK 2 52.323 25.68 52.383 25.95 ;
      RECT MASK 2 52.655 25.68 52.715 25.95 ;
      RECT MASK 2 52.987 25.68 53.047 25.95 ;
      RECT MASK 2 53.485 25.68 53.545 25.95 ;
      RECT MASK 2 53.817 25.68 53.877 25.95 ;
      RECT MASK 2 54.149 25.68 54.209 25.95 ;
      RECT MASK 2 54.647 25.68 54.707 25.95 ;
      RECT MASK 2 54.979 25.68 55.039 25.95 ;
      RECT MASK 2 55.311 25.68 55.371 25.95 ;
      RECT MASK 2 55.809 25.68 55.869 25.95 ;
      RECT MASK 2 56.141 25.68 56.201 25.95 ;
      RECT MASK 2 56.473 25.68 56.533 25.95 ;
      RECT MASK 2 58.443 25.68 58.503 25.95 ;
      RECT MASK 2 58.941 25.68 59.001 25.95 ;
      RECT MASK 2 59.273 25.68 59.333 25.95 ;
      RECT MASK 2 59.605 25.68 59.665 25.95 ;
      RECT MASK 2 60.103 25.68 60.163 25.95 ;
      RECT MASK 2 60.435 25.68 60.495 25.95 ;
      RECT MASK 2 60.767 25.68 60.827 25.95 ;
      RECT MASK 2 61.265 25.68 61.325 25.95 ;
      RECT MASK 2 61.597 25.68 61.657 25.95 ;
      RECT MASK 2 61.929 25.68 61.989 25.95 ;
      RECT MASK 2 62.427 25.68 62.487 25.95 ;
      RECT MASK 2 62.759 25.68 62.819 25.95 ;
      RECT MASK 2 63.091 25.68 63.151 25.95 ;
      RECT MASK 2 65.061 25.68 65.121 25.95 ;
      RECT MASK 2 65.559 25.68 65.619 25.95 ;
      RECT MASK 2 65.891 25.68 65.951 25.95 ;
      RECT MASK 2 66.223 25.68 66.283 25.95 ;
      RECT MASK 2 66.721 25.68 66.781 25.95 ;
      RECT MASK 2 67.053 25.68 67.113 25.95 ;
      RECT MASK 2 67.385 25.68 67.445 25.95 ;
      RECT MASK 2 67.883 25.68 67.943 25.95 ;
      RECT MASK 2 68.215 25.68 68.275 25.95 ;
      RECT MASK 2 68.547 25.68 68.607 25.95 ;
      RECT MASK 2 69.045 25.68 69.105 25.95 ;
      RECT MASK 2 69.377 25.68 69.437 25.95 ;
      RECT MASK 2 69.709 25.68 69.769 25.95 ;
      RECT MASK 2 71.679 25.68 71.739 25.95 ;
      RECT MASK 2 72.177 25.68 72.237 25.95 ;
      RECT MASK 2 72.509 25.68 72.569 25.95 ;
      RECT MASK 2 72.841 25.68 72.901 25.95 ;
      RECT MASK 2 73.339 25.68 73.399 25.95 ;
      RECT MASK 2 73.671 25.68 73.731 25.95 ;
      RECT MASK 2 74.003 25.68 74.063 25.95 ;
      RECT MASK 2 74.501 25.68 74.561 25.95 ;
      RECT MASK 2 74.833 25.68 74.893 25.95 ;
      RECT MASK 2 75.165 25.68 75.225 25.95 ;
      RECT MASK 2 75.663 25.68 75.723 25.95 ;
      RECT MASK 2 75.995 25.68 76.055 25.95 ;
      RECT MASK 2 76.327 25.68 76.387 25.95 ;
      RECT MASK 2 78.297 25.68 78.357 25.95 ;
      RECT MASK 2 78.795 25.68 78.855 25.95 ;
      RECT MASK 2 79.127 25.68 79.187 25.95 ;
      RECT MASK 2 79.459 25.68 79.519 25.95 ;
      RECT MASK 2 79.957 25.68 80.017 25.95 ;
      RECT MASK 2 80.289 25.68 80.349 25.95 ;
      RECT MASK 2 80.621 25.68 80.681 25.95 ;
      RECT MASK 2 81.119 25.68 81.179 25.95 ;
      RECT MASK 2 81.451 25.68 81.511 25.95 ;
      RECT MASK 2 81.783 25.68 81.843 25.95 ;
      RECT MASK 2 82.281 25.68 82.341 25.95 ;
      RECT MASK 2 82.613 25.68 82.673 25.95 ;
      RECT MASK 2 82.945 25.68 83.005 25.95 ;
      RECT MASK 2 84.915 25.68 84.975 25.95 ;
      RECT MASK 2 85.413 25.68 85.473 25.95 ;
      RECT MASK 2 85.745 25.68 85.805 25.95 ;
      RECT MASK 2 86.077 25.68 86.137 25.95 ;
      RECT MASK 2 86.575 25.68 86.635 25.95 ;
      RECT MASK 2 86.907 25.68 86.967 25.95 ;
      RECT MASK 2 87.239 25.68 87.299 25.95 ;
      RECT MASK 2 87.737 25.68 87.797 25.95 ;
      RECT MASK 2 88.069 25.68 88.129 25.95 ;
      RECT MASK 2 88.401 25.68 88.461 25.95 ;
      RECT MASK 2 88.899 25.68 88.959 25.95 ;
      RECT MASK 2 89.231 25.68 89.291 25.95 ;
      RECT MASK 2 89.563 25.68 89.623 25.95 ;
      RECT MASK 2 91.533 25.68 91.593 25.95 ;
      RECT MASK 2 92.031 25.68 92.091 25.95 ;
      RECT MASK 2 92.363 25.68 92.423 25.95 ;
      RECT MASK 2 92.695 25.68 92.755 25.95 ;
      RECT MASK 2 93.193 25.68 93.253 25.95 ;
      RECT MASK 2 93.525 25.68 93.585 25.95 ;
      RECT MASK 2 93.857 25.68 93.917 25.95 ;
      RECT MASK 2 94.355 25.68 94.415 25.95 ;
      RECT MASK 2 94.687 25.68 94.747 25.95 ;
      RECT MASK 2 95.019 25.68 95.079 25.95 ;
      RECT MASK 2 95.517 25.68 95.577 25.95 ;
      RECT MASK 2 95.849 25.68 95.909 25.95 ;
      RECT MASK 2 96.181 25.68 96.241 25.95 ;
      RECT MASK 2 98.151 25.68 98.211 25.95 ;
      RECT MASK 2 98.649 25.68 98.709 25.95 ;
      RECT MASK 2 98.981 25.68 99.041 25.95 ;
      RECT MASK 2 99.313 25.68 99.373 25.95 ;
      RECT MASK 2 99.811 25.68 99.871 25.95 ;
      RECT MASK 2 100.143 25.68 100.203 25.95 ;
      RECT MASK 2 100.475 25.68 100.535 25.95 ;
      RECT MASK 2 100.973 25.68 101.033 25.95 ;
      RECT MASK 2 101.305 25.68 101.365 25.95 ;
      RECT MASK 2 101.637 25.68 101.697 25.95 ;
      RECT MASK 2 102.135 25.68 102.195 25.95 ;
      RECT MASK 2 102.467 25.68 102.527 25.95 ;
      RECT MASK 2 102.799 25.68 102.859 25.95 ;
      RECT MASK 2 104.769 25.68 104.829 25.95 ;
      RECT MASK 2 105.267 25.68 105.327 25.95 ;
      RECT MASK 2 105.599 25.68 105.659 25.95 ;
      RECT MASK 2 105.931 25.68 105.991 25.95 ;
      RECT MASK 2 106.429 25.68 106.489 25.95 ;
      RECT MASK 2 106.761 25.68 106.821 25.95 ;
      RECT MASK 2 107.093 25.68 107.153 25.95 ;
      RECT MASK 2 107.591 25.68 107.651 25.95 ;
      RECT MASK 2 107.923 25.68 107.983 25.95 ;
      RECT MASK 2 108.255 25.68 108.315 25.95 ;
      RECT MASK 2 108.753 25.68 108.813 25.95 ;
      RECT MASK 2 109.085 25.68 109.145 25.95 ;
      RECT MASK 2 109.417 25.68 109.477 25.95 ;
      RECT MASK 2 2.929 26.1 3.229 77.8205 ;
      RECT MASK 2 1.839 26.156 1.919 26.476 ;
      RECT MASK 2 2.171 26.156 2.251 26.476 ;
      RECT MASK 2 2.503 26.156 2.583 26.476 ;
      RECT MASK 2 4.163 26.156 4.243 26.476 ;
      RECT MASK 2 4.495 26.156 4.575 26.476 ;
      RECT MASK 2 4.827 26.156 4.907 26.476 ;
      RECT MASK 2 5.159 26.156 5.239 26.476 ;
      RECT MASK 2 5.491 26.156 5.571 26.476 ;
      RECT MASK 2 5.823 26.156 5.903 26.476 ;
      RECT MASK 2 6.155 26.156 6.235 26.476 ;
      RECT MASK 2 6.487 26.156 6.567 26.476 ;
      RECT MASK 2 6.819 26.156 6.899 26.476 ;
      RECT MASK 2 7.151 26.156 7.231 26.476 ;
      RECT MASK 2 7.483 26.156 7.563 26.476 ;
      RECT MASK 2 7.815 26.156 7.895 26.476 ;
      RECT MASK 2 8.147 26.156 8.227 26.476 ;
      RECT MASK 2 8.479 26.156 8.559 26.476 ;
      RECT MASK 2 8.811 26.156 8.891 26.476 ;
      RECT MASK 2 9.143 26.156 9.223 26.476 ;
      RECT MASK 2 9.475 26.156 9.555 26.476 ;
      RECT MASK 2 9.807 26.156 9.887 26.476 ;
      RECT MASK 2 10.139 26.156 10.219 26.476 ;
      RECT MASK 2 10.471 26.156 10.551 26.476 ;
      RECT MASK 2 10.803 26.156 10.883 26.476 ;
      RECT MASK 2 11.135 26.156 11.215 26.476 ;
      RECT MASK 2 11.467 26.156 11.547 26.476 ;
      RECT MASK 2 11.799 26.156 11.879 26.476 ;
      RECT MASK 2 12.131 26.156 12.211 26.476 ;
      RECT MASK 2 12.463 26.156 12.543 26.476 ;
      RECT MASK 2 12.795 26.156 12.875 26.476 ;
      RECT MASK 2 13.127 26.156 13.207 26.476 ;
      RECT MASK 2 13.459 26.156 13.539 26.476 ;
      RECT MASK 2 13.791 26.156 13.871 26.476 ;
      RECT MASK 2 14.123 26.156 14.203 26.476 ;
      RECT MASK 2 14.455 26.156 14.535 26.476 ;
      RECT MASK 2 14.787 26.156 14.867 26.476 ;
      RECT MASK 2 15.119 26.156 15.199 26.476 ;
      RECT MASK 2 15.451 26.156 15.531 26.476 ;
      RECT MASK 2 15.783 26.156 15.863 26.476 ;
      RECT MASK 2 16.115 26.156 16.195 26.476 ;
      RECT MASK 2 16.447 26.156 16.527 26.476 ;
      RECT MASK 2 16.779 26.156 16.859 26.476 ;
      RECT MASK 2 17.111 26.156 17.191 26.476 ;
      RECT MASK 2 17.443 26.156 17.523 26.476 ;
      RECT MASK 2 17.775 26.156 17.855 26.476 ;
      RECT MASK 2 18.107 26.156 18.187 26.476 ;
      RECT MASK 2 18.439 26.156 18.519 26.476 ;
      RECT MASK 2 18.771 26.156 18.851 26.476 ;
      RECT MASK 2 19.103 26.156 19.183 26.476 ;
      RECT MASK 2 19.435 26.156 19.515 26.476 ;
      RECT MASK 2 19.767 26.156 19.847 26.476 ;
      RECT MASK 2 20.099 26.156 20.179 26.476 ;
      RECT MASK 2 20.431 26.156 20.511 26.476 ;
      RECT MASK 2 20.763 26.156 20.843 26.476 ;
      RECT MASK 2 21.095 26.156 21.175 26.476 ;
      RECT MASK 2 21.427 26.156 21.507 26.476 ;
      RECT MASK 2 21.759 26.156 21.839 26.476 ;
      RECT MASK 2 22.091 26.156 22.171 26.476 ;
      RECT MASK 2 22.423 26.156 22.503 26.476 ;
      RECT MASK 2 22.755 26.156 22.835 26.476 ;
      RECT MASK 2 23.087 26.156 23.167 26.476 ;
      RECT MASK 2 23.419 26.156 23.499 26.476 ;
      RECT MASK 2 23.751 26.156 23.831 26.476 ;
      RECT MASK 2 24.083 26.156 24.163 26.476 ;
      RECT MASK 2 24.415 26.156 24.495 26.476 ;
      RECT MASK 2 24.747 26.156 24.827 26.476 ;
      RECT MASK 2 25.079 26.156 25.159 26.476 ;
      RECT MASK 2 25.411 26.156 25.491 26.476 ;
      RECT MASK 2 25.743 26.156 25.823 26.476 ;
      RECT MASK 2 26.075 26.156 26.155 26.476 ;
      RECT MASK 2 26.407 26.156 26.487 26.476 ;
      RECT MASK 2 26.739 26.156 26.819 26.476 ;
      RECT MASK 2 27.071 26.156 27.151 26.476 ;
      RECT MASK 2 27.403 26.156 27.483 26.476 ;
      RECT MASK 2 27.735 26.156 27.815 26.476 ;
      RECT MASK 2 28.067 26.156 28.147 26.476 ;
      RECT MASK 2 28.399 26.156 28.479 26.476 ;
      RECT MASK 2 28.731 26.156 28.811 26.476 ;
      RECT MASK 2 29.063 26.156 29.143 26.476 ;
      RECT MASK 2 29.395 26.156 29.475 26.476 ;
      RECT MASK 2 29.727 26.156 29.807 26.476 ;
      RECT MASK 2 30.059 26.156 30.139 26.476 ;
      RECT MASK 2 30.391 26.156 30.471 26.476 ;
      RECT MASK 2 30.723 26.156 30.803 26.476 ;
      RECT MASK 2 31.055 26.156 31.135 26.476 ;
      RECT MASK 2 31.387 26.156 31.467 26.476 ;
      RECT MASK 2 31.719 26.156 31.799 26.476 ;
      RECT MASK 2 32.051 26.156 32.131 26.476 ;
      RECT MASK 2 32.383 26.156 32.463 26.476 ;
      RECT MASK 2 32.715 26.156 32.795 26.476 ;
      RECT MASK 2 33.047 26.156 33.127 26.476 ;
      RECT MASK 2 33.379 26.156 33.459 26.476 ;
      RECT MASK 2 33.711 26.156 33.791 26.476 ;
      RECT MASK 2 34.043 26.156 34.123 26.476 ;
      RECT MASK 2 34.375 26.156 34.455 26.476 ;
      RECT MASK 2 34.707 26.156 34.787 26.476 ;
      RECT MASK 2 35.039 26.156 35.119 26.476 ;
      RECT MASK 2 35.371 26.156 35.451 26.476 ;
      RECT MASK 2 35.703 26.156 35.783 26.476 ;
      RECT MASK 2 36.035 26.156 36.115 26.476 ;
      RECT MASK 2 36.367 26.156 36.447 26.476 ;
      RECT MASK 2 36.699 26.156 36.779 26.476 ;
      RECT MASK 2 37.031 26.156 37.111 26.476 ;
      RECT MASK 2 37.363 26.156 37.443 26.476 ;
      RECT MASK 2 37.695 26.156 37.775 26.476 ;
      RECT MASK 2 38.027 26.156 38.107 26.476 ;
      RECT MASK 2 38.359 26.156 38.439 26.476 ;
      RECT MASK 2 38.691 26.156 38.771 26.476 ;
      RECT MASK 2 39.023 26.156 39.103 26.476 ;
      RECT MASK 2 39.355 26.156 39.435 26.476 ;
      RECT MASK 2 39.687 26.156 39.767 26.476 ;
      RECT MASK 2 40.019 26.156 40.099 26.476 ;
      RECT MASK 2 40.351 26.156 40.431 26.476 ;
      RECT MASK 2 40.683 26.156 40.763 26.476 ;
      RECT MASK 2 41.015 26.156 41.095 26.476 ;
      RECT MASK 2 41.347 26.156 41.427 26.476 ;
      RECT MASK 2 41.679 26.156 41.759 26.476 ;
      RECT MASK 2 42.011 26.156 42.091 26.476 ;
      RECT MASK 2 42.343 26.156 42.423 26.476 ;
      RECT MASK 2 42.675 26.156 42.755 26.476 ;
      RECT MASK 2 43.007 26.156 43.087 26.476 ;
      RECT MASK 2 43.339 26.156 43.419 26.476 ;
      RECT MASK 2 43.671 26.156 43.751 26.476 ;
      RECT MASK 2 44.003 26.156 44.083 26.476 ;
      RECT MASK 2 44.335 26.156 44.415 26.476 ;
      RECT MASK 2 44.667 26.156 44.747 26.476 ;
      RECT MASK 2 44.999 26.156 45.079 26.476 ;
      RECT MASK 2 45.331 26.156 45.411 26.476 ;
      RECT MASK 2 45.663 26.156 45.743 26.476 ;
      RECT MASK 2 45.995 26.156 46.075 26.476 ;
      RECT MASK 2 46.327 26.156 46.407 26.476 ;
      RECT MASK 2 46.659 26.156 46.739 26.476 ;
      RECT MASK 2 46.991 26.156 47.071 26.476 ;
      RECT MASK 2 47.323 26.156 47.403 26.476 ;
      RECT MASK 2 47.655 26.156 47.735 26.476 ;
      RECT MASK 2 47.987 26.156 48.067 26.476 ;
      RECT MASK 2 48.319 26.156 48.399 26.476 ;
      RECT MASK 2 48.651 26.156 48.731 26.476 ;
      RECT MASK 2 48.983 26.156 49.063 26.476 ;
      RECT MASK 2 49.315 26.156 49.395 26.476 ;
      RECT MASK 2 49.647 26.156 49.727 26.476 ;
      RECT MASK 2 49.979 26.156 50.059 26.476 ;
      RECT MASK 2 50.311 26.156 50.391 26.476 ;
      RECT MASK 2 50.643 26.156 50.723 26.476 ;
      RECT MASK 2 50.975 26.156 51.055 26.476 ;
      RECT MASK 2 51.307 26.156 51.387 26.476 ;
      RECT MASK 2 51.639 26.156 51.719 26.476 ;
      RECT MASK 2 51.971 26.156 52.051 26.476 ;
      RECT MASK 2 52.303 26.156 52.383 26.476 ;
      RECT MASK 2 52.635 26.156 52.715 26.476 ;
      RECT MASK 2 52.967 26.156 53.047 26.476 ;
      RECT MASK 2 53.299 26.156 53.379 26.476 ;
      RECT MASK 2 53.631 26.156 53.711 26.476 ;
      RECT MASK 2 53.963 26.156 54.043 26.476 ;
      RECT MASK 2 54.295 26.156 54.375 26.476 ;
      RECT MASK 2 54.627 26.156 54.707 26.476 ;
      RECT MASK 2 54.959 26.156 55.039 26.476 ;
      RECT MASK 2 55.291 26.156 55.371 26.476 ;
      RECT MASK 2 55.623 26.156 55.703 26.476 ;
      RECT MASK 2 55.955 26.156 56.035 26.476 ;
      RECT MASK 2 56.287 26.156 56.367 26.476 ;
      RECT MASK 2 56.619 26.156 56.699 26.476 ;
      RECT MASK 2 56.951 26.156 57.031 26.476 ;
      RECT MASK 2 57.283 26.156 57.363 26.476 ;
      RECT MASK 2 57.615 26.156 57.695 26.476 ;
      RECT MASK 2 57.947 26.156 58.027 26.476 ;
      RECT MASK 2 58.279 26.156 58.359 26.476 ;
      RECT MASK 2 58.611 26.156 58.691 26.476 ;
      RECT MASK 2 58.943 26.156 59.023 26.476 ;
      RECT MASK 2 59.275 26.156 59.355 26.476 ;
      RECT MASK 2 59.607 26.156 59.687 26.476 ;
      RECT MASK 2 59.939 26.156 60.019 26.476 ;
      RECT MASK 2 60.271 26.156 60.351 26.476 ;
      RECT MASK 2 60.603 26.156 60.683 26.476 ;
      RECT MASK 2 60.935 26.156 61.015 26.476 ;
      RECT MASK 2 61.267 26.156 61.347 26.476 ;
      RECT MASK 2 61.599 26.156 61.679 26.476 ;
      RECT MASK 2 61.931 26.156 62.011 26.476 ;
      RECT MASK 2 62.263 26.156 62.343 26.476 ;
      RECT MASK 2 62.595 26.156 62.675 26.476 ;
      RECT MASK 2 62.927 26.156 63.007 26.476 ;
      RECT MASK 2 63.259 26.156 63.339 26.476 ;
      RECT MASK 2 63.591 26.156 63.671 26.476 ;
      RECT MASK 2 63.923 26.156 64.003 26.476 ;
      RECT MASK 2 64.255 26.156 64.335 26.476 ;
      RECT MASK 2 64.587 26.156 64.667 26.476 ;
      RECT MASK 2 64.919 26.156 64.999 26.476 ;
      RECT MASK 2 65.251 26.156 65.331 26.476 ;
      RECT MASK 2 65.583 26.156 65.663 26.476 ;
      RECT MASK 2 65.915 26.156 65.995 26.476 ;
      RECT MASK 2 66.247 26.156 66.327 26.476 ;
      RECT MASK 2 66.579 26.156 66.659 26.476 ;
      RECT MASK 2 66.911 26.156 66.991 26.476 ;
      RECT MASK 2 67.243 26.156 67.323 26.476 ;
      RECT MASK 2 67.575 26.156 67.655 26.476 ;
      RECT MASK 2 67.907 26.156 67.987 26.476 ;
      RECT MASK 2 68.239 26.156 68.319 26.476 ;
      RECT MASK 2 68.571 26.156 68.651 26.476 ;
      RECT MASK 2 68.903 26.156 68.983 26.476 ;
      RECT MASK 2 69.235 26.156 69.315 26.476 ;
      RECT MASK 2 69.567 26.156 69.647 26.476 ;
      RECT MASK 2 69.899 26.156 69.979 26.476 ;
      RECT MASK 2 70.231 26.156 70.311 26.476 ;
      RECT MASK 2 70.563 26.156 70.643 26.476 ;
      RECT MASK 2 70.895 26.156 70.975 26.476 ;
      RECT MASK 2 71.227 26.156 71.307 26.476 ;
      RECT MASK 2 71.559 26.156 71.639 26.476 ;
      RECT MASK 2 71.891 26.156 71.971 26.476 ;
      RECT MASK 2 72.223 26.156 72.303 26.476 ;
      RECT MASK 2 72.555 26.156 72.635 26.476 ;
      RECT MASK 2 72.887 26.156 72.967 26.476 ;
      RECT MASK 2 73.219 26.156 73.299 26.476 ;
      RECT MASK 2 73.551 26.156 73.631 26.476 ;
      RECT MASK 2 73.883 26.156 73.963 26.476 ;
      RECT MASK 2 74.215 26.156 74.295 26.476 ;
      RECT MASK 2 74.547 26.156 74.627 26.476 ;
      RECT MASK 2 74.879 26.156 74.959 26.476 ;
      RECT MASK 2 75.211 26.156 75.291 26.476 ;
      RECT MASK 2 75.543 26.156 75.623 26.476 ;
      RECT MASK 2 75.875 26.156 75.955 26.476 ;
      RECT MASK 2 76.207 26.156 76.287 26.476 ;
      RECT MASK 2 76.539 26.156 76.619 26.476 ;
      RECT MASK 2 76.871 26.156 76.951 26.476 ;
      RECT MASK 2 77.203 26.156 77.283 26.476 ;
      RECT MASK 2 77.535 26.156 77.615 26.476 ;
      RECT MASK 2 77.867 26.156 77.947 26.476 ;
      RECT MASK 2 78.199 26.156 78.279 26.476 ;
      RECT MASK 2 78.531 26.156 78.611 26.476 ;
      RECT MASK 2 78.863 26.156 78.943 26.476 ;
      RECT MASK 2 79.195 26.156 79.275 26.476 ;
      RECT MASK 2 79.527 26.156 79.607 26.476 ;
      RECT MASK 2 79.859 26.156 79.939 26.476 ;
      RECT MASK 2 80.191 26.156 80.271 26.476 ;
      RECT MASK 2 80.523 26.156 80.603 26.476 ;
      RECT MASK 2 80.855 26.156 80.935 26.476 ;
      RECT MASK 2 81.187 26.156 81.267 26.476 ;
      RECT MASK 2 81.519 26.156 81.599 26.476 ;
      RECT MASK 2 81.851 26.156 81.931 26.476 ;
      RECT MASK 2 82.183 26.156 82.263 26.476 ;
      RECT MASK 2 82.515 26.156 82.595 26.476 ;
      RECT MASK 2 82.847 26.156 82.927 26.476 ;
      RECT MASK 2 83.179 26.156 83.259 26.476 ;
      RECT MASK 2 83.511 26.156 83.591 26.476 ;
      RECT MASK 2 83.843 26.156 83.923 26.476 ;
      RECT MASK 2 84.175 26.156 84.255 26.476 ;
      RECT MASK 2 84.507 26.156 84.587 26.476 ;
      RECT MASK 2 84.839 26.156 84.919 26.476 ;
      RECT MASK 2 85.171 26.156 85.251 26.476 ;
      RECT MASK 2 85.503 26.156 85.583 26.476 ;
      RECT MASK 2 85.835 26.156 85.915 26.476 ;
      RECT MASK 2 86.167 26.156 86.247 26.476 ;
      RECT MASK 2 86.499 26.156 86.579 26.476 ;
      RECT MASK 2 86.831 26.156 86.911 26.476 ;
      RECT MASK 2 87.163 26.156 87.243 26.476 ;
      RECT MASK 2 87.495 26.156 87.575 26.476 ;
      RECT MASK 2 87.827 26.156 87.907 26.476 ;
      RECT MASK 2 88.159 26.156 88.239 26.476 ;
      RECT MASK 2 88.491 26.156 88.571 26.476 ;
      RECT MASK 2 88.823 26.156 88.903 26.476 ;
      RECT MASK 2 89.155 26.156 89.235 26.476 ;
      RECT MASK 2 89.487 26.156 89.567 26.476 ;
      RECT MASK 2 89.819 26.156 89.899 26.476 ;
      RECT MASK 2 90.151 26.156 90.231 26.476 ;
      RECT MASK 2 90.483 26.156 90.563 26.476 ;
      RECT MASK 2 90.815 26.156 90.895 26.476 ;
      RECT MASK 2 91.147 26.156 91.227 26.476 ;
      RECT MASK 2 91.479 26.156 91.559 26.476 ;
      RECT MASK 2 91.811 26.156 91.891 26.476 ;
      RECT MASK 2 92.143 26.156 92.223 26.476 ;
      RECT MASK 2 92.475 26.156 92.555 26.476 ;
      RECT MASK 2 92.807 26.156 92.887 26.476 ;
      RECT MASK 2 93.139 26.156 93.219 26.476 ;
      RECT MASK 2 93.471 26.156 93.551 26.476 ;
      RECT MASK 2 93.803 26.156 93.883 26.476 ;
      RECT MASK 2 94.135 26.156 94.215 26.476 ;
      RECT MASK 2 94.467 26.156 94.547 26.476 ;
      RECT MASK 2 94.799 26.156 94.879 26.476 ;
      RECT MASK 2 95.131 26.156 95.211 26.476 ;
      RECT MASK 2 95.463 26.156 95.543 26.476 ;
      RECT MASK 2 95.795 26.156 95.875 26.476 ;
      RECT MASK 2 96.127 26.156 96.207 26.476 ;
      RECT MASK 2 96.459 26.156 96.539 26.476 ;
      RECT MASK 2 96.791 26.156 96.871 26.476 ;
      RECT MASK 2 97.123 26.156 97.203 26.476 ;
      RECT MASK 2 97.455 26.156 97.535 26.476 ;
      RECT MASK 2 97.787 26.156 97.867 26.476 ;
      RECT MASK 2 98.119 26.156 98.199 26.476 ;
      RECT MASK 2 98.451 26.156 98.531 26.476 ;
      RECT MASK 2 98.783 26.156 98.863 26.476 ;
      RECT MASK 2 99.115 26.156 99.195 26.476 ;
      RECT MASK 2 99.447 26.156 99.527 26.476 ;
      RECT MASK 2 99.779 26.156 99.859 26.476 ;
      RECT MASK 2 100.111 26.156 100.191 26.476 ;
      RECT MASK 2 100.443 26.156 100.523 26.476 ;
      RECT MASK 2 100.775 26.156 100.855 26.476 ;
      RECT MASK 2 101.107 26.156 101.187 26.476 ;
      RECT MASK 2 101.439 26.156 101.519 26.476 ;
      RECT MASK 2 101.771 26.156 101.851 26.476 ;
      RECT MASK 2 102.103 26.156 102.183 26.476 ;
      RECT MASK 2 102.435 26.156 102.515 26.476 ;
      RECT MASK 2 102.767 26.156 102.847 26.476 ;
      RECT MASK 2 103.099 26.156 103.179 26.476 ;
      RECT MASK 2 103.431 26.156 103.511 26.476 ;
      RECT MASK 2 103.763 26.156 103.843 26.476 ;
      RECT MASK 2 104.095 26.156 104.175 26.476 ;
      RECT MASK 2 104.427 26.156 104.507 26.476 ;
      RECT MASK 2 104.759 26.156 104.839 26.476 ;
      RECT MASK 2 105.091 26.156 105.171 26.476 ;
      RECT MASK 2 105.423 26.156 105.503 26.476 ;
      RECT MASK 2 105.755 26.156 105.835 26.476 ;
      RECT MASK 2 106.087 26.156 106.167 26.476 ;
      RECT MASK 2 106.419 26.156 106.499 26.476 ;
      RECT MASK 2 106.751 26.156 106.831 26.476 ;
      RECT MASK 2 107.083 26.156 107.163 26.476 ;
      RECT MASK 2 107.415 26.156 107.495 26.476 ;
      RECT MASK 2 107.747 26.156 107.827 26.476 ;
      RECT MASK 2 108.079 26.156 108.159 26.476 ;
      RECT MASK 2 108.411 26.156 108.491 26.476 ;
      RECT MASK 2 108.743 26.156 108.823 26.476 ;
      RECT MASK 2 109.075 26.156 109.155 26.476 ;
      RECT MASK 2 109.407 26.156 109.487 26.476 ;
      RECT MASK 2 109.739 26.156 109.819 26.476 ;
      RECT MASK 2 110.071 26.156 110.151 26.476 ;
      RECT MASK 2 110.403 26.156 110.483 26.476 ;
      RECT MASK 2 110.735 26.156 110.815 26.476 ;
      RECT MASK 2 111.067 26.156 111.147 77.818 ;
      RECT MASK 2 111.399 26.156 111.479 77.818 ;
      RECT MASK 2 111.731 26.156 111.811 77.818 ;
      RECT MASK 2 112.063 26.156 112.143 77.818 ;
      RECT MASK 2 112.395 26.156 112.475 26.476 ;
      RECT MASK 2 112.727 26.156 112.807 26.476 ;
      RECT MASK 2 113.059 26.156 113.139 26.476 ;
      RECT MASK 2 113.391 26.156 113.471 26.476 ;
      RECT MASK 2 0.669 26.173 0.789 77.818 ;
      RECT MASK 2 1.321 26.173 1.441 77.818 ;
      RECT MASK 2 116.095 26.426 116.175 30.51 ;
      RECT MASK 2 116.427 26.426 116.507 26.728 ;
      RECT MASK 2 116.759 26.426 116.839 26.728 ;
      RECT MASK 2 117.091 26.426 117.171 26.728 ;
      RECT MASK 2 117.423 26.426 117.503 26.728 ;
      RECT MASK 2 117.755 26.426 117.835 26.728 ;
      RECT MASK 2 118.087 26.426 118.167 26.728 ;
      RECT MASK 2 118.419 26.426 118.499 26.728 ;
      RECT MASK 2 118.751 26.426 118.831 26.728 ;
      RECT MASK 2 119.083 26.426 119.163 26.728 ;
      RECT MASK 2 119.415 26.426 119.495 26.728 ;
      RECT MASK 2 119.747 26.426 119.827 26.728 ;
      RECT MASK 2 120.079 26.426 120.159 26.728 ;
      RECT MASK 2 120.411 26.426 120.491 26.728 ;
      RECT MASK 2 120.743 26.426 120.823 26.728 ;
      RECT MASK 2 121.075 26.426 121.155 26.728 ;
      RECT MASK 2 121.407 26.426 121.487 26.728 ;
      RECT MASK 2 121.739 26.426 121.819 26.728 ;
      RECT MASK 2 122.071 26.426 122.151 26.728 ;
      RECT MASK 2 122.403 26.426 122.483 26.728 ;
      RECT MASK 2 122.735 26.426 122.815 26.728 ;
      RECT MASK 2 123.067 26.426 123.147 26.728 ;
      RECT MASK 2 123.399 26.426 123.479 26.728 ;
      RECT MASK 2 123.731 26.426 123.811 26.728 ;
      RECT MASK 2 124.063 26.426 124.143 26.728 ;
      RECT MASK 2 124.395 26.426 124.475 26.728 ;
      RECT MASK 2 124.727 26.426 124.807 26.728 ;
      RECT MASK 2 125.059 26.426 125.139 26.728 ;
      RECT MASK 2 125.391 26.426 125.471 26.728 ;
      RECT MASK 2 125.723 26.426 125.803 26.728 ;
      RECT MASK 2 126.055 26.426 126.135 26.728 ;
      RECT MASK 2 126.387 26.426 126.467 30.51 ;
      RECT MASK 2 126.577 26.86 126.657 27.232 ;
      RECT MASK 2 116.427 26.94 116.507 29.758 ;
      RECT MASK 2 116.759 26.94 116.839 29.758 ;
      RECT MASK 2 117.091 26.94 117.171 29.758 ;
      RECT MASK 2 117.423 26.94 117.503 29.758 ;
      RECT MASK 2 117.755 26.94 117.835 29.758 ;
      RECT MASK 2 118.087 26.94 118.167 29.758 ;
      RECT MASK 2 118.419 26.94 118.499 29.758 ;
      RECT MASK 2 118.751 26.94 118.831 29.758 ;
      RECT MASK 2 119.083 26.94 119.163 29.758 ;
      RECT MASK 2 119.415 26.94 119.495 29.758 ;
      RECT MASK 2 119.747 26.94 119.827 29.758 ;
      RECT MASK 2 120.079 26.94 120.159 29.758 ;
      RECT MASK 2 120.411 26.94 120.491 29.758 ;
      RECT MASK 2 120.743 26.94 120.823 29.758 ;
      RECT MASK 2 121.075 26.94 121.155 29.758 ;
      RECT MASK 2 121.407 26.94 121.487 29.758 ;
      RECT MASK 2 121.739 26.94 121.819 29.758 ;
      RECT MASK 2 122.071 26.94 122.151 29.758 ;
      RECT MASK 2 122.403 26.94 122.483 29.758 ;
      RECT MASK 2 122.735 26.94 122.815 29.758 ;
      RECT MASK 2 123.067 26.94 123.147 29.758 ;
      RECT MASK 2 123.399 26.94 123.479 29.758 ;
      RECT MASK 2 123.731 26.94 123.811 29.758 ;
      RECT MASK 2 124.063 26.94 124.143 29.758 ;
      RECT MASK 2 124.395 26.94 124.475 29.758 ;
      RECT MASK 2 124.727 26.94 124.807 29.758 ;
      RECT MASK 2 125.059 26.94 125.139 29.758 ;
      RECT MASK 2 125.391 26.94 125.471 29.758 ;
      RECT MASK 2 125.723 26.94 125.803 29.758 ;
      RECT MASK 2 126.055 26.94 126.135 29.758 ;
      RECT MASK 2 126.577 27.64 126.657 28.012 ;
      RECT MASK 2 4.901 28.009 5.021 33.101 ;
      RECT MASK 2 5.341 28.009 5.461 33.101 ;
      RECT MASK 2 5.781 28.009 5.901 33.101 ;
      RECT MASK 2 6.221 28.009 6.341 33.101 ;
      RECT MASK 2 6.661 28.009 6.781 33.101 ;
      RECT MASK 2 7.101 28.009 7.221 33.101 ;
      RECT MASK 2 7.541 28.009 7.661 33.101 ;
      RECT MASK 2 7.981 28.009 8.101 33.101 ;
      RECT MASK 2 8.421 28.009 8.541 33.101 ;
      RECT MASK 2 8.861 28.009 8.981 33.101 ;
      RECT MASK 2 9.301 28.009 9.421 33.101 ;
      RECT MASK 2 9.741 28.009 9.861 33.101 ;
      RECT MASK 2 10.181 28.009 10.301 33.101 ;
      RECT MASK 2 10.621 28.009 10.741 33.101 ;
      RECT MASK 2 11.519 28.009 11.639 33.101 ;
      RECT MASK 2 11.959 28.009 12.079 33.101 ;
      RECT MASK 2 12.399 28.009 12.519 33.101 ;
      RECT MASK 2 12.839 28.009 12.959 33.101 ;
      RECT MASK 2 13.279 28.009 13.399 33.101 ;
      RECT MASK 2 13.719 28.009 13.839 33.101 ;
      RECT MASK 2 14.159 28.009 14.279 33.101 ;
      RECT MASK 2 14.599 28.009 14.719 33.101 ;
      RECT MASK 2 15.039 28.009 15.159 33.101 ;
      RECT MASK 2 15.479 28.009 15.599 33.101 ;
      RECT MASK 2 15.919 28.009 16.039 33.101 ;
      RECT MASK 2 16.359 28.009 16.479 33.101 ;
      RECT MASK 2 16.799 28.009 16.919 33.101 ;
      RECT MASK 2 17.239 28.009 17.359 33.101 ;
      RECT MASK 2 18.137 28.009 18.257 33.101 ;
      RECT MASK 2 18.577 28.009 18.697 33.101 ;
      RECT MASK 2 19.017 28.009 19.137 33.101 ;
      RECT MASK 2 19.457 28.009 19.577 33.101 ;
      RECT MASK 2 19.897 28.009 20.017 33.101 ;
      RECT MASK 2 20.337 28.009 20.457 33.101 ;
      RECT MASK 2 20.777 28.009 20.897 33.101 ;
      RECT MASK 2 21.217 28.009 21.337 33.101 ;
      RECT MASK 2 21.657 28.009 21.777 33.101 ;
      RECT MASK 2 22.097 28.009 22.217 33.101 ;
      RECT MASK 2 22.537 28.009 22.657 33.101 ;
      RECT MASK 2 22.977 28.009 23.097 33.101 ;
      RECT MASK 2 23.417 28.009 23.537 33.101 ;
      RECT MASK 2 23.857 28.009 23.977 33.101 ;
      RECT MASK 2 24.755 28.009 24.875 33.101 ;
      RECT MASK 2 25.195 28.009 25.315 33.101 ;
      RECT MASK 2 25.635 28.009 25.755 33.101 ;
      RECT MASK 2 26.075 28.009 26.195 33.101 ;
      RECT MASK 2 26.515 28.009 26.635 33.101 ;
      RECT MASK 2 26.955 28.009 27.075 33.101 ;
      RECT MASK 2 27.395 28.009 27.515 33.101 ;
      RECT MASK 2 27.835 28.009 27.955 33.101 ;
      RECT MASK 2 28.275 28.009 28.395 33.101 ;
      RECT MASK 2 28.715 28.009 28.835 33.101 ;
      RECT MASK 2 29.155 28.009 29.275 33.101 ;
      RECT MASK 2 29.595 28.009 29.715 33.101 ;
      RECT MASK 2 30.035 28.009 30.155 33.101 ;
      RECT MASK 2 30.475 28.009 30.595 33.101 ;
      RECT MASK 2 31.373 28.009 31.493 33.101 ;
      RECT MASK 2 31.813 28.009 31.933 33.101 ;
      RECT MASK 2 32.253 28.009 32.373 33.101 ;
      RECT MASK 2 32.693 28.009 32.813 33.101 ;
      RECT MASK 2 33.133 28.009 33.253 33.101 ;
      RECT MASK 2 33.573 28.009 33.693 33.101 ;
      RECT MASK 2 34.013 28.009 34.133 33.101 ;
      RECT MASK 2 34.453 28.009 34.573 33.101 ;
      RECT MASK 2 34.893 28.009 35.013 33.101 ;
      RECT MASK 2 35.333 28.009 35.453 33.101 ;
      RECT MASK 2 35.773 28.009 35.893 33.101 ;
      RECT MASK 2 36.213 28.009 36.333 33.101 ;
      RECT MASK 2 36.653 28.009 36.773 33.101 ;
      RECT MASK 2 37.093 28.009 37.213 33.101 ;
      RECT MASK 2 37.991 28.009 38.111 33.101 ;
      RECT MASK 2 38.431 28.009 38.551 33.101 ;
      RECT MASK 2 38.871 28.009 38.991 33.101 ;
      RECT MASK 2 39.311 28.009 39.431 33.101 ;
      RECT MASK 2 39.751 28.009 39.871 33.101 ;
      RECT MASK 2 40.191 28.009 40.311 33.101 ;
      RECT MASK 2 40.631 28.009 40.751 33.101 ;
      RECT MASK 2 41.071 28.009 41.191 33.101 ;
      RECT MASK 2 41.511 28.009 41.631 33.101 ;
      RECT MASK 2 41.951 28.009 42.071 33.101 ;
      RECT MASK 2 42.391 28.009 42.511 33.101 ;
      RECT MASK 2 42.831 28.009 42.951 33.101 ;
      RECT MASK 2 43.271 28.009 43.391 33.101 ;
      RECT MASK 2 43.711 28.009 43.831 33.101 ;
      RECT MASK 2 44.609 28.009 44.729 33.101 ;
      RECT MASK 2 45.049 28.009 45.169 33.101 ;
      RECT MASK 2 45.489 28.009 45.609 33.101 ;
      RECT MASK 2 45.929 28.009 46.049 33.101 ;
      RECT MASK 2 46.369 28.009 46.489 33.101 ;
      RECT MASK 2 46.809 28.009 46.929 33.101 ;
      RECT MASK 2 47.249 28.009 47.369 33.101 ;
      RECT MASK 2 47.689 28.009 47.809 33.101 ;
      RECT MASK 2 48.129 28.009 48.249 33.101 ;
      RECT MASK 2 48.569 28.009 48.689 33.101 ;
      RECT MASK 2 49.009 28.009 49.129 33.101 ;
      RECT MASK 2 49.449 28.009 49.569 33.101 ;
      RECT MASK 2 49.889 28.009 50.009 33.101 ;
      RECT MASK 2 50.329 28.009 50.449 33.101 ;
      RECT MASK 2 51.227 28.009 51.347 33.101 ;
      RECT MASK 2 51.667 28.009 51.787 33.101 ;
      RECT MASK 2 52.107 28.009 52.227 33.101 ;
      RECT MASK 2 52.547 28.009 52.667 33.101 ;
      RECT MASK 2 52.987 28.009 53.107 33.101 ;
      RECT MASK 2 53.427 28.009 53.547 33.101 ;
      RECT MASK 2 53.867 28.009 53.987 33.101 ;
      RECT MASK 2 54.307 28.009 54.427 33.101 ;
      RECT MASK 2 54.747 28.009 54.867 33.101 ;
      RECT MASK 2 55.187 28.009 55.307 33.101 ;
      RECT MASK 2 55.627 28.009 55.747 33.101 ;
      RECT MASK 2 56.067 28.009 56.187 33.101 ;
      RECT MASK 2 56.507 28.009 56.627 33.101 ;
      RECT MASK 2 56.947 28.009 57.067 33.101 ;
      RECT MASK 2 57.845 28.009 57.965 33.101 ;
      RECT MASK 2 58.285 28.009 58.405 33.101 ;
      RECT MASK 2 58.725 28.009 58.845 33.101 ;
      RECT MASK 2 59.165 28.009 59.285 33.101 ;
      RECT MASK 2 59.605 28.009 59.725 33.101 ;
      RECT MASK 2 60.045 28.009 60.165 33.101 ;
      RECT MASK 2 60.485 28.009 60.605 33.101 ;
      RECT MASK 2 60.925 28.009 61.045 33.101 ;
      RECT MASK 2 61.365 28.009 61.485 33.101 ;
      RECT MASK 2 61.805 28.009 61.925 33.101 ;
      RECT MASK 2 62.245 28.009 62.365 33.101 ;
      RECT MASK 2 62.685 28.009 62.805 33.101 ;
      RECT MASK 2 63.125 28.009 63.245 33.101 ;
      RECT MASK 2 63.565 28.009 63.685 33.101 ;
      RECT MASK 2 64.463 28.009 64.583 33.101 ;
      RECT MASK 2 64.903 28.009 65.023 33.101 ;
      RECT MASK 2 65.343 28.009 65.463 33.101 ;
      RECT MASK 2 65.783 28.009 65.903 33.101 ;
      RECT MASK 2 66.223 28.009 66.343 33.101 ;
      RECT MASK 2 66.663 28.009 66.783 33.101 ;
      RECT MASK 2 67.103 28.009 67.223 33.101 ;
      RECT MASK 2 67.543 28.009 67.663 33.101 ;
      RECT MASK 2 67.983 28.009 68.103 33.101 ;
      RECT MASK 2 68.423 28.009 68.543 33.101 ;
      RECT MASK 2 68.863 28.009 68.983 33.101 ;
      RECT MASK 2 69.303 28.009 69.423 33.101 ;
      RECT MASK 2 69.743 28.009 69.863 33.101 ;
      RECT MASK 2 70.183 28.009 70.303 33.101 ;
      RECT MASK 2 71.081 28.009 71.201 33.101 ;
      RECT MASK 2 71.521 28.009 71.641 33.101 ;
      RECT MASK 2 71.961 28.009 72.081 33.101 ;
      RECT MASK 2 72.401 28.009 72.521 33.101 ;
      RECT MASK 2 72.841 28.009 72.961 33.101 ;
      RECT MASK 2 73.281 28.009 73.401 33.101 ;
      RECT MASK 2 73.721 28.009 73.841 33.101 ;
      RECT MASK 2 74.161 28.009 74.281 33.101 ;
      RECT MASK 2 74.601 28.009 74.721 33.101 ;
      RECT MASK 2 75.041 28.009 75.161 33.101 ;
      RECT MASK 2 75.481 28.009 75.601 33.101 ;
      RECT MASK 2 75.921 28.009 76.041 33.101 ;
      RECT MASK 2 76.361 28.009 76.481 33.101 ;
      RECT MASK 2 76.801 28.009 76.921 33.101 ;
      RECT MASK 2 77.699 28.009 77.819 33.101 ;
      RECT MASK 2 78.139 28.009 78.259 33.101 ;
      RECT MASK 2 78.579 28.009 78.699 33.101 ;
      RECT MASK 2 79.019 28.009 79.139 33.101 ;
      RECT MASK 2 79.459 28.009 79.579 33.101 ;
      RECT MASK 2 79.899 28.009 80.019 33.101 ;
      RECT MASK 2 80.339 28.009 80.459 33.101 ;
      RECT MASK 2 80.779 28.009 80.899 33.101 ;
      RECT MASK 2 81.219 28.009 81.339 33.101 ;
      RECT MASK 2 81.659 28.009 81.779 33.101 ;
      RECT MASK 2 82.099 28.009 82.219 33.101 ;
      RECT MASK 2 82.539 28.009 82.659 33.101 ;
      RECT MASK 2 82.979 28.009 83.099 33.101 ;
      RECT MASK 2 83.419 28.009 83.539 33.101 ;
      RECT MASK 2 84.317 28.009 84.437 33.101 ;
      RECT MASK 2 84.757 28.009 84.877 33.101 ;
      RECT MASK 2 85.197 28.009 85.317 33.101 ;
      RECT MASK 2 85.637 28.009 85.757 33.101 ;
      RECT MASK 2 86.077 28.009 86.197 33.101 ;
      RECT MASK 2 86.517 28.009 86.637 33.101 ;
      RECT MASK 2 86.957 28.009 87.077 33.101 ;
      RECT MASK 2 87.397 28.009 87.517 33.101 ;
      RECT MASK 2 87.837 28.009 87.957 33.101 ;
      RECT MASK 2 88.277 28.009 88.397 33.101 ;
      RECT MASK 2 88.717 28.009 88.837 33.101 ;
      RECT MASK 2 89.157 28.009 89.277 33.101 ;
      RECT MASK 2 89.597 28.009 89.717 33.101 ;
      RECT MASK 2 90.037 28.009 90.157 33.101 ;
      RECT MASK 2 90.935 28.009 91.055 33.101 ;
      RECT MASK 2 91.375 28.009 91.495 33.101 ;
      RECT MASK 2 91.815 28.009 91.935 33.101 ;
      RECT MASK 2 92.255 28.009 92.375 33.101 ;
      RECT MASK 2 92.695 28.009 92.815 33.101 ;
      RECT MASK 2 93.135 28.009 93.255 33.101 ;
      RECT MASK 2 93.575 28.009 93.695 33.101 ;
      RECT MASK 2 94.015 28.009 94.135 33.101 ;
      RECT MASK 2 94.455 28.009 94.575 33.101 ;
      RECT MASK 2 94.895 28.009 95.015 33.101 ;
      RECT MASK 2 95.335 28.009 95.455 33.101 ;
      RECT MASK 2 95.775 28.009 95.895 33.101 ;
      RECT MASK 2 96.215 28.009 96.335 33.101 ;
      RECT MASK 2 96.655 28.009 96.775 33.101 ;
      RECT MASK 2 97.553 28.009 97.673 33.101 ;
      RECT MASK 2 97.993 28.009 98.113 33.101 ;
      RECT MASK 2 98.433 28.009 98.553 33.101 ;
      RECT MASK 2 98.873 28.009 98.993 33.101 ;
      RECT MASK 2 99.313 28.009 99.433 33.101 ;
      RECT MASK 2 99.753 28.009 99.873 33.101 ;
      RECT MASK 2 100.193 28.009 100.313 33.101 ;
      RECT MASK 2 100.633 28.009 100.753 33.101 ;
      RECT MASK 2 101.073 28.009 101.193 33.101 ;
      RECT MASK 2 101.513 28.009 101.633 33.101 ;
      RECT MASK 2 101.953 28.009 102.073 33.101 ;
      RECT MASK 2 102.393 28.009 102.513 33.101 ;
      RECT MASK 2 102.833 28.009 102.953 33.101 ;
      RECT MASK 2 103.273 28.009 103.393 33.101 ;
      RECT MASK 2 104.171 28.009 104.291 33.101 ;
      RECT MASK 2 104.611 28.009 104.731 33.101 ;
      RECT MASK 2 105.051 28.009 105.171 33.101 ;
      RECT MASK 2 105.491 28.009 105.611 33.101 ;
      RECT MASK 2 105.931 28.009 106.051 33.101 ;
      RECT MASK 2 106.371 28.009 106.491 33.101 ;
      RECT MASK 2 106.811 28.009 106.931 33.101 ;
      RECT MASK 2 107.251 28.009 107.371 33.101 ;
      RECT MASK 2 107.691 28.009 107.811 33.101 ;
      RECT MASK 2 108.131 28.009 108.251 33.101 ;
      RECT MASK 2 108.571 28.009 108.691 33.101 ;
      RECT MASK 2 109.011 28.009 109.131 33.101 ;
      RECT MASK 2 109.451 28.009 109.571 33.101 ;
      RECT MASK 2 109.891 28.009 110.011 33.101 ;
      RECT MASK 2 126.577 28.42 126.657 28.792 ;
      RECT MASK 2 126.577 29.2005 126.657 29.5725 ;
      RECT MASK 2 116.427 30.206 116.507 30.51 ;
      RECT MASK 2 116.759 30.206 116.839 30.51 ;
      RECT MASK 2 117.091 30.206 117.171 30.51 ;
      RECT MASK 2 117.423 30.206 117.503 30.51 ;
      RECT MASK 2 117.755 30.206 117.835 30.51 ;
      RECT MASK 2 118.087 30.206 118.167 30.51 ;
      RECT MASK 2 118.419 30.206 118.499 30.51 ;
      RECT MASK 2 118.751 30.206 118.831 30.51 ;
      RECT MASK 2 119.083 30.206 119.163 30.51 ;
      RECT MASK 2 119.415 30.206 119.495 30.51 ;
      RECT MASK 2 119.747 30.206 119.827 30.51 ;
      RECT MASK 2 120.079 30.206 120.159 30.51 ;
      RECT MASK 2 120.411 30.206 120.491 30.51 ;
      RECT MASK 2 120.743 30.206 120.823 30.51 ;
      RECT MASK 2 121.075 30.206 121.155 30.51 ;
      RECT MASK 2 121.407 30.206 121.487 30.51 ;
      RECT MASK 2 121.739 30.206 121.819 30.51 ;
      RECT MASK 2 122.071 30.206 122.151 30.51 ;
      RECT MASK 2 122.403 30.206 122.483 30.51 ;
      RECT MASK 2 122.735 30.206 122.815 30.51 ;
      RECT MASK 2 123.067 30.206 123.147 30.51 ;
      RECT MASK 2 123.399 30.206 123.479 30.51 ;
      RECT MASK 2 123.731 30.206 123.811 30.51 ;
      RECT MASK 2 124.063 30.206 124.143 30.51 ;
      RECT MASK 2 124.395 30.206 124.475 30.51 ;
      RECT MASK 2 124.727 30.206 124.807 30.51 ;
      RECT MASK 2 125.059 30.206 125.139 30.51 ;
      RECT MASK 2 125.391 30.206 125.471 30.51 ;
      RECT MASK 2 125.723 30.206 125.803 30.51 ;
      RECT MASK 2 126.055 30.206 126.135 30.51 ;
      RECT MASK 2 128.975 31.11 129.095 73.077 ;
      RECT MASK 2 114.221 31.136 114.301 31.468 ;
      RECT MASK 2 114.553 31.136 114.633 31.468 ;
      RECT MASK 2 114.885 31.136 114.965 31.468 ;
      RECT MASK 2 115.217 31.136 115.297 31.468 ;
      RECT MASK 2 115.881 31.136 115.961 31.468 ;
      RECT MASK 2 116.545 31.136 116.625 31.468 ;
      RECT MASK 2 116.877 31.136 116.957 31.468 ;
      RECT MASK 2 117.209 31.136 117.289 31.468 ;
      RECT MASK 2 117.541 31.136 117.621 31.468 ;
      RECT MASK 2 118.205 31.136 118.285 31.468 ;
      RECT MASK 2 118.869 31.136 118.949 31.468 ;
      RECT MASK 2 119.201 31.136 119.281 31.468 ;
      RECT MASK 2 119.533 31.136 119.613 31.468 ;
      RECT MASK 2 120.197 31.136 120.277 31.468 ;
      RECT MASK 2 120.861 31.136 120.941 31.468 ;
      RECT MASK 2 121.193 31.136 121.273 31.468 ;
      RECT MASK 2 121.525 31.136 121.605 31.468 ;
      RECT MASK 2 121.857 31.136 121.937 31.468 ;
      RECT MASK 2 122.521 31.136 122.601 31.468 ;
      RECT MASK 2 123.185 31.136 123.265 31.468 ;
      RECT MASK 2 123.517 31.136 123.597 31.468 ;
      RECT MASK 2 123.849 31.136 123.929 31.468 ;
      RECT MASK 2 125.509 31.136 125.589 31.468 ;
      RECT MASK 2 125.841 31.136 125.921 31.468 ;
      RECT MASK 2 126.173 31.136 126.253 31.468 ;
      RECT MASK 2 126.837 31.136 126.917 31.468 ;
      RECT MASK 2 127.501 31.136 127.581 31.468 ;
      RECT MASK 2 127.833 31.136 127.913 31.468 ;
      RECT MASK 2 128.165 31.136 128.245 31.468 ;
      RECT MASK 2 128.497 31.136 128.577 31.468 ;
      RECT MASK 2 124.2055 32.16 124.2855 71.973 ;
      RECT MASK 2 124.5375 32.16 124.6175 71.973 ;
      RECT MASK 2 124.8695 32.16 124.9495 71.973 ;
      RECT MASK 2 125.2015 32.16 125.2815 71.973 ;
      RECT MASK 2 125.5335 32.16 125.6135 71.973 ;
      RECT MASK 2 125.8655 32.16 125.9455 71.973 ;
      RECT MASK 2 126.1975 32.16 126.2775 71.973 ;
      RECT MASK 2 126.5295 32.16 126.6095 71.973 ;
      RECT MASK 2 126.8615 32.16 126.9415 71.973 ;
      RECT MASK 2 127.1935 32.16 127.2735 71.973 ;
      RECT MASK 2 127.5255 32.16 127.6055 71.973 ;
      RECT MASK 2 127.8575 32.16 127.9375 71.973 ;
      RECT MASK 2 112.5865 32.749 112.7065 34.469 ;
      RECT MASK 2 113.0265 32.749 113.1465 34.469 ;
      RECT MASK 2 113.4665 32.749 113.5865 34.469 ;
      RECT MASK 2 113.9065 32.749 114.0265 34.469 ;
      RECT MASK 2 114.3465 32.749 114.4665 34.469 ;
      RECT MASK 2 114.7865 32.749 114.9065 34.469 ;
      RECT MASK 2 115.2265 32.749 115.3465 34.469 ;
      RECT MASK 2 115.6665 32.749 115.7865 34.469 ;
      RECT MASK 2 116.1065 32.749 116.2265 34.469 ;
      RECT MASK 2 116.5465 32.749 116.6665 34.469 ;
      RECT MASK 2 117.4265 32.749 117.5465 34.469 ;
      RECT MASK 2 117.8665 32.749 117.9865 34.469 ;
      RECT MASK 2 118.3065 32.749 118.4265 34.469 ;
      RECT MASK 2 118.7465 32.749 118.8665 34.469 ;
      RECT MASK 2 119.1865 32.749 119.3065 34.469 ;
      RECT MASK 2 119.6265 32.749 119.7465 34.469 ;
      RECT MASK 2 120.0665 32.749 120.1865 34.469 ;
      RECT MASK 2 120.5065 32.749 120.6265 34.469 ;
      RECT MASK 2 120.9465 32.749 121.0665 34.469 ;
      RECT MASK 2 121.3865 32.749 121.5065 34.469 ;
      RECT MASK 2 121.8265 32.749 121.9465 34.469 ;
      RECT MASK 2 122.2665 32.749 122.3865 34.469 ;
      RECT MASK 2 122.7065 32.749 122.8265 34.469 ;
      RECT MASK 2 123.1465 32.749 123.2665 34.469 ;
      RECT MASK 2 123.5865 32.749 123.7065 34.469 ;
      RECT MASK 2 4.931 33.27 4.991 33.51 ;
      RECT MASK 2 5.371 33.27 5.431 33.51 ;
      RECT MASK 2 5.811 33.27 5.871 33.51 ;
      RECT MASK 2 6.251 33.27 6.311 33.51 ;
      RECT MASK 2 6.691 33.27 6.751 33.51 ;
      RECT MASK 2 7.131 33.27 7.191 33.51 ;
      RECT MASK 2 7.571 33.27 7.631 33.51 ;
      RECT MASK 2 8.011 33.27 8.071 33.51 ;
      RECT MASK 2 8.451 33.27 8.511 33.51 ;
      RECT MASK 2 8.891 33.27 8.951 33.51 ;
      RECT MASK 2 9.331 33.27 9.391 33.51 ;
      RECT MASK 2 9.771 33.27 9.831 33.51 ;
      RECT MASK 2 10.211 33.27 10.271 33.51 ;
      RECT MASK 2 10.651 33.27 10.711 33.51 ;
      RECT MASK 2 11.549 33.27 11.609 33.51 ;
      RECT MASK 2 11.989 33.27 12.049 33.51 ;
      RECT MASK 2 12.429 33.27 12.489 33.51 ;
      RECT MASK 2 12.869 33.27 12.929 33.51 ;
      RECT MASK 2 13.309 33.27 13.369 33.51 ;
      RECT MASK 2 13.749 33.27 13.809 33.51 ;
      RECT MASK 2 14.189 33.27 14.249 33.51 ;
      RECT MASK 2 14.629 33.27 14.689 33.51 ;
      RECT MASK 2 15.069 33.27 15.129 33.51 ;
      RECT MASK 2 15.509 33.27 15.569 33.51 ;
      RECT MASK 2 15.949 33.27 16.009 33.51 ;
      RECT MASK 2 16.389 33.27 16.449 33.51 ;
      RECT MASK 2 16.829 33.27 16.889 33.51 ;
      RECT MASK 2 17.269 33.27 17.329 33.51 ;
      RECT MASK 2 18.167 33.27 18.227 33.51 ;
      RECT MASK 2 18.607 33.27 18.667 33.51 ;
      RECT MASK 2 19.047 33.27 19.107 33.51 ;
      RECT MASK 2 19.487 33.27 19.547 33.51 ;
      RECT MASK 2 19.927 33.27 19.987 33.51 ;
      RECT MASK 2 20.367 33.27 20.427 33.51 ;
      RECT MASK 2 20.807 33.27 20.867 33.51 ;
      RECT MASK 2 21.247 33.27 21.307 33.51 ;
      RECT MASK 2 21.687 33.27 21.747 33.51 ;
      RECT MASK 2 22.127 33.27 22.187 33.51 ;
      RECT MASK 2 22.567 33.27 22.627 33.51 ;
      RECT MASK 2 23.007 33.27 23.067 33.51 ;
      RECT MASK 2 23.447 33.27 23.507 33.51 ;
      RECT MASK 2 23.887 33.27 23.947 33.51 ;
      RECT MASK 2 24.785 33.27 24.845 33.51 ;
      RECT MASK 2 25.225 33.27 25.285 33.51 ;
      RECT MASK 2 25.665 33.27 25.725 33.51 ;
      RECT MASK 2 26.105 33.27 26.165 33.51 ;
      RECT MASK 2 26.545 33.27 26.605 33.51 ;
      RECT MASK 2 26.985 33.27 27.045 33.51 ;
      RECT MASK 2 27.425 33.27 27.485 33.51 ;
      RECT MASK 2 27.865 33.27 27.925 33.51 ;
      RECT MASK 2 28.305 33.27 28.365 33.51 ;
      RECT MASK 2 28.745 33.27 28.805 33.51 ;
      RECT MASK 2 29.185 33.27 29.245 33.51 ;
      RECT MASK 2 29.625 33.27 29.685 33.51 ;
      RECT MASK 2 30.065 33.27 30.125 33.51 ;
      RECT MASK 2 30.505 33.27 30.565 33.51 ;
      RECT MASK 2 31.403 33.27 31.463 33.51 ;
      RECT MASK 2 31.843 33.27 31.903 33.51 ;
      RECT MASK 2 32.283 33.27 32.343 33.51 ;
      RECT MASK 2 32.723 33.27 32.783 33.51 ;
      RECT MASK 2 33.163 33.27 33.223 33.51 ;
      RECT MASK 2 33.603 33.27 33.663 33.51 ;
      RECT MASK 2 34.043 33.27 34.103 33.51 ;
      RECT MASK 2 34.483 33.27 34.543 33.51 ;
      RECT MASK 2 34.923 33.27 34.983 33.51 ;
      RECT MASK 2 35.363 33.27 35.423 33.51 ;
      RECT MASK 2 35.803 33.27 35.863 33.51 ;
      RECT MASK 2 36.243 33.27 36.303 33.51 ;
      RECT MASK 2 36.683 33.27 36.743 33.51 ;
      RECT MASK 2 37.123 33.27 37.183 33.51 ;
      RECT MASK 2 38.021 33.27 38.081 33.51 ;
      RECT MASK 2 38.461 33.27 38.521 33.51 ;
      RECT MASK 2 38.901 33.27 38.961 33.51 ;
      RECT MASK 2 39.341 33.27 39.401 33.51 ;
      RECT MASK 2 39.781 33.27 39.841 33.51 ;
      RECT MASK 2 40.221 33.27 40.281 33.51 ;
      RECT MASK 2 40.661 33.27 40.721 33.51 ;
      RECT MASK 2 41.101 33.27 41.161 33.51 ;
      RECT MASK 2 41.541 33.27 41.601 33.51 ;
      RECT MASK 2 42.861 33.27 42.921 33.51 ;
      RECT MASK 2 43.301 33.27 43.361 33.51 ;
      RECT MASK 2 43.741 33.27 43.801 33.51 ;
      RECT MASK 2 44.639 33.27 44.699 33.51 ;
      RECT MASK 2 45.079 33.27 45.139 33.51 ;
      RECT MASK 2 45.519 33.27 45.579 33.51 ;
      RECT MASK 2 45.959 33.27 46.019 33.51 ;
      RECT MASK 2 46.399 33.27 46.459 33.51 ;
      RECT MASK 2 46.839 33.27 46.899 33.51 ;
      RECT MASK 2 47.279 33.27 47.339 33.51 ;
      RECT MASK 2 47.719 33.27 47.779 33.51 ;
      RECT MASK 2 48.159 33.27 48.219 33.51 ;
      RECT MASK 2 48.599 33.27 48.659 33.51 ;
      RECT MASK 2 49.039 33.27 49.099 33.51 ;
      RECT MASK 2 49.479 33.27 49.539 33.51 ;
      RECT MASK 2 49.919 33.27 49.979 33.51 ;
      RECT MASK 2 50.359 33.27 50.419 33.51 ;
      RECT MASK 2 51.257 33.27 51.317 33.51 ;
      RECT MASK 2 51.697 33.27 51.757 33.51 ;
      RECT MASK 2 52.137 33.27 52.197 33.51 ;
      RECT MASK 2 52.577 33.27 52.637 33.51 ;
      RECT MASK 2 53.017 33.27 53.077 33.51 ;
      RECT MASK 2 53.457 33.27 53.517 33.51 ;
      RECT MASK 2 53.897 33.27 53.957 33.51 ;
      RECT MASK 2 54.337 33.27 54.397 33.51 ;
      RECT MASK 2 54.777 33.27 54.837 33.51 ;
      RECT MASK 2 55.217 33.27 55.277 33.51 ;
      RECT MASK 2 55.657 33.27 55.717 33.51 ;
      RECT MASK 2 56.097 33.27 56.157 33.51 ;
      RECT MASK 2 56.537 33.27 56.597 33.51 ;
      RECT MASK 2 56.977 33.27 57.037 33.51 ;
      RECT MASK 2 57.875 33.27 57.935 33.51 ;
      RECT MASK 2 58.315 33.27 58.375 33.51 ;
      RECT MASK 2 58.755 33.27 58.815 33.51 ;
      RECT MASK 2 59.195 33.27 59.255 33.51 ;
      RECT MASK 2 59.635 33.27 59.695 33.51 ;
      RECT MASK 2 60.075 33.27 60.135 33.51 ;
      RECT MASK 2 60.515 33.27 60.575 33.51 ;
      RECT MASK 2 60.955 33.27 61.015 33.51 ;
      RECT MASK 2 61.395 33.27 61.455 33.51 ;
      RECT MASK 2 61.835 33.27 61.895 33.51 ;
      RECT MASK 2 62.275 33.27 62.335 33.51 ;
      RECT MASK 2 62.715 33.27 62.775 33.51 ;
      RECT MASK 2 63.155 33.27 63.215 33.51 ;
      RECT MASK 2 63.595 33.27 63.655 33.51 ;
      RECT MASK 2 64.493 33.27 64.553 33.51 ;
      RECT MASK 2 64.933 33.27 64.993 33.51 ;
      RECT MASK 2 65.373 33.27 65.433 33.51 ;
      RECT MASK 2 65.813 33.27 65.873 33.51 ;
      RECT MASK 2 66.253 33.27 66.313 33.51 ;
      RECT MASK 2 66.693 33.27 66.753 33.51 ;
      RECT MASK 2 67.133 33.27 67.193 33.51 ;
      RECT MASK 2 67.573 33.27 67.633 33.51 ;
      RECT MASK 2 68.013 33.27 68.073 33.51 ;
      RECT MASK 2 68.453 33.27 68.513 33.51 ;
      RECT MASK 2 68.893 33.27 68.953 33.51 ;
      RECT MASK 2 69.333 33.27 69.393 33.51 ;
      RECT MASK 2 69.773 33.27 69.833 33.51 ;
      RECT MASK 2 70.213 33.27 70.273 33.51 ;
      RECT MASK 2 71.111 33.27 71.171 33.51 ;
      RECT MASK 2 71.551 33.27 71.611 33.51 ;
      RECT MASK 2 71.991 33.27 72.051 33.51 ;
      RECT MASK 2 72.431 33.27 72.491 33.51 ;
      RECT MASK 2 72.871 33.27 72.931 33.51 ;
      RECT MASK 2 73.311 33.27 73.371 33.51 ;
      RECT MASK 2 73.751 33.27 73.811 33.51 ;
      RECT MASK 2 74.191 33.27 74.251 33.51 ;
      RECT MASK 2 74.631 33.27 74.691 33.51 ;
      RECT MASK 2 75.071 33.27 75.131 33.51 ;
      RECT MASK 2 75.511 33.27 75.571 33.51 ;
      RECT MASK 2 75.951 33.27 76.011 33.51 ;
      RECT MASK 2 76.391 33.27 76.451 33.51 ;
      RECT MASK 2 76.831 33.27 76.891 33.51 ;
      RECT MASK 2 77.729 33.27 77.789 33.51 ;
      RECT MASK 2 78.169 33.27 78.229 33.51 ;
      RECT MASK 2 78.609 33.27 78.669 33.51 ;
      RECT MASK 2 79.049 33.27 79.109 33.51 ;
      RECT MASK 2 79.489 33.27 79.549 33.51 ;
      RECT MASK 2 79.929 33.27 79.989 33.51 ;
      RECT MASK 2 80.369 33.27 80.429 33.51 ;
      RECT MASK 2 80.809 33.27 80.869 33.51 ;
      RECT MASK 2 81.249 33.27 81.309 33.51 ;
      RECT MASK 2 81.689 33.27 81.749 33.51 ;
      RECT MASK 2 82.129 33.27 82.189 33.51 ;
      RECT MASK 2 83.449 33.27 83.509 33.51 ;
      RECT MASK 2 84.347 33.27 84.407 33.51 ;
      RECT MASK 2 84.787 33.27 84.847 33.51 ;
      RECT MASK 2 85.227 33.27 85.287 33.51 ;
      RECT MASK 2 85.667 33.27 85.727 33.51 ;
      RECT MASK 2 86.107 33.27 86.167 33.51 ;
      RECT MASK 2 86.547 33.27 86.607 33.51 ;
      RECT MASK 2 86.987 33.27 87.047 33.51 ;
      RECT MASK 2 87.427 33.27 87.487 33.51 ;
      RECT MASK 2 87.867 33.27 87.927 33.51 ;
      RECT MASK 2 88.307 33.27 88.367 33.51 ;
      RECT MASK 2 88.747 33.27 88.807 33.51 ;
      RECT MASK 2 89.187 33.27 89.247 33.51 ;
      RECT MASK 2 89.627 33.27 89.687 33.51 ;
      RECT MASK 2 90.067 33.27 90.127 33.51 ;
      RECT MASK 2 90.965 33.27 91.025 33.51 ;
      RECT MASK 2 91.405 33.27 91.465 33.51 ;
      RECT MASK 2 91.845 33.27 91.905 33.51 ;
      RECT MASK 2 92.285 33.27 92.345 33.51 ;
      RECT MASK 2 92.725 33.27 92.785 33.51 ;
      RECT MASK 2 93.165 33.27 93.225 33.51 ;
      RECT MASK 2 93.605 33.27 93.665 33.51 ;
      RECT MASK 2 94.045 33.27 94.105 33.51 ;
      RECT MASK 2 94.485 33.27 94.545 33.51 ;
      RECT MASK 2 94.925 33.27 94.985 33.51 ;
      RECT MASK 2 95.365 33.27 95.425 33.51 ;
      RECT MASK 2 95.805 33.27 95.865 33.51 ;
      RECT MASK 2 96.245 33.27 96.305 33.51 ;
      RECT MASK 2 96.685 33.27 96.745 33.51 ;
      RECT MASK 2 97.583 33.27 97.643 33.51 ;
      RECT MASK 2 98.023 33.27 98.083 33.51 ;
      RECT MASK 2 98.463 33.27 98.523 33.51 ;
      RECT MASK 2 98.903 33.27 98.963 33.51 ;
      RECT MASK 2 99.343 33.27 99.403 33.51 ;
      RECT MASK 2 99.783 33.27 99.843 33.51 ;
      RECT MASK 2 100.223 33.27 100.283 33.51 ;
      RECT MASK 2 100.663 33.27 100.723 33.51 ;
      RECT MASK 2 101.103 33.27 101.163 33.51 ;
      RECT MASK 2 101.543 33.27 101.603 33.51 ;
      RECT MASK 2 101.983 33.27 102.043 33.51 ;
      RECT MASK 2 102.423 33.27 102.483 33.51 ;
      RECT MASK 2 102.863 33.27 102.923 33.51 ;
      RECT MASK 2 103.303 33.27 103.363 33.51 ;
      RECT MASK 2 104.201 33.27 104.261 33.51 ;
      RECT MASK 2 104.641 33.27 104.701 33.51 ;
      RECT MASK 2 105.081 33.27 105.141 33.51 ;
      RECT MASK 2 105.521 33.27 105.581 33.51 ;
      RECT MASK 2 105.961 33.27 106.021 33.51 ;
      RECT MASK 2 106.401 33.27 106.461 33.51 ;
      RECT MASK 2 106.841 33.27 106.901 33.51 ;
      RECT MASK 2 107.281 33.27 107.341 33.51 ;
      RECT MASK 2 107.721 33.27 107.781 33.51 ;
      RECT MASK 2 108.161 33.27 108.221 33.51 ;
      RECT MASK 2 108.601 33.27 108.661 33.51 ;
      RECT MASK 2 109.041 33.27 109.101 33.51 ;
      RECT MASK 2 109.481 33.27 109.541 33.51 ;
      RECT MASK 2 109.921 33.27 109.981 33.51 ;
      RECT MASK 2 4.931 33.69 4.991 33.93 ;
      RECT MASK 2 5.371 33.69 5.431 33.93 ;
      RECT MASK 2 5.811 33.69 5.871 33.93 ;
      RECT MASK 2 6.251 33.69 6.311 33.93 ;
      RECT MASK 2 6.691 33.69 6.751 33.93 ;
      RECT MASK 2 7.131 33.69 7.191 33.93 ;
      RECT MASK 2 7.571 33.69 7.631 33.93 ;
      RECT MASK 2 8.011 33.69 8.071 33.93 ;
      RECT MASK 2 8.451 33.69 8.511 33.93 ;
      RECT MASK 2 8.891 33.69 8.951 33.93 ;
      RECT MASK 2 9.331 33.69 9.391 33.93 ;
      RECT MASK 2 9.771 33.69 9.831 33.93 ;
      RECT MASK 2 10.211 33.69 10.271 33.93 ;
      RECT MASK 2 10.651 33.69 10.711 33.93 ;
      RECT MASK 2 11.549 33.69 11.609 33.93 ;
      RECT MASK 2 11.989 33.69 12.049 33.93 ;
      RECT MASK 2 12.429 33.69 12.489 33.93 ;
      RECT MASK 2 12.869 33.69 12.929 33.93 ;
      RECT MASK 2 13.309 33.69 13.369 33.93 ;
      RECT MASK 2 13.749 33.69 13.809 33.93 ;
      RECT MASK 2 14.189 33.69 14.249 33.93 ;
      RECT MASK 2 14.629 33.69 14.689 33.93 ;
      RECT MASK 2 15.069 33.69 15.129 33.93 ;
      RECT MASK 2 15.509 33.69 15.569 33.93 ;
      RECT MASK 2 15.949 33.69 16.009 33.93 ;
      RECT MASK 2 16.389 33.69 16.449 33.93 ;
      RECT MASK 2 16.829 33.69 16.889 33.93 ;
      RECT MASK 2 17.269 33.69 17.329 33.93 ;
      RECT MASK 2 18.167 33.69 18.227 33.93 ;
      RECT MASK 2 18.607 33.69 18.667 33.93 ;
      RECT MASK 2 19.047 33.69 19.107 33.93 ;
      RECT MASK 2 19.487 33.69 19.547 33.93 ;
      RECT MASK 2 19.927 33.69 19.987 33.93 ;
      RECT MASK 2 20.367 33.69 20.427 33.93 ;
      RECT MASK 2 20.807 33.69 20.867 33.93 ;
      RECT MASK 2 21.247 33.69 21.307 33.93 ;
      RECT MASK 2 21.687 33.69 21.747 33.93 ;
      RECT MASK 2 22.127 33.69 22.187 33.93 ;
      RECT MASK 2 22.567 33.69 22.627 33.93 ;
      RECT MASK 2 23.007 33.69 23.067 33.93 ;
      RECT MASK 2 23.447 33.69 23.507 33.93 ;
      RECT MASK 2 23.887 33.69 23.947 33.93 ;
      RECT MASK 2 24.785 33.69 24.845 33.93 ;
      RECT MASK 2 25.225 33.69 25.285 33.93 ;
      RECT MASK 2 25.665 33.69 25.725 33.93 ;
      RECT MASK 2 26.105 33.69 26.165 33.93 ;
      RECT MASK 2 26.545 33.69 26.605 33.93 ;
      RECT MASK 2 26.985 33.69 27.045 33.93 ;
      RECT MASK 2 27.425 33.69 27.485 33.93 ;
      RECT MASK 2 27.865 33.69 27.925 33.93 ;
      RECT MASK 2 28.305 33.69 28.365 33.93 ;
      RECT MASK 2 28.745 33.69 28.805 33.93 ;
      RECT MASK 2 29.185 33.69 29.245 33.93 ;
      RECT MASK 2 29.625 33.69 29.685 33.93 ;
      RECT MASK 2 30.065 33.69 30.125 33.93 ;
      RECT MASK 2 30.505 33.69 30.565 33.93 ;
      RECT MASK 2 31.403 33.69 31.463 33.93 ;
      RECT MASK 2 31.843 33.69 31.903 33.93 ;
      RECT MASK 2 32.283 33.69 32.343 33.93 ;
      RECT MASK 2 32.723 33.69 32.783 33.93 ;
      RECT MASK 2 33.163 33.69 33.223 33.93 ;
      RECT MASK 2 33.603 33.69 33.663 33.93 ;
      RECT MASK 2 34.043 33.69 34.103 33.93 ;
      RECT MASK 2 34.483 33.69 34.543 33.93 ;
      RECT MASK 2 34.923 33.69 34.983 33.93 ;
      RECT MASK 2 35.363 33.69 35.423 33.93 ;
      RECT MASK 2 35.803 33.69 35.863 33.93 ;
      RECT MASK 2 36.243 33.69 36.303 33.93 ;
      RECT MASK 2 36.683 33.69 36.743 33.93 ;
      RECT MASK 2 37.123 33.69 37.183 33.93 ;
      RECT MASK 2 38.021 33.69 38.081 33.93 ;
      RECT MASK 2 38.461 33.69 38.521 33.93 ;
      RECT MASK 2 38.901 33.69 38.961 33.93 ;
      RECT MASK 2 39.341 33.69 39.401 33.93 ;
      RECT MASK 2 39.781 33.69 39.841 33.93 ;
      RECT MASK 2 40.221 33.69 40.281 33.93 ;
      RECT MASK 2 40.661 33.69 40.721 33.93 ;
      RECT MASK 2 41.101 33.69 41.161 33.93 ;
      RECT MASK 2 41.541 33.69 41.601 33.93 ;
      RECT MASK 2 42.861 33.69 42.921 33.93 ;
      RECT MASK 2 43.301 33.69 43.361 33.93 ;
      RECT MASK 2 43.741 33.69 43.801 33.93 ;
      RECT MASK 2 44.639 33.69 44.699 33.93 ;
      RECT MASK 2 45.079 33.69 45.139 33.93 ;
      RECT MASK 2 45.519 33.69 45.579 33.93 ;
      RECT MASK 2 45.959 33.69 46.019 33.93 ;
      RECT MASK 2 46.399 33.69 46.459 33.93 ;
      RECT MASK 2 46.839 33.69 46.899 33.93 ;
      RECT MASK 2 47.279 33.69 47.339 33.93 ;
      RECT MASK 2 47.719 33.69 47.779 33.93 ;
      RECT MASK 2 48.159 33.69 48.219 33.93 ;
      RECT MASK 2 48.599 33.69 48.659 33.93 ;
      RECT MASK 2 49.039 33.69 49.099 33.93 ;
      RECT MASK 2 49.479 33.69 49.539 33.93 ;
      RECT MASK 2 49.919 33.69 49.979 33.93 ;
      RECT MASK 2 50.359 33.69 50.419 33.93 ;
      RECT MASK 2 51.257 33.69 51.317 33.93 ;
      RECT MASK 2 51.697 33.69 51.757 33.93 ;
      RECT MASK 2 52.137 33.69 52.197 33.93 ;
      RECT MASK 2 52.577 33.69 52.637 33.93 ;
      RECT MASK 2 53.017 33.69 53.077 33.93 ;
      RECT MASK 2 53.457 33.69 53.517 33.93 ;
      RECT MASK 2 53.897 33.69 53.957 33.93 ;
      RECT MASK 2 54.337 33.69 54.397 33.93 ;
      RECT MASK 2 54.777 33.69 54.837 33.93 ;
      RECT MASK 2 55.217 33.69 55.277 33.93 ;
      RECT MASK 2 55.657 33.69 55.717 33.93 ;
      RECT MASK 2 56.097 33.69 56.157 33.93 ;
      RECT MASK 2 56.537 33.69 56.597 33.93 ;
      RECT MASK 2 56.977 33.69 57.037 33.93 ;
      RECT MASK 2 57.875 33.69 57.935 33.93 ;
      RECT MASK 2 58.315 33.69 58.375 33.93 ;
      RECT MASK 2 58.755 33.69 58.815 33.93 ;
      RECT MASK 2 59.195 33.69 59.255 33.93 ;
      RECT MASK 2 59.635 33.69 59.695 33.93 ;
      RECT MASK 2 60.075 33.69 60.135 33.93 ;
      RECT MASK 2 60.515 33.69 60.575 33.93 ;
      RECT MASK 2 60.955 33.69 61.015 33.93 ;
      RECT MASK 2 61.395 33.69 61.455 33.93 ;
      RECT MASK 2 61.835 33.69 61.895 33.93 ;
      RECT MASK 2 62.275 33.69 62.335 33.93 ;
      RECT MASK 2 62.715 33.69 62.775 33.93 ;
      RECT MASK 2 63.155 33.69 63.215 33.93 ;
      RECT MASK 2 63.595 33.69 63.655 33.93 ;
      RECT MASK 2 64.493 33.69 64.553 33.93 ;
      RECT MASK 2 64.933 33.69 64.993 33.93 ;
      RECT MASK 2 65.373 33.69 65.433 33.93 ;
      RECT MASK 2 65.813 33.69 65.873 33.93 ;
      RECT MASK 2 66.253 33.69 66.313 33.93 ;
      RECT MASK 2 66.693 33.69 66.753 33.93 ;
      RECT MASK 2 67.133 33.69 67.193 33.93 ;
      RECT MASK 2 67.573 33.69 67.633 33.93 ;
      RECT MASK 2 68.013 33.69 68.073 33.93 ;
      RECT MASK 2 68.453 33.69 68.513 33.93 ;
      RECT MASK 2 68.893 33.69 68.953 33.93 ;
      RECT MASK 2 69.333 33.69 69.393 33.93 ;
      RECT MASK 2 69.773 33.69 69.833 33.93 ;
      RECT MASK 2 70.213 33.69 70.273 33.93 ;
      RECT MASK 2 71.111 33.69 71.171 33.93 ;
      RECT MASK 2 71.551 33.69 71.611 33.93 ;
      RECT MASK 2 71.991 33.69 72.051 33.93 ;
      RECT MASK 2 72.431 33.69 72.491 33.93 ;
      RECT MASK 2 72.871 33.69 72.931 33.93 ;
      RECT MASK 2 73.311 33.69 73.371 33.93 ;
      RECT MASK 2 73.751 33.69 73.811 33.93 ;
      RECT MASK 2 74.191 33.69 74.251 33.93 ;
      RECT MASK 2 74.631 33.69 74.691 33.93 ;
      RECT MASK 2 75.071 33.69 75.131 33.93 ;
      RECT MASK 2 75.511 33.69 75.571 33.93 ;
      RECT MASK 2 75.951 33.69 76.011 33.93 ;
      RECT MASK 2 76.391 33.69 76.451 33.93 ;
      RECT MASK 2 76.831 33.69 76.891 33.93 ;
      RECT MASK 2 77.729 33.69 77.789 33.93 ;
      RECT MASK 2 78.169 33.69 78.229 33.93 ;
      RECT MASK 2 78.609 33.69 78.669 33.93 ;
      RECT MASK 2 79.049 33.69 79.109 33.93 ;
      RECT MASK 2 79.489 33.69 79.549 33.93 ;
      RECT MASK 2 79.929 33.69 79.989 33.93 ;
      RECT MASK 2 80.369 33.69 80.429 33.93 ;
      RECT MASK 2 80.809 33.69 80.869 33.93 ;
      RECT MASK 2 81.249 33.69 81.309 33.93 ;
      RECT MASK 2 81.689 33.69 81.749 33.93 ;
      RECT MASK 2 82.129 33.69 82.189 33.93 ;
      RECT MASK 2 83.449 33.69 83.509 33.93 ;
      RECT MASK 2 84.347 33.69 84.407 33.93 ;
      RECT MASK 2 84.787 33.69 84.847 33.93 ;
      RECT MASK 2 85.227 33.69 85.287 33.93 ;
      RECT MASK 2 85.667 33.69 85.727 33.93 ;
      RECT MASK 2 86.107 33.69 86.167 33.93 ;
      RECT MASK 2 86.547 33.69 86.607 33.93 ;
      RECT MASK 2 86.987 33.69 87.047 33.93 ;
      RECT MASK 2 87.427 33.69 87.487 33.93 ;
      RECT MASK 2 87.867 33.69 87.927 33.93 ;
      RECT MASK 2 88.307 33.69 88.367 33.93 ;
      RECT MASK 2 88.747 33.69 88.807 33.93 ;
      RECT MASK 2 89.187 33.69 89.247 33.93 ;
      RECT MASK 2 89.627 33.69 89.687 33.93 ;
      RECT MASK 2 90.067 33.69 90.127 33.93 ;
      RECT MASK 2 90.965 33.69 91.025 33.93 ;
      RECT MASK 2 91.405 33.69 91.465 33.93 ;
      RECT MASK 2 91.845 33.69 91.905 33.93 ;
      RECT MASK 2 92.285 33.69 92.345 33.93 ;
      RECT MASK 2 92.725 33.69 92.785 33.93 ;
      RECT MASK 2 93.165 33.69 93.225 33.93 ;
      RECT MASK 2 93.605 33.69 93.665 33.93 ;
      RECT MASK 2 94.045 33.69 94.105 33.93 ;
      RECT MASK 2 94.485 33.69 94.545 33.93 ;
      RECT MASK 2 94.925 33.69 94.985 33.93 ;
      RECT MASK 2 95.365 33.69 95.425 33.93 ;
      RECT MASK 2 95.805 33.69 95.865 33.93 ;
      RECT MASK 2 96.245 33.69 96.305 33.93 ;
      RECT MASK 2 96.685 33.69 96.745 33.93 ;
      RECT MASK 2 97.583 33.69 97.643 33.93 ;
      RECT MASK 2 98.023 33.69 98.083 33.93 ;
      RECT MASK 2 98.463 33.69 98.523 33.93 ;
      RECT MASK 2 98.903 33.69 98.963 33.93 ;
      RECT MASK 2 99.343 33.69 99.403 33.93 ;
      RECT MASK 2 99.783 33.69 99.843 33.93 ;
      RECT MASK 2 100.223 33.69 100.283 33.93 ;
      RECT MASK 2 100.663 33.69 100.723 33.93 ;
      RECT MASK 2 101.103 33.69 101.163 33.93 ;
      RECT MASK 2 101.543 33.69 101.603 33.93 ;
      RECT MASK 2 101.983 33.69 102.043 33.93 ;
      RECT MASK 2 102.423 33.69 102.483 33.93 ;
      RECT MASK 2 102.863 33.69 102.923 33.93 ;
      RECT MASK 2 103.303 33.69 103.363 33.93 ;
      RECT MASK 2 104.201 33.69 104.261 33.93 ;
      RECT MASK 2 104.641 33.69 104.701 33.93 ;
      RECT MASK 2 105.081 33.69 105.141 33.93 ;
      RECT MASK 2 105.521 33.69 105.581 33.93 ;
      RECT MASK 2 105.961 33.69 106.021 33.93 ;
      RECT MASK 2 106.401 33.69 106.461 33.93 ;
      RECT MASK 2 106.841 33.69 106.901 33.93 ;
      RECT MASK 2 107.281 33.69 107.341 33.93 ;
      RECT MASK 2 107.721 33.69 107.781 33.93 ;
      RECT MASK 2 108.161 33.69 108.221 33.93 ;
      RECT MASK 2 108.601 33.69 108.661 33.93 ;
      RECT MASK 2 109.041 33.69 109.101 33.93 ;
      RECT MASK 2 109.481 33.69 109.541 33.93 ;
      RECT MASK 2 109.921 33.69 109.981 33.93 ;
      RECT MASK 2 4.901 34.099 5.021 45.311 ;
      RECT MASK 2 5.341 34.099 5.461 45.311 ;
      RECT MASK 2 5.781 34.099 5.901 45.311 ;
      RECT MASK 2 6.221 34.099 6.341 45.311 ;
      RECT MASK 2 6.661 34.099 6.781 45.311 ;
      RECT MASK 2 7.101 34.099 7.221 45.311 ;
      RECT MASK 2 7.541 34.099 7.661 45.311 ;
      RECT MASK 2 7.981 34.099 8.101 45.311 ;
      RECT MASK 2 8.421 34.099 8.541 45.311 ;
      RECT MASK 2 8.861 34.099 8.981 45.311 ;
      RECT MASK 2 9.301 34.099 9.421 45.311 ;
      RECT MASK 2 9.741 34.099 9.861 45.311 ;
      RECT MASK 2 10.181 34.099 10.301 45.311 ;
      RECT MASK 2 10.621 34.099 10.741 45.311 ;
      RECT MASK 2 11.519 34.099 11.639 45.311 ;
      RECT MASK 2 11.959 34.099 12.079 45.311 ;
      RECT MASK 2 12.399 34.099 12.519 45.311 ;
      RECT MASK 2 12.839 34.099 12.959 45.311 ;
      RECT MASK 2 13.279 34.099 13.399 45.311 ;
      RECT MASK 2 13.719 34.099 13.839 45.311 ;
      RECT MASK 2 14.159 34.099 14.279 45.311 ;
      RECT MASK 2 14.599 34.099 14.719 45.311 ;
      RECT MASK 2 15.039 34.099 15.159 45.311 ;
      RECT MASK 2 15.479 34.099 15.599 45.311 ;
      RECT MASK 2 15.919 34.099 16.039 45.311 ;
      RECT MASK 2 16.359 34.099 16.479 45.311 ;
      RECT MASK 2 16.799 34.099 16.919 45.311 ;
      RECT MASK 2 17.239 34.099 17.359 45.311 ;
      RECT MASK 2 18.137 34.099 18.257 45.311 ;
      RECT MASK 2 18.577 34.099 18.697 45.311 ;
      RECT MASK 2 19.017 34.099 19.137 45.311 ;
      RECT MASK 2 19.457 34.099 19.577 45.311 ;
      RECT MASK 2 19.897 34.099 20.017 45.311 ;
      RECT MASK 2 20.337 34.099 20.457 45.311 ;
      RECT MASK 2 20.777 34.099 20.897 45.311 ;
      RECT MASK 2 21.217 34.099 21.337 45.311 ;
      RECT MASK 2 21.657 34.099 21.777 45.311 ;
      RECT MASK 2 22.097 34.099 22.217 45.311 ;
      RECT MASK 2 22.537 34.099 22.657 45.311 ;
      RECT MASK 2 22.977 34.099 23.097 45.311 ;
      RECT MASK 2 23.417 34.099 23.537 45.311 ;
      RECT MASK 2 23.857 34.099 23.977 45.311 ;
      RECT MASK 2 24.755 34.099 24.875 45.311 ;
      RECT MASK 2 25.195 34.099 25.315 45.311 ;
      RECT MASK 2 25.635 34.099 25.755 45.311 ;
      RECT MASK 2 26.075 34.099 26.195 45.311 ;
      RECT MASK 2 26.515 34.099 26.635 45.311 ;
      RECT MASK 2 26.955 34.099 27.075 45.311 ;
      RECT MASK 2 27.395 34.099 27.515 45.311 ;
      RECT MASK 2 27.835 34.099 27.955 45.311 ;
      RECT MASK 2 28.275 34.099 28.395 45.311 ;
      RECT MASK 2 28.715 34.099 28.835 45.311 ;
      RECT MASK 2 29.155 34.099 29.275 45.311 ;
      RECT MASK 2 29.595 34.099 29.715 45.311 ;
      RECT MASK 2 30.035 34.099 30.155 45.311 ;
      RECT MASK 2 30.475 34.099 30.595 45.311 ;
      RECT MASK 2 31.373 34.099 31.493 45.311 ;
      RECT MASK 2 31.813 34.099 31.933 45.311 ;
      RECT MASK 2 32.253 34.099 32.373 45.311 ;
      RECT MASK 2 32.693 34.099 32.813 45.311 ;
      RECT MASK 2 33.133 34.099 33.253 45.311 ;
      RECT MASK 2 33.573 34.099 33.693 45.311 ;
      RECT MASK 2 34.013 34.099 34.133 45.311 ;
      RECT MASK 2 34.453 34.099 34.573 45.311 ;
      RECT MASK 2 34.893 34.099 35.013 45.311 ;
      RECT MASK 2 35.333 34.099 35.453 45.311 ;
      RECT MASK 2 35.773 34.099 35.893 45.311 ;
      RECT MASK 2 36.213 34.099 36.333 45.311 ;
      RECT MASK 2 36.653 34.099 36.773 45.311 ;
      RECT MASK 2 37.093 34.099 37.213 45.311 ;
      RECT MASK 2 37.991 34.099 38.111 45.311 ;
      RECT MASK 2 38.431 34.099 38.551 45.311 ;
      RECT MASK 2 38.871 34.099 38.991 45.311 ;
      RECT MASK 2 39.311 34.099 39.431 45.311 ;
      RECT MASK 2 39.751 34.099 39.871 45.311 ;
      RECT MASK 2 40.191 34.099 40.311 45.311 ;
      RECT MASK 2 40.631 34.099 40.751 45.311 ;
      RECT MASK 2 41.071 34.099 41.191 45.311 ;
      RECT MASK 2 41.511 34.099 41.631 45.311 ;
      RECT MASK 2 41.951 34.099 42.071 45.311 ;
      RECT MASK 2 42.391 34.099 42.511 45.311 ;
      RECT MASK 2 42.831 34.099 42.951 45.311 ;
      RECT MASK 2 43.271 34.099 43.391 45.311 ;
      RECT MASK 2 43.711 34.099 43.831 45.311 ;
      RECT MASK 2 44.609 34.099 44.729 45.311 ;
      RECT MASK 2 45.049 34.099 45.169 45.311 ;
      RECT MASK 2 45.489 34.099 45.609 45.311 ;
      RECT MASK 2 45.929 34.099 46.049 45.311 ;
      RECT MASK 2 46.369 34.099 46.489 45.311 ;
      RECT MASK 2 46.809 34.099 46.929 45.311 ;
      RECT MASK 2 47.249 34.099 47.369 45.311 ;
      RECT MASK 2 47.689 34.099 47.809 45.311 ;
      RECT MASK 2 48.129 34.099 48.249 45.311 ;
      RECT MASK 2 48.569 34.099 48.689 45.311 ;
      RECT MASK 2 49.009 34.099 49.129 45.311 ;
      RECT MASK 2 49.449 34.099 49.569 45.311 ;
      RECT MASK 2 49.889 34.099 50.009 45.311 ;
      RECT MASK 2 50.329 34.099 50.449 45.311 ;
      RECT MASK 2 51.227 34.099 51.347 45.311 ;
      RECT MASK 2 51.667 34.099 51.787 45.311 ;
      RECT MASK 2 52.107 34.099 52.227 45.311 ;
      RECT MASK 2 52.547 34.099 52.667 45.311 ;
      RECT MASK 2 52.987 34.099 53.107 45.311 ;
      RECT MASK 2 53.427 34.099 53.547 45.311 ;
      RECT MASK 2 53.867 34.099 53.987 45.311 ;
      RECT MASK 2 54.307 34.099 54.427 45.311 ;
      RECT MASK 2 54.747 34.099 54.867 45.311 ;
      RECT MASK 2 55.187 34.099 55.307 45.311 ;
      RECT MASK 2 55.627 34.099 55.747 45.311 ;
      RECT MASK 2 56.067 34.099 56.187 45.311 ;
      RECT MASK 2 56.507 34.099 56.627 45.311 ;
      RECT MASK 2 56.947 34.099 57.067 45.311 ;
      RECT MASK 2 57.845 34.099 57.965 45.311 ;
      RECT MASK 2 58.285 34.099 58.405 45.311 ;
      RECT MASK 2 58.725 34.099 58.845 45.311 ;
      RECT MASK 2 59.165 34.099 59.285 45.311 ;
      RECT MASK 2 59.605 34.099 59.725 45.311 ;
      RECT MASK 2 60.045 34.099 60.165 45.311 ;
      RECT MASK 2 60.485 34.099 60.605 45.311 ;
      RECT MASK 2 60.925 34.099 61.045 45.311 ;
      RECT MASK 2 61.365 34.099 61.485 45.311 ;
      RECT MASK 2 61.805 34.099 61.925 45.311 ;
      RECT MASK 2 62.245 34.099 62.365 45.311 ;
      RECT MASK 2 62.685 34.099 62.805 45.311 ;
      RECT MASK 2 63.125 34.099 63.245 45.311 ;
      RECT MASK 2 63.565 34.099 63.685 45.311 ;
      RECT MASK 2 64.463 34.099 64.583 45.311 ;
      RECT MASK 2 64.903 34.099 65.023 45.311 ;
      RECT MASK 2 65.343 34.099 65.463 45.311 ;
      RECT MASK 2 65.783 34.099 65.903 45.311 ;
      RECT MASK 2 66.223 34.099 66.343 45.311 ;
      RECT MASK 2 66.663 34.099 66.783 45.311 ;
      RECT MASK 2 67.103 34.099 67.223 45.311 ;
      RECT MASK 2 67.543 34.099 67.663 45.311 ;
      RECT MASK 2 67.983 34.099 68.103 45.311 ;
      RECT MASK 2 68.423 34.099 68.543 45.311 ;
      RECT MASK 2 68.863 34.099 68.983 45.311 ;
      RECT MASK 2 69.303 34.099 69.423 45.311 ;
      RECT MASK 2 69.743 34.099 69.863 45.311 ;
      RECT MASK 2 70.183 34.099 70.303 45.311 ;
      RECT MASK 2 71.081 34.099 71.201 45.311 ;
      RECT MASK 2 71.521 34.099 71.641 45.311 ;
      RECT MASK 2 71.961 34.099 72.081 45.311 ;
      RECT MASK 2 72.401 34.099 72.521 45.311 ;
      RECT MASK 2 72.841 34.099 72.961 45.311 ;
      RECT MASK 2 73.281 34.099 73.401 45.311 ;
      RECT MASK 2 73.721 34.099 73.841 45.311 ;
      RECT MASK 2 74.161 34.099 74.281 45.311 ;
      RECT MASK 2 74.601 34.099 74.721 45.311 ;
      RECT MASK 2 75.041 34.099 75.161 45.311 ;
      RECT MASK 2 75.481 34.099 75.601 45.311 ;
      RECT MASK 2 75.921 34.099 76.041 45.311 ;
      RECT MASK 2 76.361 34.099 76.481 45.311 ;
      RECT MASK 2 76.801 34.099 76.921 45.311 ;
      RECT MASK 2 77.699 34.099 77.819 45.311 ;
      RECT MASK 2 78.139 34.099 78.259 45.311 ;
      RECT MASK 2 78.579 34.099 78.699 45.311 ;
      RECT MASK 2 79.019 34.099 79.139 45.311 ;
      RECT MASK 2 79.459 34.099 79.579 45.311 ;
      RECT MASK 2 79.899 34.099 80.019 45.311 ;
      RECT MASK 2 80.339 34.099 80.459 45.311 ;
      RECT MASK 2 80.779 34.099 80.899 45.311 ;
      RECT MASK 2 81.219 34.099 81.339 45.311 ;
      RECT MASK 2 81.659 34.099 81.779 45.311 ;
      RECT MASK 2 82.099 34.099 82.219 45.311 ;
      RECT MASK 2 82.539 34.099 82.659 45.311 ;
      RECT MASK 2 82.979 34.099 83.099 45.311 ;
      RECT MASK 2 83.419 34.099 83.539 45.311 ;
      RECT MASK 2 84.317 34.099 84.437 45.311 ;
      RECT MASK 2 84.757 34.099 84.877 45.311 ;
      RECT MASK 2 85.197 34.099 85.317 45.311 ;
      RECT MASK 2 85.637 34.099 85.757 45.311 ;
      RECT MASK 2 86.077 34.099 86.197 45.311 ;
      RECT MASK 2 86.517 34.099 86.637 45.311 ;
      RECT MASK 2 86.957 34.099 87.077 45.311 ;
      RECT MASK 2 87.397 34.099 87.517 45.311 ;
      RECT MASK 2 87.837 34.099 87.957 45.311 ;
      RECT MASK 2 88.277 34.099 88.397 45.311 ;
      RECT MASK 2 88.717 34.099 88.837 45.311 ;
      RECT MASK 2 89.157 34.099 89.277 45.311 ;
      RECT MASK 2 89.597 34.099 89.717 45.311 ;
      RECT MASK 2 90.037 34.099 90.157 45.311 ;
      RECT MASK 2 90.935 34.099 91.055 45.311 ;
      RECT MASK 2 91.375 34.099 91.495 45.311 ;
      RECT MASK 2 91.815 34.099 91.935 45.311 ;
      RECT MASK 2 92.255 34.099 92.375 45.311 ;
      RECT MASK 2 92.695 34.099 92.815 45.311 ;
      RECT MASK 2 93.135 34.099 93.255 45.311 ;
      RECT MASK 2 93.575 34.099 93.695 45.311 ;
      RECT MASK 2 94.015 34.099 94.135 45.311 ;
      RECT MASK 2 94.455 34.099 94.575 45.311 ;
      RECT MASK 2 94.895 34.099 95.015 45.311 ;
      RECT MASK 2 95.335 34.099 95.455 45.311 ;
      RECT MASK 2 95.775 34.099 95.895 45.311 ;
      RECT MASK 2 96.215 34.099 96.335 45.311 ;
      RECT MASK 2 96.655 34.099 96.775 45.311 ;
      RECT MASK 2 97.553 34.099 97.673 45.311 ;
      RECT MASK 2 97.993 34.099 98.113 45.311 ;
      RECT MASK 2 98.433 34.099 98.553 45.311 ;
      RECT MASK 2 98.873 34.099 98.993 45.311 ;
      RECT MASK 2 99.313 34.099 99.433 45.311 ;
      RECT MASK 2 99.753 34.099 99.873 45.311 ;
      RECT MASK 2 100.193 34.099 100.313 45.311 ;
      RECT MASK 2 100.633 34.099 100.753 45.311 ;
      RECT MASK 2 101.073 34.099 101.193 45.311 ;
      RECT MASK 2 101.513 34.099 101.633 45.311 ;
      RECT MASK 2 101.953 34.099 102.073 45.311 ;
      RECT MASK 2 102.393 34.099 102.513 45.311 ;
      RECT MASK 2 102.833 34.099 102.953 45.311 ;
      RECT MASK 2 103.273 34.099 103.393 45.311 ;
      RECT MASK 2 104.171 34.099 104.291 45.311 ;
      RECT MASK 2 104.611 34.099 104.731 45.311 ;
      RECT MASK 2 105.051 34.099 105.171 45.311 ;
      RECT MASK 2 105.491 34.099 105.611 45.311 ;
      RECT MASK 2 105.931 34.099 106.051 45.311 ;
      RECT MASK 2 106.371 34.099 106.491 45.311 ;
      RECT MASK 2 106.811 34.099 106.931 45.311 ;
      RECT MASK 2 107.251 34.099 107.371 45.311 ;
      RECT MASK 2 107.691 34.099 107.811 45.311 ;
      RECT MASK 2 108.131 34.099 108.251 45.311 ;
      RECT MASK 2 108.571 34.099 108.691 45.311 ;
      RECT MASK 2 109.011 34.099 109.131 45.311 ;
      RECT MASK 2 109.451 34.099 109.571 45.311 ;
      RECT MASK 2 109.891 34.099 110.011 45.311 ;
      RECT MASK 2 112.5865 34.729 112.7065 35.819 ;
      RECT MASK 2 113.0265 34.729 113.1465 35.819 ;
      RECT MASK 2 113.4665 34.729 113.5865 35.819 ;
      RECT MASK 2 113.9065 34.729 114.0265 35.819 ;
      RECT MASK 2 114.3465 34.729 114.4665 35.819 ;
      RECT MASK 2 114.7865 34.729 114.9065 35.819 ;
      RECT MASK 2 115.2265 34.729 115.3465 35.819 ;
      RECT MASK 2 115.6665 34.729 115.7865 35.819 ;
      RECT MASK 2 116.1065 34.729 116.2265 35.819 ;
      RECT MASK 2 116.5465 34.729 116.6665 35.819 ;
      RECT MASK 2 117.4265 34.729 117.5465 35.819 ;
      RECT MASK 2 117.8665 34.729 117.9865 35.819 ;
      RECT MASK 2 118.3065 34.729 118.4265 35.819 ;
      RECT MASK 2 118.7465 34.729 118.8665 35.819 ;
      RECT MASK 2 119.1865 34.729 119.3065 35.819 ;
      RECT MASK 2 119.6265 34.729 119.7465 35.819 ;
      RECT MASK 2 120.0665 34.729 120.1865 35.819 ;
      RECT MASK 2 120.5065 34.729 120.6265 35.819 ;
      RECT MASK 2 120.9465 34.729 121.0665 35.819 ;
      RECT MASK 2 121.3865 34.729 121.5065 35.819 ;
      RECT MASK 2 121.8265 34.729 121.9465 35.819 ;
      RECT MASK 2 122.2665 34.729 122.3865 35.819 ;
      RECT MASK 2 122.7065 34.729 122.8265 35.819 ;
      RECT MASK 2 123.1465 34.729 123.2665 35.819 ;
      RECT MASK 2 123.5865 34.729 123.7065 35.819 ;
      RECT MASK 2 112.5865 36.079 112.7065 37.169 ;
      RECT MASK 2 113.0265 36.079 113.1465 37.169 ;
      RECT MASK 2 113.4665 36.079 113.5865 37.169 ;
      RECT MASK 2 113.9065 36.079 114.0265 37.169 ;
      RECT MASK 2 114.3465 36.079 114.4665 37.169 ;
      RECT MASK 2 114.7865 36.079 114.9065 37.169 ;
      RECT MASK 2 115.2265 36.079 115.3465 37.169 ;
      RECT MASK 2 115.6665 36.079 115.7865 37.169 ;
      RECT MASK 2 116.1065 36.079 116.2265 37.169 ;
      RECT MASK 2 116.5465 36.079 116.6665 37.169 ;
      RECT MASK 2 117.4265 36.079 117.5465 37.169 ;
      RECT MASK 2 117.8665 36.079 117.9865 37.169 ;
      RECT MASK 2 118.3065 36.079 118.4265 37.169 ;
      RECT MASK 2 118.7465 36.079 118.8665 37.169 ;
      RECT MASK 2 119.1865 36.079 119.3065 37.169 ;
      RECT MASK 2 119.6265 36.079 119.7465 37.169 ;
      RECT MASK 2 120.0665 36.079 120.1865 37.169 ;
      RECT MASK 2 120.5065 36.079 120.6265 37.169 ;
      RECT MASK 2 120.9465 36.079 121.0665 37.169 ;
      RECT MASK 2 121.3865 36.079 121.5065 37.169 ;
      RECT MASK 2 121.8265 36.079 121.9465 37.169 ;
      RECT MASK 2 122.2665 36.079 122.3865 37.169 ;
      RECT MASK 2 122.7065 36.079 122.8265 37.169 ;
      RECT MASK 2 123.1465 36.079 123.2665 37.169 ;
      RECT MASK 2 123.5865 36.079 123.7065 37.169 ;
      RECT MASK 2 112.5865 37.429 112.7065 38.519 ;
      RECT MASK 2 113.0265 37.429 113.1465 38.519 ;
      RECT MASK 2 113.4665 37.429 113.5865 38.519 ;
      RECT MASK 2 113.9065 37.429 114.0265 38.519 ;
      RECT MASK 2 114.3465 37.429 114.4665 38.519 ;
      RECT MASK 2 114.7865 37.429 114.9065 38.519 ;
      RECT MASK 2 115.2265 37.429 115.3465 38.519 ;
      RECT MASK 2 115.6665 37.429 115.7865 38.519 ;
      RECT MASK 2 116.1065 37.429 116.2265 38.519 ;
      RECT MASK 2 116.5465 37.429 116.6665 38.519 ;
      RECT MASK 2 117.4265 37.429 117.5465 38.519 ;
      RECT MASK 2 117.8665 37.429 117.9865 38.519 ;
      RECT MASK 2 118.3065 37.429 118.4265 38.519 ;
      RECT MASK 2 118.7465 37.429 118.8665 38.519 ;
      RECT MASK 2 119.1865 37.429 119.3065 38.519 ;
      RECT MASK 2 119.6265 37.429 119.7465 38.519 ;
      RECT MASK 2 120.0665 37.429 120.1865 38.519 ;
      RECT MASK 2 120.5065 37.429 120.6265 38.519 ;
      RECT MASK 2 120.9465 37.429 121.0665 38.519 ;
      RECT MASK 2 121.3865 37.429 121.5065 38.519 ;
      RECT MASK 2 121.8265 37.429 121.9465 38.519 ;
      RECT MASK 2 122.2665 37.429 122.3865 38.519 ;
      RECT MASK 2 122.7065 37.429 122.8265 38.519 ;
      RECT MASK 2 123.1465 37.429 123.2665 38.519 ;
      RECT MASK 2 123.5865 37.429 123.7065 38.519 ;
      RECT MASK 2 112.5865 38.779 112.7065 40.619 ;
      RECT MASK 2 113.0265 38.779 113.1465 40.619 ;
      RECT MASK 2 113.4665 38.779 113.5865 40.619 ;
      RECT MASK 2 113.9065 38.779 114.0265 40.619 ;
      RECT MASK 2 114.3465 38.779 114.4665 40.619 ;
      RECT MASK 2 114.7865 38.779 114.9065 40.619 ;
      RECT MASK 2 115.2265 38.779 115.3465 40.619 ;
      RECT MASK 2 115.6665 38.779 115.7865 40.619 ;
      RECT MASK 2 116.1065 38.779 116.2265 40.619 ;
      RECT MASK 2 116.5465 38.779 116.6665 40.619 ;
      RECT MASK 2 117.4265 38.779 117.5465 40.619 ;
      RECT MASK 2 117.8665 38.779 117.9865 40.619 ;
      RECT MASK 2 118.3065 38.779 118.4265 40.619 ;
      RECT MASK 2 118.7465 38.779 118.8665 40.619 ;
      RECT MASK 2 119.1865 38.779 119.3065 40.619 ;
      RECT MASK 2 119.6265 38.779 119.7465 40.619 ;
      RECT MASK 2 120.0665 38.779 120.1865 40.619 ;
      RECT MASK 2 120.5065 38.779 120.6265 40.619 ;
      RECT MASK 2 120.9465 38.779 121.0665 40.619 ;
      RECT MASK 2 121.3865 38.779 121.5065 40.619 ;
      RECT MASK 2 121.8265 38.779 121.9465 40.619 ;
      RECT MASK 2 122.2665 38.779 122.3865 40.619 ;
      RECT MASK 2 122.7065 38.779 122.8265 40.619 ;
      RECT MASK 2 123.1465 38.779 123.2665 40.619 ;
      RECT MASK 2 123.5865 38.779 123.7065 40.619 ;
      RECT MASK 2 112.5865 40.879 112.7065 41.939 ;
      RECT MASK 2 113.0265 40.879 113.1465 41.939 ;
      RECT MASK 2 113.4665 40.879 113.5865 41.939 ;
      RECT MASK 2 113.9065 40.879 114.0265 41.939 ;
      RECT MASK 2 114.3465 40.879 114.4665 41.939 ;
      RECT MASK 2 114.7865 40.879 114.9065 41.939 ;
      RECT MASK 2 115.2265 40.879 115.3465 41.939 ;
      RECT MASK 2 115.6665 40.879 115.7865 41.939 ;
      RECT MASK 2 116.1065 40.879 116.2265 41.939 ;
      RECT MASK 2 116.5465 40.879 116.6665 41.939 ;
      RECT MASK 2 117.4265 40.879 117.5465 41.939 ;
      RECT MASK 2 117.8665 40.879 117.9865 41.939 ;
      RECT MASK 2 118.3065 40.879 118.4265 41.939 ;
      RECT MASK 2 118.7465 40.879 118.8665 41.939 ;
      RECT MASK 2 119.1865 40.879 119.3065 41.939 ;
      RECT MASK 2 119.6265 40.879 119.7465 41.939 ;
      RECT MASK 2 120.0665 40.879 120.1865 41.939 ;
      RECT MASK 2 120.5065 40.879 120.6265 41.939 ;
      RECT MASK 2 120.9465 40.879 121.0665 41.939 ;
      RECT MASK 2 121.3865 40.879 121.5065 41.939 ;
      RECT MASK 2 121.8265 40.879 121.9465 41.939 ;
      RECT MASK 2 122.2665 40.879 122.3865 41.939 ;
      RECT MASK 2 122.7065 40.879 122.8265 41.939 ;
      RECT MASK 2 123.1465 40.879 123.2665 41.939 ;
      RECT MASK 2 123.5865 40.879 123.7065 41.939 ;
      RECT MASK 2 112.5865 42.199 112.7065 43.289 ;
      RECT MASK 2 113.0265 42.199 113.1465 43.289 ;
      RECT MASK 2 113.4665 42.199 113.5865 43.289 ;
      RECT MASK 2 113.9065 42.199 114.0265 43.289 ;
      RECT MASK 2 114.3465 42.199 114.4665 43.289 ;
      RECT MASK 2 114.7865 42.199 114.9065 43.289 ;
      RECT MASK 2 115.2265 42.199 115.3465 43.289 ;
      RECT MASK 2 115.6665 42.199 115.7865 43.289 ;
      RECT MASK 2 116.1065 42.199 116.2265 43.289 ;
      RECT MASK 2 116.5465 42.199 116.6665 43.289 ;
      RECT MASK 2 117.4265 42.199 117.5465 43.289 ;
      RECT MASK 2 117.8665 42.199 117.9865 43.289 ;
      RECT MASK 2 118.3065 42.199 118.4265 43.289 ;
      RECT MASK 2 118.7465 42.199 118.8665 43.289 ;
      RECT MASK 2 119.1865 42.199 119.3065 43.289 ;
      RECT MASK 2 119.6265 42.199 119.7465 43.289 ;
      RECT MASK 2 120.0665 42.199 120.1865 43.289 ;
      RECT MASK 2 120.5065 42.199 120.6265 43.289 ;
      RECT MASK 2 120.9465 42.199 121.0665 43.289 ;
      RECT MASK 2 121.3865 42.199 121.5065 43.289 ;
      RECT MASK 2 121.8265 42.199 121.9465 43.289 ;
      RECT MASK 2 122.2665 42.199 122.3865 43.289 ;
      RECT MASK 2 122.7065 42.199 122.8265 43.289 ;
      RECT MASK 2 123.1465 42.199 123.2665 43.289 ;
      RECT MASK 2 123.5865 42.199 123.7065 43.289 ;
      RECT MASK 2 112.5865 43.549 112.7065 44.639 ;
      RECT MASK 2 113.0265 43.549 113.1465 44.639 ;
      RECT MASK 2 113.4665 43.549 113.5865 44.639 ;
      RECT MASK 2 113.9065 43.549 114.0265 44.639 ;
      RECT MASK 2 114.3465 43.549 114.4665 44.639 ;
      RECT MASK 2 114.7865 43.549 114.9065 44.639 ;
      RECT MASK 2 115.2265 43.549 115.3465 44.639 ;
      RECT MASK 2 115.6665 43.549 115.7865 44.639 ;
      RECT MASK 2 116.1065 43.549 116.2265 44.639 ;
      RECT MASK 2 116.5465 43.549 116.6665 44.639 ;
      RECT MASK 2 117.4265 43.549 117.5465 44.639 ;
      RECT MASK 2 117.8665 43.549 117.9865 44.639 ;
      RECT MASK 2 118.3065 43.549 118.4265 44.639 ;
      RECT MASK 2 118.7465 43.549 118.8665 44.639 ;
      RECT MASK 2 119.1865 43.549 119.3065 44.639 ;
      RECT MASK 2 119.6265 43.549 119.7465 44.639 ;
      RECT MASK 2 120.0665 43.549 120.1865 44.639 ;
      RECT MASK 2 120.5065 43.549 120.6265 44.639 ;
      RECT MASK 2 120.9465 43.549 121.0665 44.639 ;
      RECT MASK 2 121.3865 43.549 121.5065 44.639 ;
      RECT MASK 2 121.8265 43.549 121.9465 44.639 ;
      RECT MASK 2 122.2665 43.549 122.3865 44.639 ;
      RECT MASK 2 122.7065 43.549 122.8265 44.639 ;
      RECT MASK 2 123.1465 43.549 123.2665 44.639 ;
      RECT MASK 2 123.5865 43.549 123.7065 44.639 ;
      RECT MASK 2 112.5865 44.899 112.7065 46.709 ;
      RECT MASK 2 113.0265 44.899 113.1465 46.709 ;
      RECT MASK 2 113.4665 44.899 113.5865 46.709 ;
      RECT MASK 2 113.9065 44.899 114.0265 46.709 ;
      RECT MASK 2 114.3465 44.899 114.4665 46.709 ;
      RECT MASK 2 114.7865 44.899 114.9065 46.709 ;
      RECT MASK 2 115.2265 44.899 115.3465 46.709 ;
      RECT MASK 2 115.6665 44.899 115.7865 46.709 ;
      RECT MASK 2 116.1065 44.899 116.2265 46.709 ;
      RECT MASK 2 116.5465 44.899 116.6665 46.709 ;
      RECT MASK 2 117.4265 44.899 117.5465 46.709 ;
      RECT MASK 2 117.8665 44.899 117.9865 46.709 ;
      RECT MASK 2 118.3065 44.899 118.4265 46.709 ;
      RECT MASK 2 118.7465 44.899 118.8665 46.709 ;
      RECT MASK 2 119.1865 44.899 119.3065 46.709 ;
      RECT MASK 2 119.6265 44.899 119.7465 46.709 ;
      RECT MASK 2 120.0665 44.899 120.1865 46.709 ;
      RECT MASK 2 120.5065 44.899 120.6265 46.709 ;
      RECT MASK 2 120.9465 44.899 121.0665 46.709 ;
      RECT MASK 2 121.3865 44.899 121.5065 46.709 ;
      RECT MASK 2 121.8265 44.899 121.9465 46.709 ;
      RECT MASK 2 122.2665 44.899 122.3865 46.709 ;
      RECT MASK 2 122.7065 44.899 122.8265 46.709 ;
      RECT MASK 2 123.1465 44.899 123.2665 46.709 ;
      RECT MASK 2 123.5865 44.899 123.7065 46.709 ;
      RECT MASK 2 4.931 45.48 4.991 45.72 ;
      RECT MASK 2 5.371 45.48 5.431 45.72 ;
      RECT MASK 2 5.811 45.48 5.871 45.72 ;
      RECT MASK 2 6.251 45.48 6.311 45.72 ;
      RECT MASK 2 6.691 45.48 6.751 45.72 ;
      RECT MASK 2 7.131 45.48 7.191 45.72 ;
      RECT MASK 2 7.571 45.48 7.631 45.72 ;
      RECT MASK 2 8.011 45.48 8.071 45.72 ;
      RECT MASK 2 8.451 45.48 8.511 45.72 ;
      RECT MASK 2 8.891 45.48 8.951 45.72 ;
      RECT MASK 2 9.331 45.48 9.391 45.72 ;
      RECT MASK 2 9.771 45.48 9.831 45.72 ;
      RECT MASK 2 10.211 45.48 10.271 45.72 ;
      RECT MASK 2 10.651 45.48 10.711 45.72 ;
      RECT MASK 2 11.549 45.48 11.609 45.72 ;
      RECT MASK 2 11.989 45.48 12.049 45.72 ;
      RECT MASK 2 12.429 45.48 12.489 45.72 ;
      RECT MASK 2 12.869 45.48 12.929 45.72 ;
      RECT MASK 2 13.309 45.48 13.369 45.72 ;
      RECT MASK 2 13.749 45.48 13.809 45.72 ;
      RECT MASK 2 14.189 45.48 14.249 45.72 ;
      RECT MASK 2 14.629 45.48 14.689 45.72 ;
      RECT MASK 2 15.069 45.48 15.129 45.72 ;
      RECT MASK 2 15.509 45.48 15.569 45.72 ;
      RECT MASK 2 15.949 45.48 16.009 45.72 ;
      RECT MASK 2 16.389 45.48 16.449 45.72 ;
      RECT MASK 2 16.829 45.48 16.889 45.72 ;
      RECT MASK 2 17.269 45.48 17.329 45.72 ;
      RECT MASK 2 18.167 45.48 18.227 45.72 ;
      RECT MASK 2 18.607 45.48 18.667 45.72 ;
      RECT MASK 2 19.047 45.48 19.107 45.72 ;
      RECT MASK 2 19.487 45.48 19.547 45.72 ;
      RECT MASK 2 19.927 45.48 19.987 45.72 ;
      RECT MASK 2 20.367 45.48 20.427 45.72 ;
      RECT MASK 2 20.807 45.48 20.867 45.72 ;
      RECT MASK 2 21.247 45.48 21.307 45.72 ;
      RECT MASK 2 21.687 45.48 21.747 45.72 ;
      RECT MASK 2 22.127 45.48 22.187 45.72 ;
      RECT MASK 2 22.567 45.48 22.627 45.72 ;
      RECT MASK 2 23.007 45.48 23.067 45.72 ;
      RECT MASK 2 23.447 45.48 23.507 45.72 ;
      RECT MASK 2 23.887 45.48 23.947 45.72 ;
      RECT MASK 2 24.785 45.48 24.845 45.72 ;
      RECT MASK 2 25.225 45.48 25.285 45.72 ;
      RECT MASK 2 25.665 45.48 25.725 45.72 ;
      RECT MASK 2 26.105 45.48 26.165 45.72 ;
      RECT MASK 2 26.545 45.48 26.605 45.72 ;
      RECT MASK 2 26.985 45.48 27.045 45.72 ;
      RECT MASK 2 27.425 45.48 27.485 45.72 ;
      RECT MASK 2 27.865 45.48 27.925 45.72 ;
      RECT MASK 2 28.305 45.48 28.365 45.72 ;
      RECT MASK 2 28.745 45.48 28.805 45.72 ;
      RECT MASK 2 29.185 45.48 29.245 45.72 ;
      RECT MASK 2 29.625 45.48 29.685 45.72 ;
      RECT MASK 2 30.065 45.48 30.125 45.72 ;
      RECT MASK 2 30.505 45.48 30.565 45.72 ;
      RECT MASK 2 31.403 45.48 31.463 45.72 ;
      RECT MASK 2 31.843 45.48 31.903 45.72 ;
      RECT MASK 2 32.283 45.48 32.343 45.72 ;
      RECT MASK 2 32.723 45.48 32.783 45.72 ;
      RECT MASK 2 33.163 45.48 33.223 45.72 ;
      RECT MASK 2 33.603 45.48 33.663 45.72 ;
      RECT MASK 2 34.043 45.48 34.103 45.72 ;
      RECT MASK 2 34.483 45.48 34.543 45.72 ;
      RECT MASK 2 34.923 45.48 34.983 45.72 ;
      RECT MASK 2 35.363 45.48 35.423 45.72 ;
      RECT MASK 2 35.803 45.48 35.863 45.72 ;
      RECT MASK 2 36.243 45.48 36.303 45.72 ;
      RECT MASK 2 36.683 45.48 36.743 45.72 ;
      RECT MASK 2 37.123 45.48 37.183 45.72 ;
      RECT MASK 2 38.021 45.48 38.081 45.72 ;
      RECT MASK 2 38.461 45.48 38.521 45.72 ;
      RECT MASK 2 38.901 45.48 38.961 45.72 ;
      RECT MASK 2 39.341 45.48 39.401 45.72 ;
      RECT MASK 2 39.781 45.48 39.841 45.72 ;
      RECT MASK 2 40.221 45.48 40.281 45.72 ;
      RECT MASK 2 40.661 45.48 40.721 45.72 ;
      RECT MASK 2 41.101 45.48 41.161 45.72 ;
      RECT MASK 2 41.541 45.48 41.601 45.72 ;
      RECT MASK 2 42.861 45.48 42.921 45.72 ;
      RECT MASK 2 43.301 45.48 43.361 45.72 ;
      RECT MASK 2 43.741 45.48 43.801 45.72 ;
      RECT MASK 2 44.639 45.48 44.699 45.72 ;
      RECT MASK 2 45.079 45.48 45.139 45.72 ;
      RECT MASK 2 45.519 45.48 45.579 45.72 ;
      RECT MASK 2 45.959 45.48 46.019 45.72 ;
      RECT MASK 2 46.399 45.48 46.459 45.72 ;
      RECT MASK 2 46.839 45.48 46.899 45.72 ;
      RECT MASK 2 47.279 45.48 47.339 45.72 ;
      RECT MASK 2 47.719 45.48 47.779 45.72 ;
      RECT MASK 2 48.159 45.48 48.219 45.72 ;
      RECT MASK 2 48.599 45.48 48.659 45.72 ;
      RECT MASK 2 49.039 45.48 49.099 45.72 ;
      RECT MASK 2 49.479 45.48 49.539 45.72 ;
      RECT MASK 2 49.919 45.48 49.979 45.72 ;
      RECT MASK 2 50.359 45.48 50.419 45.72 ;
      RECT MASK 2 51.257 45.48 51.317 45.72 ;
      RECT MASK 2 51.697 45.48 51.757 45.72 ;
      RECT MASK 2 52.137 45.48 52.197 45.72 ;
      RECT MASK 2 52.577 45.48 52.637 45.72 ;
      RECT MASK 2 53.017 45.48 53.077 45.72 ;
      RECT MASK 2 53.457 45.48 53.517 45.72 ;
      RECT MASK 2 53.897 45.48 53.957 45.72 ;
      RECT MASK 2 54.337 45.48 54.397 45.72 ;
      RECT MASK 2 54.777 45.48 54.837 45.72 ;
      RECT MASK 2 55.217 45.48 55.277 45.72 ;
      RECT MASK 2 55.657 45.48 55.717 45.72 ;
      RECT MASK 2 56.097 45.48 56.157 45.72 ;
      RECT MASK 2 56.537 45.48 56.597 45.72 ;
      RECT MASK 2 56.977 45.48 57.037 45.72 ;
      RECT MASK 2 57.875 45.48 57.935 45.72 ;
      RECT MASK 2 58.315 45.48 58.375 45.72 ;
      RECT MASK 2 58.755 45.48 58.815 45.72 ;
      RECT MASK 2 59.195 45.48 59.255 45.72 ;
      RECT MASK 2 59.635 45.48 59.695 45.72 ;
      RECT MASK 2 60.075 45.48 60.135 45.72 ;
      RECT MASK 2 60.515 45.48 60.575 45.72 ;
      RECT MASK 2 60.955 45.48 61.015 45.72 ;
      RECT MASK 2 61.395 45.48 61.455 45.72 ;
      RECT MASK 2 61.835 45.48 61.895 45.72 ;
      RECT MASK 2 62.275 45.48 62.335 45.72 ;
      RECT MASK 2 62.715 45.48 62.775 45.72 ;
      RECT MASK 2 63.155 45.48 63.215 45.72 ;
      RECT MASK 2 63.595 45.48 63.655 45.72 ;
      RECT MASK 2 64.493 45.48 64.553 45.72 ;
      RECT MASK 2 64.933 45.48 64.993 45.72 ;
      RECT MASK 2 65.373 45.48 65.433 45.72 ;
      RECT MASK 2 65.813 45.48 65.873 45.72 ;
      RECT MASK 2 66.253 45.48 66.313 45.72 ;
      RECT MASK 2 66.693 45.48 66.753 45.72 ;
      RECT MASK 2 67.133 45.48 67.193 45.72 ;
      RECT MASK 2 67.573 45.48 67.633 45.72 ;
      RECT MASK 2 68.013 45.48 68.073 45.72 ;
      RECT MASK 2 68.453 45.48 68.513 45.72 ;
      RECT MASK 2 68.893 45.48 68.953 45.72 ;
      RECT MASK 2 69.333 45.48 69.393 45.72 ;
      RECT MASK 2 69.773 45.48 69.833 45.72 ;
      RECT MASK 2 70.213 45.48 70.273 45.72 ;
      RECT MASK 2 71.111 45.48 71.171 45.72 ;
      RECT MASK 2 71.551 45.48 71.611 45.72 ;
      RECT MASK 2 71.991 45.48 72.051 45.72 ;
      RECT MASK 2 72.431 45.48 72.491 45.72 ;
      RECT MASK 2 72.871 45.48 72.931 45.72 ;
      RECT MASK 2 73.311 45.48 73.371 45.72 ;
      RECT MASK 2 73.751 45.48 73.811 45.72 ;
      RECT MASK 2 74.191 45.48 74.251 45.72 ;
      RECT MASK 2 74.631 45.48 74.691 45.72 ;
      RECT MASK 2 75.071 45.48 75.131 45.72 ;
      RECT MASK 2 75.511 45.48 75.571 45.72 ;
      RECT MASK 2 75.951 45.48 76.011 45.72 ;
      RECT MASK 2 76.391 45.48 76.451 45.72 ;
      RECT MASK 2 76.831 45.48 76.891 45.72 ;
      RECT MASK 2 77.729 45.48 77.789 45.72 ;
      RECT MASK 2 78.169 45.48 78.229 45.72 ;
      RECT MASK 2 78.609 45.48 78.669 45.72 ;
      RECT MASK 2 79.049 45.48 79.109 45.72 ;
      RECT MASK 2 79.489 45.48 79.549 45.72 ;
      RECT MASK 2 79.929 45.48 79.989 45.72 ;
      RECT MASK 2 80.369 45.48 80.429 45.72 ;
      RECT MASK 2 80.809 45.48 80.869 45.72 ;
      RECT MASK 2 81.249 45.48 81.309 45.72 ;
      RECT MASK 2 81.689 45.48 81.749 45.72 ;
      RECT MASK 2 82.129 45.48 82.189 45.72 ;
      RECT MASK 2 83.449 45.48 83.509 45.72 ;
      RECT MASK 2 84.347 45.48 84.407 45.72 ;
      RECT MASK 2 84.787 45.48 84.847 45.72 ;
      RECT MASK 2 85.227 45.48 85.287 45.72 ;
      RECT MASK 2 85.667 45.48 85.727 45.72 ;
      RECT MASK 2 86.107 45.48 86.167 45.72 ;
      RECT MASK 2 86.547 45.48 86.607 45.72 ;
      RECT MASK 2 86.987 45.48 87.047 45.72 ;
      RECT MASK 2 87.427 45.48 87.487 45.72 ;
      RECT MASK 2 87.867 45.48 87.927 45.72 ;
      RECT MASK 2 88.307 45.48 88.367 45.72 ;
      RECT MASK 2 88.747 45.48 88.807 45.72 ;
      RECT MASK 2 89.187 45.48 89.247 45.72 ;
      RECT MASK 2 89.627 45.48 89.687 45.72 ;
      RECT MASK 2 90.067 45.48 90.127 45.72 ;
      RECT MASK 2 90.965 45.48 91.025 45.72 ;
      RECT MASK 2 91.405 45.48 91.465 45.72 ;
      RECT MASK 2 91.845 45.48 91.905 45.72 ;
      RECT MASK 2 92.285 45.48 92.345 45.72 ;
      RECT MASK 2 92.725 45.48 92.785 45.72 ;
      RECT MASK 2 93.165 45.48 93.225 45.72 ;
      RECT MASK 2 93.605 45.48 93.665 45.72 ;
      RECT MASK 2 94.045 45.48 94.105 45.72 ;
      RECT MASK 2 94.485 45.48 94.545 45.72 ;
      RECT MASK 2 94.925 45.48 94.985 45.72 ;
      RECT MASK 2 95.365 45.48 95.425 45.72 ;
      RECT MASK 2 95.805 45.48 95.865 45.72 ;
      RECT MASK 2 96.245 45.48 96.305 45.72 ;
      RECT MASK 2 96.685 45.48 96.745 45.72 ;
      RECT MASK 2 97.583 45.48 97.643 45.72 ;
      RECT MASK 2 98.023 45.48 98.083 45.72 ;
      RECT MASK 2 98.463 45.48 98.523 45.72 ;
      RECT MASK 2 98.903 45.48 98.963 45.72 ;
      RECT MASK 2 99.343 45.48 99.403 45.72 ;
      RECT MASK 2 99.783 45.48 99.843 45.72 ;
      RECT MASK 2 100.223 45.48 100.283 45.72 ;
      RECT MASK 2 100.663 45.48 100.723 45.72 ;
      RECT MASK 2 101.103 45.48 101.163 45.72 ;
      RECT MASK 2 101.543 45.48 101.603 45.72 ;
      RECT MASK 2 101.983 45.48 102.043 45.72 ;
      RECT MASK 2 102.423 45.48 102.483 45.72 ;
      RECT MASK 2 102.863 45.48 102.923 45.72 ;
      RECT MASK 2 103.303 45.48 103.363 45.72 ;
      RECT MASK 2 104.201 45.48 104.261 45.72 ;
      RECT MASK 2 104.641 45.48 104.701 45.72 ;
      RECT MASK 2 105.081 45.48 105.141 45.72 ;
      RECT MASK 2 105.521 45.48 105.581 45.72 ;
      RECT MASK 2 105.961 45.48 106.021 45.72 ;
      RECT MASK 2 106.401 45.48 106.461 45.72 ;
      RECT MASK 2 106.841 45.48 106.901 45.72 ;
      RECT MASK 2 107.281 45.48 107.341 45.72 ;
      RECT MASK 2 107.721 45.48 107.781 45.72 ;
      RECT MASK 2 108.161 45.48 108.221 45.72 ;
      RECT MASK 2 108.601 45.48 108.661 45.72 ;
      RECT MASK 2 109.041 45.48 109.101 45.72 ;
      RECT MASK 2 109.481 45.48 109.541 45.72 ;
      RECT MASK 2 109.921 45.48 109.981 45.72 ;
      RECT MASK 2 4.931 45.9 4.991 46.14 ;
      RECT MASK 2 5.371 45.9 5.431 46.14 ;
      RECT MASK 2 5.811 45.9 5.871 46.14 ;
      RECT MASK 2 6.251 45.9 6.311 46.14 ;
      RECT MASK 2 6.691 45.9 6.751 46.14 ;
      RECT MASK 2 7.131 45.9 7.191 46.14 ;
      RECT MASK 2 7.571 45.9 7.631 46.14 ;
      RECT MASK 2 8.011 45.9 8.071 46.14 ;
      RECT MASK 2 8.451 45.9 8.511 46.14 ;
      RECT MASK 2 8.891 45.9 8.951 46.14 ;
      RECT MASK 2 9.331 45.9 9.391 46.14 ;
      RECT MASK 2 9.771 45.9 9.831 46.14 ;
      RECT MASK 2 10.211 45.9 10.271 46.14 ;
      RECT MASK 2 10.651 45.9 10.711 46.14 ;
      RECT MASK 2 11.549 45.9 11.609 46.14 ;
      RECT MASK 2 11.989 45.9 12.049 46.14 ;
      RECT MASK 2 12.429 45.9 12.489 46.14 ;
      RECT MASK 2 12.869 45.9 12.929 46.14 ;
      RECT MASK 2 13.309 45.9 13.369 46.14 ;
      RECT MASK 2 13.749 45.9 13.809 46.14 ;
      RECT MASK 2 14.189 45.9 14.249 46.14 ;
      RECT MASK 2 14.629 45.9 14.689 46.14 ;
      RECT MASK 2 15.069 45.9 15.129 46.14 ;
      RECT MASK 2 15.509 45.9 15.569 46.14 ;
      RECT MASK 2 15.949 45.9 16.009 46.14 ;
      RECT MASK 2 16.389 45.9 16.449 46.14 ;
      RECT MASK 2 16.829 45.9 16.889 46.14 ;
      RECT MASK 2 17.269 45.9 17.329 46.14 ;
      RECT MASK 2 18.167 45.9 18.227 46.14 ;
      RECT MASK 2 18.607 45.9 18.667 46.14 ;
      RECT MASK 2 19.047 45.9 19.107 46.14 ;
      RECT MASK 2 19.487 45.9 19.547 46.14 ;
      RECT MASK 2 19.927 45.9 19.987 46.14 ;
      RECT MASK 2 20.367 45.9 20.427 46.14 ;
      RECT MASK 2 20.807 45.9 20.867 46.14 ;
      RECT MASK 2 21.247 45.9 21.307 46.14 ;
      RECT MASK 2 21.687 45.9 21.747 46.14 ;
      RECT MASK 2 22.127 45.9 22.187 46.14 ;
      RECT MASK 2 22.567 45.9 22.627 46.14 ;
      RECT MASK 2 23.007 45.9 23.067 46.14 ;
      RECT MASK 2 23.447 45.9 23.507 46.14 ;
      RECT MASK 2 23.887 45.9 23.947 46.14 ;
      RECT MASK 2 24.785 45.9 24.845 46.14 ;
      RECT MASK 2 25.225 45.9 25.285 46.14 ;
      RECT MASK 2 25.665 45.9 25.725 46.14 ;
      RECT MASK 2 26.105 45.9 26.165 46.14 ;
      RECT MASK 2 26.545 45.9 26.605 46.14 ;
      RECT MASK 2 26.985 45.9 27.045 46.14 ;
      RECT MASK 2 27.425 45.9 27.485 46.14 ;
      RECT MASK 2 27.865 45.9 27.925 46.14 ;
      RECT MASK 2 28.305 45.9 28.365 46.14 ;
      RECT MASK 2 28.745 45.9 28.805 46.14 ;
      RECT MASK 2 29.185 45.9 29.245 46.14 ;
      RECT MASK 2 29.625 45.9 29.685 46.14 ;
      RECT MASK 2 30.065 45.9 30.125 46.14 ;
      RECT MASK 2 30.505 45.9 30.565 46.14 ;
      RECT MASK 2 31.403 45.9 31.463 46.14 ;
      RECT MASK 2 31.843 45.9 31.903 46.14 ;
      RECT MASK 2 32.283 45.9 32.343 46.14 ;
      RECT MASK 2 32.723 45.9 32.783 46.14 ;
      RECT MASK 2 33.163 45.9 33.223 46.14 ;
      RECT MASK 2 33.603 45.9 33.663 46.14 ;
      RECT MASK 2 34.043 45.9 34.103 46.14 ;
      RECT MASK 2 34.483 45.9 34.543 46.14 ;
      RECT MASK 2 34.923 45.9 34.983 46.14 ;
      RECT MASK 2 35.363 45.9 35.423 46.14 ;
      RECT MASK 2 35.803 45.9 35.863 46.14 ;
      RECT MASK 2 36.243 45.9 36.303 46.14 ;
      RECT MASK 2 36.683 45.9 36.743 46.14 ;
      RECT MASK 2 37.123 45.9 37.183 46.14 ;
      RECT MASK 2 38.021 45.9 38.081 46.14 ;
      RECT MASK 2 38.461 45.9 38.521 46.14 ;
      RECT MASK 2 38.901 45.9 38.961 46.14 ;
      RECT MASK 2 39.341 45.9 39.401 46.14 ;
      RECT MASK 2 39.781 45.9 39.841 46.14 ;
      RECT MASK 2 40.221 45.9 40.281 46.14 ;
      RECT MASK 2 40.661 45.9 40.721 46.14 ;
      RECT MASK 2 41.101 45.9 41.161 46.14 ;
      RECT MASK 2 41.541 45.9 41.601 46.14 ;
      RECT MASK 2 42.861 45.9 42.921 46.14 ;
      RECT MASK 2 43.301 45.9 43.361 46.14 ;
      RECT MASK 2 43.741 45.9 43.801 46.14 ;
      RECT MASK 2 44.639 45.9 44.699 46.14 ;
      RECT MASK 2 45.079 45.9 45.139 46.14 ;
      RECT MASK 2 45.519 45.9 45.579 46.14 ;
      RECT MASK 2 45.959 45.9 46.019 46.14 ;
      RECT MASK 2 46.399 45.9 46.459 46.14 ;
      RECT MASK 2 46.839 45.9 46.899 46.14 ;
      RECT MASK 2 47.279 45.9 47.339 46.14 ;
      RECT MASK 2 47.719 45.9 47.779 46.14 ;
      RECT MASK 2 48.159 45.9 48.219 46.14 ;
      RECT MASK 2 48.599 45.9 48.659 46.14 ;
      RECT MASK 2 49.039 45.9 49.099 46.14 ;
      RECT MASK 2 49.479 45.9 49.539 46.14 ;
      RECT MASK 2 49.919 45.9 49.979 46.14 ;
      RECT MASK 2 50.359 45.9 50.419 46.14 ;
      RECT MASK 2 51.257 45.9 51.317 46.14 ;
      RECT MASK 2 51.697 45.9 51.757 46.14 ;
      RECT MASK 2 52.137 45.9 52.197 46.14 ;
      RECT MASK 2 52.577 45.9 52.637 46.14 ;
      RECT MASK 2 53.017 45.9 53.077 46.14 ;
      RECT MASK 2 53.457 45.9 53.517 46.14 ;
      RECT MASK 2 53.897 45.9 53.957 46.14 ;
      RECT MASK 2 54.337 45.9 54.397 46.14 ;
      RECT MASK 2 54.777 45.9 54.837 46.14 ;
      RECT MASK 2 55.217 45.9 55.277 46.14 ;
      RECT MASK 2 55.657 45.9 55.717 46.14 ;
      RECT MASK 2 56.097 45.9 56.157 46.14 ;
      RECT MASK 2 56.537 45.9 56.597 46.14 ;
      RECT MASK 2 56.977 45.9 57.037 46.14 ;
      RECT MASK 2 57.875 45.9 57.935 46.14 ;
      RECT MASK 2 58.315 45.9 58.375 46.14 ;
      RECT MASK 2 58.755 45.9 58.815 46.14 ;
      RECT MASK 2 59.195 45.9 59.255 46.14 ;
      RECT MASK 2 59.635 45.9 59.695 46.14 ;
      RECT MASK 2 60.075 45.9 60.135 46.14 ;
      RECT MASK 2 60.515 45.9 60.575 46.14 ;
      RECT MASK 2 60.955 45.9 61.015 46.14 ;
      RECT MASK 2 61.395 45.9 61.455 46.14 ;
      RECT MASK 2 61.835 45.9 61.895 46.14 ;
      RECT MASK 2 62.275 45.9 62.335 46.14 ;
      RECT MASK 2 62.715 45.9 62.775 46.14 ;
      RECT MASK 2 63.155 45.9 63.215 46.14 ;
      RECT MASK 2 63.595 45.9 63.655 46.14 ;
      RECT MASK 2 64.493 45.9 64.553 46.14 ;
      RECT MASK 2 64.933 45.9 64.993 46.14 ;
      RECT MASK 2 65.373 45.9 65.433 46.14 ;
      RECT MASK 2 65.813 45.9 65.873 46.14 ;
      RECT MASK 2 66.253 45.9 66.313 46.14 ;
      RECT MASK 2 66.693 45.9 66.753 46.14 ;
      RECT MASK 2 67.133 45.9 67.193 46.14 ;
      RECT MASK 2 67.573 45.9 67.633 46.14 ;
      RECT MASK 2 68.013 45.9 68.073 46.14 ;
      RECT MASK 2 68.453 45.9 68.513 46.14 ;
      RECT MASK 2 68.893 45.9 68.953 46.14 ;
      RECT MASK 2 69.333 45.9 69.393 46.14 ;
      RECT MASK 2 69.773 45.9 69.833 46.14 ;
      RECT MASK 2 70.213 45.9 70.273 46.14 ;
      RECT MASK 2 71.111 45.9 71.171 46.14 ;
      RECT MASK 2 71.551 45.9 71.611 46.14 ;
      RECT MASK 2 71.991 45.9 72.051 46.14 ;
      RECT MASK 2 72.431 45.9 72.491 46.14 ;
      RECT MASK 2 72.871 45.9 72.931 46.14 ;
      RECT MASK 2 73.311 45.9 73.371 46.14 ;
      RECT MASK 2 73.751 45.9 73.811 46.14 ;
      RECT MASK 2 74.191 45.9 74.251 46.14 ;
      RECT MASK 2 74.631 45.9 74.691 46.14 ;
      RECT MASK 2 75.071 45.9 75.131 46.14 ;
      RECT MASK 2 75.511 45.9 75.571 46.14 ;
      RECT MASK 2 75.951 45.9 76.011 46.14 ;
      RECT MASK 2 76.391 45.9 76.451 46.14 ;
      RECT MASK 2 76.831 45.9 76.891 46.14 ;
      RECT MASK 2 77.729 45.9 77.789 46.14 ;
      RECT MASK 2 78.169 45.9 78.229 46.14 ;
      RECT MASK 2 78.609 45.9 78.669 46.14 ;
      RECT MASK 2 79.049 45.9 79.109 46.14 ;
      RECT MASK 2 79.489 45.9 79.549 46.14 ;
      RECT MASK 2 79.929 45.9 79.989 46.14 ;
      RECT MASK 2 80.369 45.9 80.429 46.14 ;
      RECT MASK 2 80.809 45.9 80.869 46.14 ;
      RECT MASK 2 81.249 45.9 81.309 46.14 ;
      RECT MASK 2 81.689 45.9 81.749 46.14 ;
      RECT MASK 2 82.129 45.9 82.189 46.14 ;
      RECT MASK 2 83.449 45.9 83.509 46.14 ;
      RECT MASK 2 84.347 45.9 84.407 46.14 ;
      RECT MASK 2 84.787 45.9 84.847 46.14 ;
      RECT MASK 2 85.227 45.9 85.287 46.14 ;
      RECT MASK 2 85.667 45.9 85.727 46.14 ;
      RECT MASK 2 86.107 45.9 86.167 46.14 ;
      RECT MASK 2 86.547 45.9 86.607 46.14 ;
      RECT MASK 2 86.987 45.9 87.047 46.14 ;
      RECT MASK 2 87.427 45.9 87.487 46.14 ;
      RECT MASK 2 87.867 45.9 87.927 46.14 ;
      RECT MASK 2 88.307 45.9 88.367 46.14 ;
      RECT MASK 2 88.747 45.9 88.807 46.14 ;
      RECT MASK 2 89.187 45.9 89.247 46.14 ;
      RECT MASK 2 89.627 45.9 89.687 46.14 ;
      RECT MASK 2 90.067 45.9 90.127 46.14 ;
      RECT MASK 2 90.965 45.9 91.025 46.14 ;
      RECT MASK 2 91.405 45.9 91.465 46.14 ;
      RECT MASK 2 91.845 45.9 91.905 46.14 ;
      RECT MASK 2 92.285 45.9 92.345 46.14 ;
      RECT MASK 2 92.725 45.9 92.785 46.14 ;
      RECT MASK 2 93.165 45.9 93.225 46.14 ;
      RECT MASK 2 93.605 45.9 93.665 46.14 ;
      RECT MASK 2 94.045 45.9 94.105 46.14 ;
      RECT MASK 2 94.485 45.9 94.545 46.14 ;
      RECT MASK 2 94.925 45.9 94.985 46.14 ;
      RECT MASK 2 95.365 45.9 95.425 46.14 ;
      RECT MASK 2 95.805 45.9 95.865 46.14 ;
      RECT MASK 2 96.245 45.9 96.305 46.14 ;
      RECT MASK 2 96.685 45.9 96.745 46.14 ;
      RECT MASK 2 97.583 45.9 97.643 46.14 ;
      RECT MASK 2 98.023 45.9 98.083 46.14 ;
      RECT MASK 2 98.463 45.9 98.523 46.14 ;
      RECT MASK 2 98.903 45.9 98.963 46.14 ;
      RECT MASK 2 99.343 45.9 99.403 46.14 ;
      RECT MASK 2 99.783 45.9 99.843 46.14 ;
      RECT MASK 2 100.223 45.9 100.283 46.14 ;
      RECT MASK 2 100.663 45.9 100.723 46.14 ;
      RECT MASK 2 101.103 45.9 101.163 46.14 ;
      RECT MASK 2 101.543 45.9 101.603 46.14 ;
      RECT MASK 2 101.983 45.9 102.043 46.14 ;
      RECT MASK 2 102.423 45.9 102.483 46.14 ;
      RECT MASK 2 102.863 45.9 102.923 46.14 ;
      RECT MASK 2 103.303 45.9 103.363 46.14 ;
      RECT MASK 2 104.201 45.9 104.261 46.14 ;
      RECT MASK 2 104.641 45.9 104.701 46.14 ;
      RECT MASK 2 105.081 45.9 105.141 46.14 ;
      RECT MASK 2 105.521 45.9 105.581 46.14 ;
      RECT MASK 2 105.961 45.9 106.021 46.14 ;
      RECT MASK 2 106.401 45.9 106.461 46.14 ;
      RECT MASK 2 106.841 45.9 106.901 46.14 ;
      RECT MASK 2 107.281 45.9 107.341 46.14 ;
      RECT MASK 2 107.721 45.9 107.781 46.14 ;
      RECT MASK 2 108.161 45.9 108.221 46.14 ;
      RECT MASK 2 108.601 45.9 108.661 46.14 ;
      RECT MASK 2 109.041 45.9 109.101 46.14 ;
      RECT MASK 2 109.481 45.9 109.541 46.14 ;
      RECT MASK 2 109.921 45.9 109.981 46.14 ;
      RECT MASK 2 4.901 46.339 5.021 57.551 ;
      RECT MASK 2 5.341 46.339 5.461 57.551 ;
      RECT MASK 2 5.781 46.339 5.901 57.551 ;
      RECT MASK 2 6.221 46.339 6.341 57.551 ;
      RECT MASK 2 6.661 46.339 6.781 57.551 ;
      RECT MASK 2 7.101 46.339 7.221 57.551 ;
      RECT MASK 2 7.541 46.339 7.661 57.551 ;
      RECT MASK 2 7.981 46.339 8.101 57.551 ;
      RECT MASK 2 8.421 46.339 8.541 57.551 ;
      RECT MASK 2 8.861 46.339 8.981 57.551 ;
      RECT MASK 2 9.301 46.339 9.421 57.551 ;
      RECT MASK 2 9.741 46.339 9.861 57.551 ;
      RECT MASK 2 10.181 46.339 10.301 57.551 ;
      RECT MASK 2 10.621 46.339 10.741 57.551 ;
      RECT MASK 2 11.519 46.339 11.639 51.431 ;
      RECT MASK 2 11.959 46.339 12.079 51.431 ;
      RECT MASK 2 12.399 46.339 12.519 51.431 ;
      RECT MASK 2 12.839 46.339 12.959 51.431 ;
      RECT MASK 2 13.279 46.339 13.399 51.431 ;
      RECT MASK 2 13.719 46.339 13.839 51.431 ;
      RECT MASK 2 14.159 46.339 14.279 51.431 ;
      RECT MASK 2 14.599 46.339 14.719 51.431 ;
      RECT MASK 2 15.039 46.339 15.159 51.431 ;
      RECT MASK 2 15.479 46.339 15.599 51.431 ;
      RECT MASK 2 15.919 46.339 16.039 51.431 ;
      RECT MASK 2 16.359 46.339 16.479 51.431 ;
      RECT MASK 2 16.799 46.339 16.919 51.431 ;
      RECT MASK 2 17.239 46.339 17.359 51.431 ;
      RECT MASK 2 18.137 46.339 18.257 51.431 ;
      RECT MASK 2 18.577 46.339 18.697 51.431 ;
      RECT MASK 2 19.017 46.339 19.137 51.431 ;
      RECT MASK 2 19.457 46.339 19.577 51.431 ;
      RECT MASK 2 19.897 46.339 20.017 51.431 ;
      RECT MASK 2 20.337 46.339 20.457 51.431 ;
      RECT MASK 2 20.777 46.339 20.897 51.431 ;
      RECT MASK 2 21.217 46.339 21.337 51.431 ;
      RECT MASK 2 21.657 46.339 21.777 51.431 ;
      RECT MASK 2 22.097 46.339 22.217 51.431 ;
      RECT MASK 2 22.537 46.339 22.657 51.431 ;
      RECT MASK 2 22.977 46.339 23.097 51.431 ;
      RECT MASK 2 23.417 46.339 23.537 51.431 ;
      RECT MASK 2 23.857 46.339 23.977 51.431 ;
      RECT MASK 2 24.755 46.339 24.875 51.431 ;
      RECT MASK 2 25.195 46.339 25.315 51.431 ;
      RECT MASK 2 25.635 46.339 25.755 51.431 ;
      RECT MASK 2 26.075 46.339 26.195 51.431 ;
      RECT MASK 2 26.515 46.339 26.635 51.431 ;
      RECT MASK 2 26.955 46.339 27.075 51.431 ;
      RECT MASK 2 27.395 46.339 27.515 51.431 ;
      RECT MASK 2 27.835 46.339 27.955 51.431 ;
      RECT MASK 2 28.275 46.339 28.395 51.431 ;
      RECT MASK 2 28.715 46.339 28.835 51.431 ;
      RECT MASK 2 29.155 46.339 29.275 51.431 ;
      RECT MASK 2 29.595 46.339 29.715 51.431 ;
      RECT MASK 2 30.035 46.339 30.155 51.431 ;
      RECT MASK 2 30.475 46.339 30.595 51.431 ;
      RECT MASK 2 31.373 46.339 31.493 51.431 ;
      RECT MASK 2 31.813 46.339 31.933 51.431 ;
      RECT MASK 2 32.253 46.339 32.373 51.431 ;
      RECT MASK 2 32.693 46.339 32.813 51.431 ;
      RECT MASK 2 33.133 46.339 33.253 51.431 ;
      RECT MASK 2 33.573 46.339 33.693 51.431 ;
      RECT MASK 2 34.013 46.339 34.133 51.431 ;
      RECT MASK 2 34.453 46.339 34.573 51.431 ;
      RECT MASK 2 34.893 46.339 35.013 51.431 ;
      RECT MASK 2 35.333 46.339 35.453 51.431 ;
      RECT MASK 2 35.773 46.339 35.893 51.431 ;
      RECT MASK 2 36.213 46.339 36.333 51.431 ;
      RECT MASK 2 36.653 46.339 36.773 51.431 ;
      RECT MASK 2 37.093 46.339 37.213 51.431 ;
      RECT MASK 2 37.991 46.339 38.111 51.431 ;
      RECT MASK 2 38.431 46.339 38.551 51.431 ;
      RECT MASK 2 38.871 46.339 38.991 51.431 ;
      RECT MASK 2 39.311 46.339 39.431 51.431 ;
      RECT MASK 2 39.751 46.339 39.871 51.431 ;
      RECT MASK 2 40.191 46.339 40.311 51.431 ;
      RECT MASK 2 40.631 46.339 40.751 51.431 ;
      RECT MASK 2 41.071 46.339 41.191 51.431 ;
      RECT MASK 2 41.511 46.339 41.631 51.431 ;
      RECT MASK 2 41.951 46.339 42.071 51.431 ;
      RECT MASK 2 42.391 46.339 42.511 51.431 ;
      RECT MASK 2 42.831 46.339 42.951 51.431 ;
      RECT MASK 2 43.271 46.339 43.391 51.431 ;
      RECT MASK 2 43.711 46.339 43.831 51.431 ;
      RECT MASK 2 44.609 46.339 44.729 51.431 ;
      RECT MASK 2 45.049 46.339 45.169 51.431 ;
      RECT MASK 2 45.489 46.339 45.609 51.431 ;
      RECT MASK 2 45.929 46.339 46.049 51.431 ;
      RECT MASK 2 46.369 46.339 46.489 51.431 ;
      RECT MASK 2 46.809 46.339 46.929 51.431 ;
      RECT MASK 2 47.249 46.339 47.369 51.431 ;
      RECT MASK 2 47.689 46.339 47.809 51.431 ;
      RECT MASK 2 48.129 46.339 48.249 51.431 ;
      RECT MASK 2 48.569 46.339 48.689 51.431 ;
      RECT MASK 2 49.009 46.339 49.129 51.431 ;
      RECT MASK 2 49.449 46.339 49.569 51.431 ;
      RECT MASK 2 49.889 46.339 50.009 51.431 ;
      RECT MASK 2 50.329 46.339 50.449 51.431 ;
      RECT MASK 2 51.227 46.339 51.347 51.431 ;
      RECT MASK 2 51.667 46.339 51.787 51.431 ;
      RECT MASK 2 52.107 46.339 52.227 51.431 ;
      RECT MASK 2 52.547 46.339 52.667 51.431 ;
      RECT MASK 2 52.987 46.339 53.107 51.431 ;
      RECT MASK 2 53.427 46.339 53.547 51.431 ;
      RECT MASK 2 53.867 46.339 53.987 51.431 ;
      RECT MASK 2 54.307 46.339 54.427 51.431 ;
      RECT MASK 2 54.747 46.339 54.867 51.431 ;
      RECT MASK 2 55.187 46.339 55.307 51.431 ;
      RECT MASK 2 55.627 46.339 55.747 51.431 ;
      RECT MASK 2 56.067 46.339 56.187 51.431 ;
      RECT MASK 2 56.507 46.339 56.627 51.431 ;
      RECT MASK 2 56.947 46.339 57.067 51.431 ;
      RECT MASK 2 57.845 46.339 57.965 51.431 ;
      RECT MASK 2 58.285 46.339 58.405 51.431 ;
      RECT MASK 2 58.725 46.339 58.845 51.431 ;
      RECT MASK 2 59.165 46.339 59.285 51.431 ;
      RECT MASK 2 59.605 46.339 59.725 51.431 ;
      RECT MASK 2 60.045 46.339 60.165 51.431 ;
      RECT MASK 2 60.485 46.339 60.605 51.431 ;
      RECT MASK 2 60.925 46.339 61.045 51.431 ;
      RECT MASK 2 61.365 46.339 61.485 51.431 ;
      RECT MASK 2 61.805 46.339 61.925 51.431 ;
      RECT MASK 2 62.245 46.339 62.365 51.431 ;
      RECT MASK 2 62.685 46.339 62.805 51.431 ;
      RECT MASK 2 63.125 46.339 63.245 51.431 ;
      RECT MASK 2 63.565 46.339 63.685 51.431 ;
      RECT MASK 2 64.463 46.339 64.583 51.431 ;
      RECT MASK 2 64.903 46.339 65.023 51.431 ;
      RECT MASK 2 65.343 46.339 65.463 51.431 ;
      RECT MASK 2 65.783 46.339 65.903 51.431 ;
      RECT MASK 2 66.223 46.339 66.343 51.431 ;
      RECT MASK 2 66.663 46.339 66.783 51.431 ;
      RECT MASK 2 67.103 46.339 67.223 51.431 ;
      RECT MASK 2 67.543 46.339 67.663 51.431 ;
      RECT MASK 2 67.983 46.339 68.103 51.431 ;
      RECT MASK 2 68.423 46.339 68.543 51.431 ;
      RECT MASK 2 68.863 46.339 68.983 51.431 ;
      RECT MASK 2 69.303 46.339 69.423 51.431 ;
      RECT MASK 2 69.743 46.339 69.863 51.431 ;
      RECT MASK 2 70.183 46.339 70.303 51.431 ;
      RECT MASK 2 71.081 46.339 71.201 51.431 ;
      RECT MASK 2 71.521 46.339 71.641 51.431 ;
      RECT MASK 2 71.961 46.339 72.081 51.431 ;
      RECT MASK 2 72.401 46.339 72.521 51.431 ;
      RECT MASK 2 72.841 46.339 72.961 51.431 ;
      RECT MASK 2 73.281 46.339 73.401 51.431 ;
      RECT MASK 2 73.721 46.339 73.841 51.431 ;
      RECT MASK 2 74.161 46.339 74.281 51.431 ;
      RECT MASK 2 74.601 46.339 74.721 51.431 ;
      RECT MASK 2 75.041 46.339 75.161 51.431 ;
      RECT MASK 2 75.481 46.339 75.601 51.431 ;
      RECT MASK 2 75.921 46.339 76.041 51.431 ;
      RECT MASK 2 76.361 46.339 76.481 51.431 ;
      RECT MASK 2 76.801 46.339 76.921 51.431 ;
      RECT MASK 2 77.699 46.339 77.819 51.431 ;
      RECT MASK 2 78.139 46.339 78.259 51.431 ;
      RECT MASK 2 78.579 46.339 78.699 51.431 ;
      RECT MASK 2 79.019 46.339 79.139 51.431 ;
      RECT MASK 2 79.459 46.339 79.579 51.431 ;
      RECT MASK 2 79.899 46.339 80.019 51.431 ;
      RECT MASK 2 80.339 46.339 80.459 51.431 ;
      RECT MASK 2 80.779 46.339 80.899 51.431 ;
      RECT MASK 2 81.219 46.339 81.339 51.431 ;
      RECT MASK 2 81.659 46.339 81.779 51.431 ;
      RECT MASK 2 82.099 46.339 82.219 51.431 ;
      RECT MASK 2 82.539 46.339 82.659 51.431 ;
      RECT MASK 2 82.979 46.339 83.099 51.431 ;
      RECT MASK 2 83.419 46.339 83.539 51.431 ;
      RECT MASK 2 84.317 46.339 84.437 51.431 ;
      RECT MASK 2 84.757 46.339 84.877 51.431 ;
      RECT MASK 2 85.197 46.339 85.317 51.431 ;
      RECT MASK 2 85.637 46.339 85.757 51.431 ;
      RECT MASK 2 86.077 46.339 86.197 51.431 ;
      RECT MASK 2 86.517 46.339 86.637 51.431 ;
      RECT MASK 2 86.957 46.339 87.077 51.431 ;
      RECT MASK 2 87.397 46.339 87.517 51.431 ;
      RECT MASK 2 87.837 46.339 87.957 51.431 ;
      RECT MASK 2 88.277 46.339 88.397 51.431 ;
      RECT MASK 2 88.717 46.339 88.837 51.431 ;
      RECT MASK 2 89.157 46.339 89.277 51.431 ;
      RECT MASK 2 89.597 46.339 89.717 51.431 ;
      RECT MASK 2 90.037 46.339 90.157 51.431 ;
      RECT MASK 2 90.935 46.339 91.055 51.431 ;
      RECT MASK 2 91.375 46.339 91.495 51.431 ;
      RECT MASK 2 91.815 46.339 91.935 51.431 ;
      RECT MASK 2 92.255 46.339 92.375 51.431 ;
      RECT MASK 2 92.695 46.339 92.815 51.431 ;
      RECT MASK 2 93.135 46.339 93.255 51.431 ;
      RECT MASK 2 93.575 46.339 93.695 51.431 ;
      RECT MASK 2 94.015 46.339 94.135 51.431 ;
      RECT MASK 2 94.455 46.339 94.575 51.431 ;
      RECT MASK 2 94.895 46.339 95.015 51.431 ;
      RECT MASK 2 95.335 46.339 95.455 51.431 ;
      RECT MASK 2 95.775 46.339 95.895 51.431 ;
      RECT MASK 2 96.215 46.339 96.335 51.431 ;
      RECT MASK 2 96.655 46.339 96.775 51.431 ;
      RECT MASK 2 97.553 46.339 97.673 51.431 ;
      RECT MASK 2 97.993 46.339 98.113 51.431 ;
      RECT MASK 2 98.433 46.339 98.553 51.431 ;
      RECT MASK 2 98.873 46.339 98.993 51.431 ;
      RECT MASK 2 99.313 46.339 99.433 51.431 ;
      RECT MASK 2 99.753 46.339 99.873 51.431 ;
      RECT MASK 2 100.193 46.339 100.313 51.431 ;
      RECT MASK 2 100.633 46.339 100.753 51.431 ;
      RECT MASK 2 101.073 46.339 101.193 51.431 ;
      RECT MASK 2 101.513 46.339 101.633 51.431 ;
      RECT MASK 2 101.953 46.339 102.073 51.431 ;
      RECT MASK 2 102.393 46.339 102.513 51.431 ;
      RECT MASK 2 102.833 46.339 102.953 51.431 ;
      RECT MASK 2 103.273 46.339 103.393 51.431 ;
      RECT MASK 2 104.171 46.339 104.291 51.431 ;
      RECT MASK 2 104.611 46.339 104.731 51.431 ;
      RECT MASK 2 105.051 46.339 105.171 51.431 ;
      RECT MASK 2 105.491 46.339 105.611 51.431 ;
      RECT MASK 2 105.931 46.339 106.051 51.431 ;
      RECT MASK 2 106.371 46.339 106.491 51.431 ;
      RECT MASK 2 106.811 46.339 106.931 51.431 ;
      RECT MASK 2 107.251 46.339 107.371 51.431 ;
      RECT MASK 2 107.691 46.339 107.811 51.431 ;
      RECT MASK 2 108.131 46.339 108.251 51.431 ;
      RECT MASK 2 108.571 46.339 108.691 51.431 ;
      RECT MASK 2 109.011 46.339 109.131 51.431 ;
      RECT MASK 2 109.451 46.339 109.571 51.431 ;
      RECT MASK 2 109.891 46.339 110.011 51.431 ;
      RECT MASK 2 112.5865 46.969 112.7065 48.119 ;
      RECT MASK 2 113.0265 46.969 113.1465 48.119 ;
      RECT MASK 2 113.4665 46.969 113.5865 48.119 ;
      RECT MASK 2 113.9065 46.969 114.0265 48.119 ;
      RECT MASK 2 114.3465 46.969 114.4665 48.119 ;
      RECT MASK 2 114.7865 46.969 114.9065 48.119 ;
      RECT MASK 2 115.2265 46.969 115.3465 48.119 ;
      RECT MASK 2 115.6665 46.969 115.7865 48.119 ;
      RECT MASK 2 116.1065 46.969 116.2265 48.119 ;
      RECT MASK 2 116.5465 46.969 116.6665 48.119 ;
      RECT MASK 2 117.4265 46.969 117.5465 48.059 ;
      RECT MASK 2 117.8665 46.969 117.9865 48.059 ;
      RECT MASK 2 118.3065 46.969 118.4265 48.059 ;
      RECT MASK 2 118.7465 46.969 118.8665 48.059 ;
      RECT MASK 2 119.1865 46.969 119.3065 48.059 ;
      RECT MASK 2 119.6265 46.969 119.7465 48.059 ;
      RECT MASK 2 120.0665 46.969 120.1865 48.059 ;
      RECT MASK 2 120.5065 46.969 120.6265 48.059 ;
      RECT MASK 2 120.9465 46.969 121.0665 48.059 ;
      RECT MASK 2 121.3865 46.969 121.5065 48.059 ;
      RECT MASK 2 121.8265 46.969 121.9465 48.059 ;
      RECT MASK 2 122.2665 46.969 122.3865 48.059 ;
      RECT MASK 2 122.7065 46.969 122.8265 48.059 ;
      RECT MASK 2 123.1465 46.969 123.2665 48.059 ;
      RECT MASK 2 123.5865 46.969 123.7065 48.059 ;
      RECT MASK 2 112.5865 48.379 112.7065 49.409 ;
      RECT MASK 2 113.0265 48.379 113.1465 49.409 ;
      RECT MASK 2 113.4665 48.379 113.5865 49.409 ;
      RECT MASK 2 113.9065 48.379 114.0265 49.409 ;
      RECT MASK 2 114.3465 48.379 114.4665 49.409 ;
      RECT MASK 2 114.7865 48.379 114.9065 49.409 ;
      RECT MASK 2 115.2265 48.379 115.3465 49.409 ;
      RECT MASK 2 115.6665 48.379 115.7865 49.409 ;
      RECT MASK 2 116.1065 48.379 116.2265 49.409 ;
      RECT MASK 2 116.5465 48.379 116.6665 49.409 ;
      RECT MASK 2 117.4265 49.269 117.5465 50.759 ;
      RECT MASK 2 117.8665 49.269 117.9865 50.759 ;
      RECT MASK 2 118.3065 49.269 118.4265 50.759 ;
      RECT MASK 2 118.7465 49.269 118.8665 50.759 ;
      RECT MASK 2 119.1865 49.269 119.3065 50.759 ;
      RECT MASK 2 119.6265 49.269 119.7465 50.759 ;
      RECT MASK 2 120.0665 49.269 120.1865 50.759 ;
      RECT MASK 2 120.5065 49.269 120.6265 50.759 ;
      RECT MASK 2 120.9465 49.269 121.0665 50.759 ;
      RECT MASK 2 121.3865 49.269 121.5065 50.759 ;
      RECT MASK 2 121.8265 49.269 121.9465 50.759 ;
      RECT MASK 2 122.2665 49.269 122.3865 50.759 ;
      RECT MASK 2 122.7065 49.269 122.8265 50.759 ;
      RECT MASK 2 123.1465 49.269 123.2665 50.759 ;
      RECT MASK 2 112.5865 49.669 112.7065 50.759 ;
      RECT MASK 2 113.0265 49.669 113.1465 50.759 ;
      RECT MASK 2 113.4665 49.669 113.5865 50.759 ;
      RECT MASK 2 113.9065 49.669 114.0265 50.759 ;
      RECT MASK 2 114.3465 49.669 114.4665 50.759 ;
      RECT MASK 2 114.7865 49.669 114.9065 50.759 ;
      RECT MASK 2 115.2265 49.669 115.3465 50.759 ;
      RECT MASK 2 115.6665 49.669 115.7865 50.759 ;
      RECT MASK 2 116.1065 49.669 116.2265 50.759 ;
      RECT MASK 2 116.5465 49.669 116.6665 50.759 ;
      RECT MASK 2 11.519 52.459 11.639 57.551 ;
      RECT MASK 2 11.959 52.459 12.079 57.551 ;
      RECT MASK 2 12.399 52.459 12.519 57.551 ;
      RECT MASK 2 12.839 52.459 12.959 57.551 ;
      RECT MASK 2 13.279 52.459 13.399 57.551 ;
      RECT MASK 2 13.719 52.459 13.839 57.551 ;
      RECT MASK 2 14.159 52.459 14.279 57.551 ;
      RECT MASK 2 14.599 52.459 14.719 57.551 ;
      RECT MASK 2 15.039 52.459 15.159 57.551 ;
      RECT MASK 2 15.479 52.459 15.599 57.551 ;
      RECT MASK 2 15.919 52.459 16.039 57.551 ;
      RECT MASK 2 16.359 52.459 16.479 57.551 ;
      RECT MASK 2 16.799 52.459 16.919 57.551 ;
      RECT MASK 2 17.239 52.459 17.359 57.551 ;
      RECT MASK 2 18.137 52.459 18.257 57.551 ;
      RECT MASK 2 18.577 52.459 18.697 57.551 ;
      RECT MASK 2 19.017 52.459 19.137 57.551 ;
      RECT MASK 2 19.457 52.459 19.577 57.551 ;
      RECT MASK 2 19.897 52.459 20.017 57.551 ;
      RECT MASK 2 20.337 52.459 20.457 57.551 ;
      RECT MASK 2 20.777 52.459 20.897 57.551 ;
      RECT MASK 2 21.217 52.459 21.337 57.551 ;
      RECT MASK 2 21.657 52.459 21.777 57.551 ;
      RECT MASK 2 22.097 52.459 22.217 57.551 ;
      RECT MASK 2 22.537 52.459 22.657 57.551 ;
      RECT MASK 2 22.977 52.459 23.097 57.551 ;
      RECT MASK 2 23.417 52.459 23.537 57.551 ;
      RECT MASK 2 23.857 52.459 23.977 57.551 ;
      RECT MASK 2 24.755 52.459 24.875 57.551 ;
      RECT MASK 2 25.195 52.459 25.315 57.551 ;
      RECT MASK 2 25.635 52.459 25.755 57.551 ;
      RECT MASK 2 26.075 52.459 26.195 57.551 ;
      RECT MASK 2 26.515 52.459 26.635 57.551 ;
      RECT MASK 2 26.955 52.459 27.075 57.551 ;
      RECT MASK 2 27.395 52.459 27.515 57.551 ;
      RECT MASK 2 27.835 52.459 27.955 57.551 ;
      RECT MASK 2 28.275 52.459 28.395 57.551 ;
      RECT MASK 2 28.715 52.459 28.835 57.551 ;
      RECT MASK 2 29.155 52.459 29.275 57.551 ;
      RECT MASK 2 29.595 52.459 29.715 57.551 ;
      RECT MASK 2 30.035 52.459 30.155 57.551 ;
      RECT MASK 2 30.475 52.459 30.595 57.551 ;
      RECT MASK 2 31.373 52.459 31.493 57.551 ;
      RECT MASK 2 31.813 52.459 31.933 57.551 ;
      RECT MASK 2 32.253 52.459 32.373 57.551 ;
      RECT MASK 2 32.693 52.459 32.813 57.551 ;
      RECT MASK 2 33.133 52.459 33.253 57.551 ;
      RECT MASK 2 33.573 52.459 33.693 57.551 ;
      RECT MASK 2 34.013 52.459 34.133 57.551 ;
      RECT MASK 2 34.453 52.459 34.573 57.551 ;
      RECT MASK 2 34.893 52.459 35.013 57.551 ;
      RECT MASK 2 35.333 52.459 35.453 57.551 ;
      RECT MASK 2 35.773 52.459 35.893 57.551 ;
      RECT MASK 2 36.213 52.459 36.333 57.551 ;
      RECT MASK 2 36.653 52.459 36.773 57.551 ;
      RECT MASK 2 37.093 52.459 37.213 57.551 ;
      RECT MASK 2 37.991 52.459 38.111 57.551 ;
      RECT MASK 2 38.431 52.459 38.551 57.551 ;
      RECT MASK 2 38.871 52.459 38.991 57.551 ;
      RECT MASK 2 39.311 52.459 39.431 57.551 ;
      RECT MASK 2 39.751 52.459 39.871 57.551 ;
      RECT MASK 2 40.191 52.459 40.311 57.551 ;
      RECT MASK 2 40.631 52.459 40.751 57.551 ;
      RECT MASK 2 41.071 52.459 41.191 57.551 ;
      RECT MASK 2 41.511 52.459 41.631 57.551 ;
      RECT MASK 2 41.951 52.459 42.071 57.551 ;
      RECT MASK 2 42.391 52.459 42.511 57.551 ;
      RECT MASK 2 42.831 52.459 42.951 57.551 ;
      RECT MASK 2 43.271 52.459 43.391 57.551 ;
      RECT MASK 2 43.711 52.459 43.831 57.551 ;
      RECT MASK 2 44.609 52.459 44.729 57.551 ;
      RECT MASK 2 45.049 52.459 45.169 57.551 ;
      RECT MASK 2 45.489 52.459 45.609 57.551 ;
      RECT MASK 2 45.929 52.459 46.049 57.551 ;
      RECT MASK 2 46.369 52.459 46.489 57.551 ;
      RECT MASK 2 46.809 52.459 46.929 57.551 ;
      RECT MASK 2 47.249 52.459 47.369 57.551 ;
      RECT MASK 2 47.689 52.459 47.809 57.551 ;
      RECT MASK 2 48.129 52.459 48.249 57.551 ;
      RECT MASK 2 48.569 52.459 48.689 57.551 ;
      RECT MASK 2 49.009 52.459 49.129 57.551 ;
      RECT MASK 2 49.449 52.459 49.569 57.551 ;
      RECT MASK 2 49.889 52.459 50.009 57.551 ;
      RECT MASK 2 50.329 52.459 50.449 57.551 ;
      RECT MASK 2 51.227 52.459 51.347 57.551 ;
      RECT MASK 2 51.667 52.459 51.787 57.551 ;
      RECT MASK 2 52.107 52.459 52.227 57.551 ;
      RECT MASK 2 52.547 52.459 52.667 57.551 ;
      RECT MASK 2 52.987 52.459 53.107 57.551 ;
      RECT MASK 2 53.427 52.459 53.547 57.551 ;
      RECT MASK 2 53.867 52.459 53.987 57.551 ;
      RECT MASK 2 54.307 52.459 54.427 57.551 ;
      RECT MASK 2 54.747 52.459 54.867 57.551 ;
      RECT MASK 2 55.187 52.459 55.307 57.551 ;
      RECT MASK 2 55.627 52.459 55.747 57.551 ;
      RECT MASK 2 56.067 52.459 56.187 57.551 ;
      RECT MASK 2 56.507 52.459 56.627 57.551 ;
      RECT MASK 2 56.947 52.459 57.067 57.551 ;
      RECT MASK 2 57.845 52.459 57.965 57.551 ;
      RECT MASK 2 58.285 52.459 58.405 57.551 ;
      RECT MASK 2 58.725 52.459 58.845 57.551 ;
      RECT MASK 2 59.165 52.459 59.285 57.551 ;
      RECT MASK 2 59.605 52.459 59.725 57.551 ;
      RECT MASK 2 60.045 52.459 60.165 57.551 ;
      RECT MASK 2 60.485 52.459 60.605 57.551 ;
      RECT MASK 2 60.925 52.459 61.045 57.551 ;
      RECT MASK 2 61.365 52.459 61.485 57.551 ;
      RECT MASK 2 61.805 52.459 61.925 57.551 ;
      RECT MASK 2 62.245 52.459 62.365 57.551 ;
      RECT MASK 2 62.685 52.459 62.805 57.551 ;
      RECT MASK 2 63.125 52.459 63.245 57.551 ;
      RECT MASK 2 63.565 52.459 63.685 57.551 ;
      RECT MASK 2 64.463 52.459 64.583 57.551 ;
      RECT MASK 2 64.903 52.459 65.023 57.551 ;
      RECT MASK 2 65.343 52.459 65.463 57.551 ;
      RECT MASK 2 65.783 52.459 65.903 57.551 ;
      RECT MASK 2 66.223 52.459 66.343 57.551 ;
      RECT MASK 2 66.663 52.459 66.783 57.551 ;
      RECT MASK 2 67.103 52.459 67.223 57.551 ;
      RECT MASK 2 67.543 52.459 67.663 57.551 ;
      RECT MASK 2 67.983 52.459 68.103 57.551 ;
      RECT MASK 2 68.423 52.459 68.543 57.551 ;
      RECT MASK 2 68.863 52.459 68.983 57.551 ;
      RECT MASK 2 69.303 52.459 69.423 57.551 ;
      RECT MASK 2 69.743 52.459 69.863 57.551 ;
      RECT MASK 2 70.183 52.459 70.303 57.551 ;
      RECT MASK 2 71.081 52.459 71.201 57.551 ;
      RECT MASK 2 71.521 52.459 71.641 57.551 ;
      RECT MASK 2 71.961 52.459 72.081 57.551 ;
      RECT MASK 2 72.401 52.459 72.521 57.551 ;
      RECT MASK 2 72.841 52.459 72.961 57.551 ;
      RECT MASK 2 73.281 52.459 73.401 57.551 ;
      RECT MASK 2 73.721 52.459 73.841 57.551 ;
      RECT MASK 2 74.161 52.459 74.281 57.551 ;
      RECT MASK 2 74.601 52.459 74.721 57.551 ;
      RECT MASK 2 75.041 52.459 75.161 57.551 ;
      RECT MASK 2 75.481 52.459 75.601 57.551 ;
      RECT MASK 2 75.921 52.459 76.041 57.551 ;
      RECT MASK 2 76.361 52.459 76.481 57.551 ;
      RECT MASK 2 76.801 52.459 76.921 57.551 ;
      RECT MASK 2 77.699 52.459 77.819 57.551 ;
      RECT MASK 2 78.139 52.459 78.259 57.551 ;
      RECT MASK 2 78.579 52.459 78.699 57.551 ;
      RECT MASK 2 79.019 52.459 79.139 57.551 ;
      RECT MASK 2 79.459 52.459 79.579 57.551 ;
      RECT MASK 2 79.899 52.459 80.019 57.551 ;
      RECT MASK 2 80.339 52.459 80.459 57.551 ;
      RECT MASK 2 80.779 52.459 80.899 57.551 ;
      RECT MASK 2 81.219 52.459 81.339 57.551 ;
      RECT MASK 2 81.659 52.459 81.779 57.551 ;
      RECT MASK 2 82.099 52.459 82.219 57.551 ;
      RECT MASK 2 82.539 52.459 82.659 57.551 ;
      RECT MASK 2 82.979 52.459 83.099 57.551 ;
      RECT MASK 2 83.419 52.459 83.539 57.551 ;
      RECT MASK 2 84.317 52.459 84.437 57.551 ;
      RECT MASK 2 84.757 52.459 84.877 57.551 ;
      RECT MASK 2 85.197 52.459 85.317 57.551 ;
      RECT MASK 2 85.637 52.459 85.757 57.551 ;
      RECT MASK 2 86.077 52.459 86.197 57.551 ;
      RECT MASK 2 86.517 52.459 86.637 57.551 ;
      RECT MASK 2 86.957 52.459 87.077 57.551 ;
      RECT MASK 2 87.397 52.459 87.517 57.551 ;
      RECT MASK 2 87.837 52.459 87.957 57.551 ;
      RECT MASK 2 88.277 52.459 88.397 57.551 ;
      RECT MASK 2 88.717 52.459 88.837 57.551 ;
      RECT MASK 2 89.157 52.459 89.277 57.551 ;
      RECT MASK 2 89.597 52.459 89.717 57.551 ;
      RECT MASK 2 90.037 52.459 90.157 57.551 ;
      RECT MASK 2 90.935 52.459 91.055 57.551 ;
      RECT MASK 2 91.375 52.459 91.495 57.551 ;
      RECT MASK 2 91.815 52.459 91.935 57.551 ;
      RECT MASK 2 92.255 52.459 92.375 57.551 ;
      RECT MASK 2 92.695 52.459 92.815 57.551 ;
      RECT MASK 2 93.135 52.459 93.255 57.551 ;
      RECT MASK 2 93.575 52.459 93.695 57.551 ;
      RECT MASK 2 94.015 52.459 94.135 57.551 ;
      RECT MASK 2 94.455 52.459 94.575 57.551 ;
      RECT MASK 2 94.895 52.459 95.015 57.551 ;
      RECT MASK 2 95.335 52.459 95.455 57.551 ;
      RECT MASK 2 95.775 52.459 95.895 57.551 ;
      RECT MASK 2 96.215 52.459 96.335 57.551 ;
      RECT MASK 2 96.655 52.459 96.775 57.551 ;
      RECT MASK 2 97.553 52.459 97.673 57.551 ;
      RECT MASK 2 97.993 52.459 98.113 57.551 ;
      RECT MASK 2 98.433 52.459 98.553 57.551 ;
      RECT MASK 2 98.873 52.459 98.993 57.551 ;
      RECT MASK 2 99.313 52.459 99.433 57.551 ;
      RECT MASK 2 99.753 52.459 99.873 57.551 ;
      RECT MASK 2 100.193 52.459 100.313 57.551 ;
      RECT MASK 2 100.633 52.459 100.753 57.551 ;
      RECT MASK 2 101.073 52.459 101.193 57.551 ;
      RECT MASK 2 101.513 52.459 101.633 57.551 ;
      RECT MASK 2 101.953 52.459 102.073 57.551 ;
      RECT MASK 2 102.393 52.459 102.513 57.551 ;
      RECT MASK 2 102.833 52.459 102.953 57.551 ;
      RECT MASK 2 103.273 52.459 103.393 57.551 ;
      RECT MASK 2 104.171 52.459 104.291 57.551 ;
      RECT MASK 2 104.611 52.459 104.731 57.551 ;
      RECT MASK 2 105.051 52.459 105.171 57.551 ;
      RECT MASK 2 105.491 52.459 105.611 57.551 ;
      RECT MASK 2 105.931 52.459 106.051 57.551 ;
      RECT MASK 2 106.371 52.459 106.491 57.551 ;
      RECT MASK 2 106.811 52.459 106.931 57.551 ;
      RECT MASK 2 107.251 52.459 107.371 57.551 ;
      RECT MASK 2 107.691 52.459 107.811 57.551 ;
      RECT MASK 2 108.131 52.459 108.251 57.551 ;
      RECT MASK 2 108.571 52.459 108.691 57.551 ;
      RECT MASK 2 109.011 52.459 109.131 57.551 ;
      RECT MASK 2 109.451 52.459 109.571 57.551 ;
      RECT MASK 2 109.891 52.459 110.011 57.551 ;
      RECT MASK 2 112.5865 53.149 112.7065 54.179 ;
      RECT MASK 2 113.0265 53.149 113.1465 54.179 ;
      RECT MASK 2 113.4665 53.149 113.5865 54.179 ;
      RECT MASK 2 113.9065 53.149 114.0265 54.179 ;
      RECT MASK 2 114.3465 53.149 114.4665 54.179 ;
      RECT MASK 2 114.7865 53.149 114.9065 54.179 ;
      RECT MASK 2 115.2265 53.149 115.3465 54.179 ;
      RECT MASK 2 115.6665 53.149 115.7865 54.179 ;
      RECT MASK 2 116.1065 53.149 116.2265 54.179 ;
      RECT MASK 2 116.5465 53.149 116.6665 54.179 ;
      RECT MASK 2 117.4265 54.41 117.5465 55.78 ;
      RECT MASK 2 117.8665 54.41 117.9865 55.78 ;
      RECT MASK 2 118.3065 54.41 118.4265 55.78 ;
      RECT MASK 2 118.7465 54.41 118.8665 55.78 ;
      RECT MASK 2 119.1865 54.41 119.3065 55.78 ;
      RECT MASK 2 119.6265 54.41 119.7465 55.78 ;
      RECT MASK 2 120.0665 54.41 120.1865 55.78 ;
      RECT MASK 2 120.5065 54.41 120.6265 55.78 ;
      RECT MASK 2 120.9465 54.41 121.0665 55.78 ;
      RECT MASK 2 121.3865 54.41 121.5065 55.78 ;
      RECT MASK 2 121.8265 54.41 121.9465 55.78 ;
      RECT MASK 2 122.2665 54.41 122.3865 55.78 ;
      RECT MASK 2 122.7065 54.41 122.8265 55.78 ;
      RECT MASK 2 123.1465 54.41 123.2665 55.78 ;
      RECT MASK 2 112.5865 54.499 112.7065 55.529 ;
      RECT MASK 2 113.0265 54.499 113.1465 55.529 ;
      RECT MASK 2 113.4665 54.499 113.5865 55.529 ;
      RECT MASK 2 113.9065 54.499 114.0265 55.529 ;
      RECT MASK 2 114.3465 54.499 114.4665 55.529 ;
      RECT MASK 2 114.7865 54.499 114.9065 55.529 ;
      RECT MASK 2 115.2265 54.499 115.3465 55.529 ;
      RECT MASK 2 115.6665 54.499 115.7865 55.529 ;
      RECT MASK 2 116.1065 54.499 116.2265 55.529 ;
      RECT MASK 2 116.5465 54.499 116.6665 55.529 ;
      RECT MASK 2 112.5865 55.789 112.7065 56.879 ;
      RECT MASK 2 113.0265 55.789 113.1465 56.879 ;
      RECT MASK 2 113.4665 55.789 113.5865 56.879 ;
      RECT MASK 2 113.9065 55.789 114.0265 56.879 ;
      RECT MASK 2 114.3465 55.789 114.4665 56.879 ;
      RECT MASK 2 114.7865 55.789 114.9065 56.879 ;
      RECT MASK 2 115.2265 55.789 115.3465 56.879 ;
      RECT MASK 2 115.6665 55.789 115.7865 56.879 ;
      RECT MASK 2 116.1065 55.789 116.2265 56.879 ;
      RECT MASK 2 116.5465 55.789 116.6665 56.879 ;
      RECT MASK 2 123.5865 55.849 123.7065 56.879 ;
      RECT MASK 2 112.5865 57.139 112.7065 58.949 ;
      RECT MASK 2 113.0265 57.139 113.1465 58.949 ;
      RECT MASK 2 113.4665 57.139 113.5865 58.949 ;
      RECT MASK 2 113.9065 57.139 114.0265 58.949 ;
      RECT MASK 2 114.3465 57.139 114.4665 58.949 ;
      RECT MASK 2 114.7865 57.139 114.9065 58.949 ;
      RECT MASK 2 115.2265 57.139 115.3465 58.949 ;
      RECT MASK 2 115.6665 57.139 115.7865 58.949 ;
      RECT MASK 2 116.1065 57.139 116.2265 58.949 ;
      RECT MASK 2 116.5465 57.139 116.6665 58.949 ;
      RECT MASK 2 117.4265 57.199 117.5465 58.949 ;
      RECT MASK 2 117.8665 57.199 117.9865 58.949 ;
      RECT MASK 2 118.3065 57.199 118.4265 58.949 ;
      RECT MASK 2 118.7465 57.199 118.8665 58.949 ;
      RECT MASK 2 119.1865 57.199 119.3065 58.949 ;
      RECT MASK 2 119.6265 57.199 119.7465 58.949 ;
      RECT MASK 2 120.0665 57.199 120.1865 58.949 ;
      RECT MASK 2 120.5065 57.199 120.6265 58.949 ;
      RECT MASK 2 120.9465 57.199 121.0665 58.949 ;
      RECT MASK 2 121.3865 57.199 121.5065 58.949 ;
      RECT MASK 2 121.8265 57.199 121.9465 58.949 ;
      RECT MASK 2 122.2665 57.199 122.3865 58.949 ;
      RECT MASK 2 122.7065 57.199 122.8265 58.949 ;
      RECT MASK 2 123.1465 57.199 123.2665 58.949 ;
      RECT MASK 2 123.5865 57.199 123.7065 58.949 ;
      RECT MASK 2 4.931 57.72 4.991 57.96 ;
      RECT MASK 2 5.371 57.72 5.431 57.96 ;
      RECT MASK 2 5.811 57.72 5.871 57.96 ;
      RECT MASK 2 6.251 57.72 6.311 57.96 ;
      RECT MASK 2 6.691 57.72 6.751 57.96 ;
      RECT MASK 2 7.131 57.72 7.191 57.96 ;
      RECT MASK 2 7.571 57.72 7.631 57.96 ;
      RECT MASK 2 8.011 57.72 8.071 57.96 ;
      RECT MASK 2 8.451 57.72 8.511 57.96 ;
      RECT MASK 2 8.891 57.72 8.951 57.96 ;
      RECT MASK 2 9.331 57.72 9.391 57.96 ;
      RECT MASK 2 9.771 57.72 9.831 57.96 ;
      RECT MASK 2 10.211 57.72 10.271 57.96 ;
      RECT MASK 2 10.651 57.72 10.711 57.96 ;
      RECT MASK 2 11.549 57.72 11.609 57.96 ;
      RECT MASK 2 11.989 57.72 12.049 57.96 ;
      RECT MASK 2 12.429 57.72 12.489 57.96 ;
      RECT MASK 2 12.869 57.72 12.929 57.96 ;
      RECT MASK 2 13.309 57.72 13.369 57.96 ;
      RECT MASK 2 13.749 57.72 13.809 57.96 ;
      RECT MASK 2 14.189 57.72 14.249 57.96 ;
      RECT MASK 2 14.629 57.72 14.689 57.96 ;
      RECT MASK 2 15.069 57.72 15.129 57.96 ;
      RECT MASK 2 15.509 57.72 15.569 57.96 ;
      RECT MASK 2 15.949 57.72 16.009 57.96 ;
      RECT MASK 2 16.389 57.72 16.449 57.96 ;
      RECT MASK 2 16.829 57.72 16.889 57.96 ;
      RECT MASK 2 17.269 57.72 17.329 57.96 ;
      RECT MASK 2 18.167 57.72 18.227 57.96 ;
      RECT MASK 2 18.607 57.72 18.667 57.96 ;
      RECT MASK 2 19.047 57.72 19.107 57.96 ;
      RECT MASK 2 19.487 57.72 19.547 57.96 ;
      RECT MASK 2 19.927 57.72 19.987 57.96 ;
      RECT MASK 2 20.367 57.72 20.427 57.96 ;
      RECT MASK 2 20.807 57.72 20.867 57.96 ;
      RECT MASK 2 21.247 57.72 21.307 57.96 ;
      RECT MASK 2 21.687 57.72 21.747 57.96 ;
      RECT MASK 2 22.127 57.72 22.187 57.96 ;
      RECT MASK 2 22.567 57.72 22.627 57.96 ;
      RECT MASK 2 23.007 57.72 23.067 57.96 ;
      RECT MASK 2 23.447 57.72 23.507 57.96 ;
      RECT MASK 2 23.887 57.72 23.947 57.96 ;
      RECT MASK 2 24.785 57.72 24.845 57.96 ;
      RECT MASK 2 25.225 57.72 25.285 57.96 ;
      RECT MASK 2 25.665 57.72 25.725 57.96 ;
      RECT MASK 2 26.105 57.72 26.165 57.96 ;
      RECT MASK 2 26.545 57.72 26.605 57.96 ;
      RECT MASK 2 26.985 57.72 27.045 57.96 ;
      RECT MASK 2 27.425 57.72 27.485 57.96 ;
      RECT MASK 2 27.865 57.72 27.925 57.96 ;
      RECT MASK 2 28.305 57.72 28.365 57.96 ;
      RECT MASK 2 28.745 57.72 28.805 57.96 ;
      RECT MASK 2 29.185 57.72 29.245 57.96 ;
      RECT MASK 2 29.625 57.72 29.685 57.96 ;
      RECT MASK 2 30.065 57.72 30.125 57.96 ;
      RECT MASK 2 30.505 57.72 30.565 57.96 ;
      RECT MASK 2 31.403 57.72 31.463 57.96 ;
      RECT MASK 2 31.843 57.72 31.903 57.96 ;
      RECT MASK 2 32.283 57.72 32.343 57.96 ;
      RECT MASK 2 32.723 57.72 32.783 57.96 ;
      RECT MASK 2 33.163 57.72 33.223 57.96 ;
      RECT MASK 2 33.603 57.72 33.663 57.96 ;
      RECT MASK 2 34.043 57.72 34.103 57.96 ;
      RECT MASK 2 34.483 57.72 34.543 57.96 ;
      RECT MASK 2 34.923 57.72 34.983 57.96 ;
      RECT MASK 2 35.363 57.72 35.423 57.96 ;
      RECT MASK 2 35.803 57.72 35.863 57.96 ;
      RECT MASK 2 36.243 57.72 36.303 57.96 ;
      RECT MASK 2 36.683 57.72 36.743 57.96 ;
      RECT MASK 2 37.123 57.72 37.183 57.96 ;
      RECT MASK 2 38.021 57.72 38.081 57.96 ;
      RECT MASK 2 38.461 57.72 38.521 57.96 ;
      RECT MASK 2 38.901 57.72 38.961 57.96 ;
      RECT MASK 2 39.341 57.72 39.401 57.96 ;
      RECT MASK 2 39.781 57.72 39.841 57.96 ;
      RECT MASK 2 40.221 57.72 40.281 57.96 ;
      RECT MASK 2 40.661 57.72 40.721 57.96 ;
      RECT MASK 2 41.101 57.72 41.161 57.96 ;
      RECT MASK 2 41.541 57.72 41.601 57.96 ;
      RECT MASK 2 42.861 57.72 42.921 57.96 ;
      RECT MASK 2 43.301 57.72 43.361 57.96 ;
      RECT MASK 2 43.741 57.72 43.801 57.96 ;
      RECT MASK 2 44.639 57.72 44.699 57.96 ;
      RECT MASK 2 45.079 57.72 45.139 57.96 ;
      RECT MASK 2 45.519 57.72 45.579 57.96 ;
      RECT MASK 2 45.959 57.72 46.019 57.96 ;
      RECT MASK 2 46.399 57.72 46.459 57.96 ;
      RECT MASK 2 46.839 57.72 46.899 57.96 ;
      RECT MASK 2 47.279 57.72 47.339 57.96 ;
      RECT MASK 2 47.719 57.72 47.779 57.96 ;
      RECT MASK 2 48.159 57.72 48.219 57.96 ;
      RECT MASK 2 48.599 57.72 48.659 57.96 ;
      RECT MASK 2 49.039 57.72 49.099 57.96 ;
      RECT MASK 2 49.479 57.72 49.539 57.96 ;
      RECT MASK 2 49.919 57.72 49.979 57.96 ;
      RECT MASK 2 50.359 57.72 50.419 57.96 ;
      RECT MASK 2 51.257 57.72 51.317 57.96 ;
      RECT MASK 2 51.697 57.72 51.757 57.96 ;
      RECT MASK 2 52.137 57.72 52.197 57.96 ;
      RECT MASK 2 52.577 57.72 52.637 57.96 ;
      RECT MASK 2 53.017 57.72 53.077 57.96 ;
      RECT MASK 2 53.457 57.72 53.517 57.96 ;
      RECT MASK 2 53.897 57.72 53.957 57.96 ;
      RECT MASK 2 54.337 57.72 54.397 57.96 ;
      RECT MASK 2 54.777 57.72 54.837 57.96 ;
      RECT MASK 2 55.217 57.72 55.277 57.96 ;
      RECT MASK 2 55.657 57.72 55.717 57.96 ;
      RECT MASK 2 56.097 57.72 56.157 57.96 ;
      RECT MASK 2 56.537 57.72 56.597 57.96 ;
      RECT MASK 2 56.977 57.72 57.037 57.96 ;
      RECT MASK 2 57.875 57.72 57.935 57.96 ;
      RECT MASK 2 58.315 57.72 58.375 57.96 ;
      RECT MASK 2 58.755 57.72 58.815 57.96 ;
      RECT MASK 2 59.195 57.72 59.255 57.96 ;
      RECT MASK 2 59.635 57.72 59.695 57.96 ;
      RECT MASK 2 60.075 57.72 60.135 57.96 ;
      RECT MASK 2 60.515 57.72 60.575 57.96 ;
      RECT MASK 2 60.955 57.72 61.015 57.96 ;
      RECT MASK 2 61.395 57.72 61.455 57.96 ;
      RECT MASK 2 61.835 57.72 61.895 57.96 ;
      RECT MASK 2 62.275 57.72 62.335 57.96 ;
      RECT MASK 2 62.715 57.72 62.775 57.96 ;
      RECT MASK 2 63.155 57.72 63.215 57.96 ;
      RECT MASK 2 63.595 57.72 63.655 57.96 ;
      RECT MASK 2 64.493 57.72 64.553 57.96 ;
      RECT MASK 2 64.933 57.72 64.993 57.96 ;
      RECT MASK 2 65.373 57.72 65.433 57.96 ;
      RECT MASK 2 65.813 57.72 65.873 57.96 ;
      RECT MASK 2 66.253 57.72 66.313 57.96 ;
      RECT MASK 2 66.693 57.72 66.753 57.96 ;
      RECT MASK 2 67.133 57.72 67.193 57.96 ;
      RECT MASK 2 67.573 57.72 67.633 57.96 ;
      RECT MASK 2 68.013 57.72 68.073 57.96 ;
      RECT MASK 2 68.453 57.72 68.513 57.96 ;
      RECT MASK 2 68.893 57.72 68.953 57.96 ;
      RECT MASK 2 69.333 57.72 69.393 57.96 ;
      RECT MASK 2 69.773 57.72 69.833 57.96 ;
      RECT MASK 2 70.213 57.72 70.273 57.96 ;
      RECT MASK 2 71.111 57.72 71.171 57.96 ;
      RECT MASK 2 71.551 57.72 71.611 57.96 ;
      RECT MASK 2 71.991 57.72 72.051 57.96 ;
      RECT MASK 2 72.431 57.72 72.491 57.96 ;
      RECT MASK 2 72.871 57.72 72.931 57.96 ;
      RECT MASK 2 73.311 57.72 73.371 57.96 ;
      RECT MASK 2 73.751 57.72 73.811 57.96 ;
      RECT MASK 2 74.191 57.72 74.251 57.96 ;
      RECT MASK 2 74.631 57.72 74.691 57.96 ;
      RECT MASK 2 75.071 57.72 75.131 57.96 ;
      RECT MASK 2 75.511 57.72 75.571 57.96 ;
      RECT MASK 2 75.951 57.72 76.011 57.96 ;
      RECT MASK 2 76.391 57.72 76.451 57.96 ;
      RECT MASK 2 76.831 57.72 76.891 57.96 ;
      RECT MASK 2 77.729 57.72 77.789 57.96 ;
      RECT MASK 2 78.169 57.72 78.229 57.96 ;
      RECT MASK 2 78.609 57.72 78.669 57.96 ;
      RECT MASK 2 79.049 57.72 79.109 57.96 ;
      RECT MASK 2 79.489 57.72 79.549 57.96 ;
      RECT MASK 2 79.929 57.72 79.989 57.96 ;
      RECT MASK 2 80.369 57.72 80.429 57.96 ;
      RECT MASK 2 80.809 57.72 80.869 57.96 ;
      RECT MASK 2 81.249 57.72 81.309 57.96 ;
      RECT MASK 2 81.689 57.72 81.749 57.96 ;
      RECT MASK 2 82.129 57.72 82.189 57.96 ;
      RECT MASK 2 83.449 57.72 83.509 57.96 ;
      RECT MASK 2 84.347 57.72 84.407 57.96 ;
      RECT MASK 2 84.787 57.72 84.847 57.96 ;
      RECT MASK 2 85.227 57.72 85.287 57.96 ;
      RECT MASK 2 85.667 57.72 85.727 57.96 ;
      RECT MASK 2 86.107 57.72 86.167 57.96 ;
      RECT MASK 2 86.547 57.72 86.607 57.96 ;
      RECT MASK 2 86.987 57.72 87.047 57.96 ;
      RECT MASK 2 87.427 57.72 87.487 57.96 ;
      RECT MASK 2 87.867 57.72 87.927 57.96 ;
      RECT MASK 2 88.307 57.72 88.367 57.96 ;
      RECT MASK 2 88.747 57.72 88.807 57.96 ;
      RECT MASK 2 89.187 57.72 89.247 57.96 ;
      RECT MASK 2 89.627 57.72 89.687 57.96 ;
      RECT MASK 2 90.067 57.72 90.127 57.96 ;
      RECT MASK 2 90.965 57.72 91.025 57.96 ;
      RECT MASK 2 91.405 57.72 91.465 57.96 ;
      RECT MASK 2 91.845 57.72 91.905 57.96 ;
      RECT MASK 2 92.285 57.72 92.345 57.96 ;
      RECT MASK 2 92.725 57.72 92.785 57.96 ;
      RECT MASK 2 93.165 57.72 93.225 57.96 ;
      RECT MASK 2 93.605 57.72 93.665 57.96 ;
      RECT MASK 2 94.045 57.72 94.105 57.96 ;
      RECT MASK 2 94.485 57.72 94.545 57.96 ;
      RECT MASK 2 94.925 57.72 94.985 57.96 ;
      RECT MASK 2 95.365 57.72 95.425 57.96 ;
      RECT MASK 2 95.805 57.72 95.865 57.96 ;
      RECT MASK 2 96.245 57.72 96.305 57.96 ;
      RECT MASK 2 96.685 57.72 96.745 57.96 ;
      RECT MASK 2 97.583 57.72 97.643 57.96 ;
      RECT MASK 2 98.023 57.72 98.083 57.96 ;
      RECT MASK 2 98.463 57.72 98.523 57.96 ;
      RECT MASK 2 98.903 57.72 98.963 57.96 ;
      RECT MASK 2 99.343 57.72 99.403 57.96 ;
      RECT MASK 2 99.783 57.72 99.843 57.96 ;
      RECT MASK 2 100.223 57.72 100.283 57.96 ;
      RECT MASK 2 100.663 57.72 100.723 57.96 ;
      RECT MASK 2 101.103 57.72 101.163 57.96 ;
      RECT MASK 2 101.543 57.72 101.603 57.96 ;
      RECT MASK 2 101.983 57.72 102.043 57.96 ;
      RECT MASK 2 102.423 57.72 102.483 57.96 ;
      RECT MASK 2 102.863 57.72 102.923 57.96 ;
      RECT MASK 2 103.303 57.72 103.363 57.96 ;
      RECT MASK 2 104.201 57.72 104.261 57.96 ;
      RECT MASK 2 104.641 57.72 104.701 57.96 ;
      RECT MASK 2 105.081 57.72 105.141 57.96 ;
      RECT MASK 2 105.521 57.72 105.581 57.96 ;
      RECT MASK 2 105.961 57.72 106.021 57.96 ;
      RECT MASK 2 106.401 57.72 106.461 57.96 ;
      RECT MASK 2 106.841 57.72 106.901 57.96 ;
      RECT MASK 2 107.281 57.72 107.341 57.96 ;
      RECT MASK 2 107.721 57.72 107.781 57.96 ;
      RECT MASK 2 108.161 57.72 108.221 57.96 ;
      RECT MASK 2 108.601 57.72 108.661 57.96 ;
      RECT MASK 2 109.041 57.72 109.101 57.96 ;
      RECT MASK 2 109.481 57.72 109.541 57.96 ;
      RECT MASK 2 109.921 57.72 109.981 57.96 ;
      RECT MASK 2 4.931 58.14 4.991 58.38 ;
      RECT MASK 2 5.371 58.14 5.431 58.38 ;
      RECT MASK 2 5.811 58.14 5.871 58.38 ;
      RECT MASK 2 6.251 58.14 6.311 58.38 ;
      RECT MASK 2 6.691 58.14 6.751 58.38 ;
      RECT MASK 2 7.131 58.14 7.191 58.38 ;
      RECT MASK 2 7.571 58.14 7.631 58.38 ;
      RECT MASK 2 8.011 58.14 8.071 58.38 ;
      RECT MASK 2 8.451 58.14 8.511 58.38 ;
      RECT MASK 2 8.891 58.14 8.951 58.38 ;
      RECT MASK 2 9.331 58.14 9.391 58.38 ;
      RECT MASK 2 9.771 58.14 9.831 58.38 ;
      RECT MASK 2 10.211 58.14 10.271 58.38 ;
      RECT MASK 2 10.651 58.14 10.711 58.38 ;
      RECT MASK 2 11.549 58.14 11.609 58.38 ;
      RECT MASK 2 11.989 58.14 12.049 58.38 ;
      RECT MASK 2 12.429 58.14 12.489 58.38 ;
      RECT MASK 2 12.869 58.14 12.929 58.38 ;
      RECT MASK 2 13.309 58.14 13.369 58.38 ;
      RECT MASK 2 13.749 58.14 13.809 58.38 ;
      RECT MASK 2 14.189 58.14 14.249 58.38 ;
      RECT MASK 2 14.629 58.14 14.689 58.38 ;
      RECT MASK 2 15.069 58.14 15.129 58.38 ;
      RECT MASK 2 15.509 58.14 15.569 58.38 ;
      RECT MASK 2 15.949 58.14 16.009 58.38 ;
      RECT MASK 2 16.389 58.14 16.449 58.38 ;
      RECT MASK 2 16.829 58.14 16.889 58.38 ;
      RECT MASK 2 17.269 58.14 17.329 58.38 ;
      RECT MASK 2 18.167 58.14 18.227 58.38 ;
      RECT MASK 2 18.607 58.14 18.667 58.38 ;
      RECT MASK 2 19.047 58.14 19.107 58.38 ;
      RECT MASK 2 19.487 58.14 19.547 58.38 ;
      RECT MASK 2 19.927 58.14 19.987 58.38 ;
      RECT MASK 2 20.367 58.14 20.427 58.38 ;
      RECT MASK 2 20.807 58.14 20.867 58.38 ;
      RECT MASK 2 21.247 58.14 21.307 58.38 ;
      RECT MASK 2 21.687 58.14 21.747 58.38 ;
      RECT MASK 2 22.127 58.14 22.187 58.38 ;
      RECT MASK 2 22.567 58.14 22.627 58.38 ;
      RECT MASK 2 23.007 58.14 23.067 58.38 ;
      RECT MASK 2 23.447 58.14 23.507 58.38 ;
      RECT MASK 2 23.887 58.14 23.947 58.38 ;
      RECT MASK 2 24.785 58.14 24.845 58.38 ;
      RECT MASK 2 25.225 58.14 25.285 58.38 ;
      RECT MASK 2 25.665 58.14 25.725 58.38 ;
      RECT MASK 2 26.105 58.14 26.165 58.38 ;
      RECT MASK 2 26.545 58.14 26.605 58.38 ;
      RECT MASK 2 26.985 58.14 27.045 58.38 ;
      RECT MASK 2 27.425 58.14 27.485 58.38 ;
      RECT MASK 2 27.865 58.14 27.925 58.38 ;
      RECT MASK 2 28.305 58.14 28.365 58.38 ;
      RECT MASK 2 28.745 58.14 28.805 58.38 ;
      RECT MASK 2 29.185 58.14 29.245 58.38 ;
      RECT MASK 2 29.625 58.14 29.685 58.38 ;
      RECT MASK 2 30.065 58.14 30.125 58.38 ;
      RECT MASK 2 30.505 58.14 30.565 58.38 ;
      RECT MASK 2 31.403 58.14 31.463 58.38 ;
      RECT MASK 2 31.843 58.14 31.903 58.38 ;
      RECT MASK 2 32.283 58.14 32.343 58.38 ;
      RECT MASK 2 32.723 58.14 32.783 58.38 ;
      RECT MASK 2 33.163 58.14 33.223 58.38 ;
      RECT MASK 2 33.603 58.14 33.663 58.38 ;
      RECT MASK 2 34.043 58.14 34.103 58.38 ;
      RECT MASK 2 34.483 58.14 34.543 58.38 ;
      RECT MASK 2 34.923 58.14 34.983 58.38 ;
      RECT MASK 2 35.363 58.14 35.423 58.38 ;
      RECT MASK 2 35.803 58.14 35.863 58.38 ;
      RECT MASK 2 36.243 58.14 36.303 58.38 ;
      RECT MASK 2 36.683 58.14 36.743 58.38 ;
      RECT MASK 2 37.123 58.14 37.183 58.38 ;
      RECT MASK 2 38.021 58.14 38.081 58.38 ;
      RECT MASK 2 38.461 58.14 38.521 58.38 ;
      RECT MASK 2 38.901 58.14 38.961 58.38 ;
      RECT MASK 2 39.341 58.14 39.401 58.38 ;
      RECT MASK 2 39.781 58.14 39.841 58.38 ;
      RECT MASK 2 40.221 58.14 40.281 58.38 ;
      RECT MASK 2 40.661 58.14 40.721 58.38 ;
      RECT MASK 2 41.101 58.14 41.161 58.38 ;
      RECT MASK 2 41.541 58.14 41.601 58.38 ;
      RECT MASK 2 42.861 58.14 42.921 58.38 ;
      RECT MASK 2 43.301 58.14 43.361 58.38 ;
      RECT MASK 2 43.741 58.14 43.801 58.38 ;
      RECT MASK 2 44.639 58.14 44.699 58.38 ;
      RECT MASK 2 45.079 58.14 45.139 58.38 ;
      RECT MASK 2 45.519 58.14 45.579 58.38 ;
      RECT MASK 2 45.959 58.14 46.019 58.38 ;
      RECT MASK 2 46.399 58.14 46.459 58.38 ;
      RECT MASK 2 46.839 58.14 46.899 58.38 ;
      RECT MASK 2 47.279 58.14 47.339 58.38 ;
      RECT MASK 2 47.719 58.14 47.779 58.38 ;
      RECT MASK 2 48.159 58.14 48.219 58.38 ;
      RECT MASK 2 48.599 58.14 48.659 58.38 ;
      RECT MASK 2 49.039 58.14 49.099 58.38 ;
      RECT MASK 2 49.479 58.14 49.539 58.38 ;
      RECT MASK 2 49.919 58.14 49.979 58.38 ;
      RECT MASK 2 50.359 58.14 50.419 58.38 ;
      RECT MASK 2 51.257 58.14 51.317 58.38 ;
      RECT MASK 2 51.697 58.14 51.757 58.38 ;
      RECT MASK 2 52.137 58.14 52.197 58.38 ;
      RECT MASK 2 52.577 58.14 52.637 58.38 ;
      RECT MASK 2 53.017 58.14 53.077 58.38 ;
      RECT MASK 2 53.457 58.14 53.517 58.38 ;
      RECT MASK 2 53.897 58.14 53.957 58.38 ;
      RECT MASK 2 54.337 58.14 54.397 58.38 ;
      RECT MASK 2 54.777 58.14 54.837 58.38 ;
      RECT MASK 2 55.217 58.14 55.277 58.38 ;
      RECT MASK 2 55.657 58.14 55.717 58.38 ;
      RECT MASK 2 56.097 58.14 56.157 58.38 ;
      RECT MASK 2 56.537 58.14 56.597 58.38 ;
      RECT MASK 2 56.977 58.14 57.037 58.38 ;
      RECT MASK 2 57.875 58.14 57.935 58.38 ;
      RECT MASK 2 58.315 58.14 58.375 58.38 ;
      RECT MASK 2 58.755 58.14 58.815 58.38 ;
      RECT MASK 2 59.195 58.14 59.255 58.38 ;
      RECT MASK 2 59.635 58.14 59.695 58.38 ;
      RECT MASK 2 60.075 58.14 60.135 58.38 ;
      RECT MASK 2 60.515 58.14 60.575 58.38 ;
      RECT MASK 2 60.955 58.14 61.015 58.38 ;
      RECT MASK 2 61.395 58.14 61.455 58.38 ;
      RECT MASK 2 61.835 58.14 61.895 58.38 ;
      RECT MASK 2 62.275 58.14 62.335 58.38 ;
      RECT MASK 2 62.715 58.14 62.775 58.38 ;
      RECT MASK 2 63.155 58.14 63.215 58.38 ;
      RECT MASK 2 63.595 58.14 63.655 58.38 ;
      RECT MASK 2 64.493 58.14 64.553 58.38 ;
      RECT MASK 2 64.933 58.14 64.993 58.38 ;
      RECT MASK 2 65.373 58.14 65.433 58.38 ;
      RECT MASK 2 65.813 58.14 65.873 58.38 ;
      RECT MASK 2 66.253 58.14 66.313 58.38 ;
      RECT MASK 2 66.693 58.14 66.753 58.38 ;
      RECT MASK 2 67.133 58.14 67.193 58.38 ;
      RECT MASK 2 67.573 58.14 67.633 58.38 ;
      RECT MASK 2 68.013 58.14 68.073 58.38 ;
      RECT MASK 2 68.453 58.14 68.513 58.38 ;
      RECT MASK 2 68.893 58.14 68.953 58.38 ;
      RECT MASK 2 69.333 58.14 69.393 58.38 ;
      RECT MASK 2 69.773 58.14 69.833 58.38 ;
      RECT MASK 2 70.213 58.14 70.273 58.38 ;
      RECT MASK 2 71.111 58.14 71.171 58.38 ;
      RECT MASK 2 71.551 58.14 71.611 58.38 ;
      RECT MASK 2 71.991 58.14 72.051 58.38 ;
      RECT MASK 2 72.431 58.14 72.491 58.38 ;
      RECT MASK 2 72.871 58.14 72.931 58.38 ;
      RECT MASK 2 73.311 58.14 73.371 58.38 ;
      RECT MASK 2 73.751 58.14 73.811 58.38 ;
      RECT MASK 2 74.191 58.14 74.251 58.38 ;
      RECT MASK 2 74.631 58.14 74.691 58.38 ;
      RECT MASK 2 75.071 58.14 75.131 58.38 ;
      RECT MASK 2 75.511 58.14 75.571 58.38 ;
      RECT MASK 2 75.951 58.14 76.011 58.38 ;
      RECT MASK 2 76.391 58.14 76.451 58.38 ;
      RECT MASK 2 76.831 58.14 76.891 58.38 ;
      RECT MASK 2 77.729 58.14 77.789 58.38 ;
      RECT MASK 2 78.169 58.14 78.229 58.38 ;
      RECT MASK 2 78.609 58.14 78.669 58.38 ;
      RECT MASK 2 79.049 58.14 79.109 58.38 ;
      RECT MASK 2 79.489 58.14 79.549 58.38 ;
      RECT MASK 2 79.929 58.14 79.989 58.38 ;
      RECT MASK 2 80.369 58.14 80.429 58.38 ;
      RECT MASK 2 80.809 58.14 80.869 58.38 ;
      RECT MASK 2 81.249 58.14 81.309 58.38 ;
      RECT MASK 2 81.689 58.14 81.749 58.38 ;
      RECT MASK 2 82.129 58.14 82.189 58.38 ;
      RECT MASK 2 83.449 58.14 83.509 58.38 ;
      RECT MASK 2 84.347 58.14 84.407 58.38 ;
      RECT MASK 2 84.787 58.14 84.847 58.38 ;
      RECT MASK 2 85.227 58.14 85.287 58.38 ;
      RECT MASK 2 85.667 58.14 85.727 58.38 ;
      RECT MASK 2 86.107 58.14 86.167 58.38 ;
      RECT MASK 2 86.547 58.14 86.607 58.38 ;
      RECT MASK 2 86.987 58.14 87.047 58.38 ;
      RECT MASK 2 87.427 58.14 87.487 58.38 ;
      RECT MASK 2 87.867 58.14 87.927 58.38 ;
      RECT MASK 2 88.307 58.14 88.367 58.38 ;
      RECT MASK 2 88.747 58.14 88.807 58.38 ;
      RECT MASK 2 89.187 58.14 89.247 58.38 ;
      RECT MASK 2 89.627 58.14 89.687 58.38 ;
      RECT MASK 2 90.067 58.14 90.127 58.38 ;
      RECT MASK 2 90.965 58.14 91.025 58.38 ;
      RECT MASK 2 91.405 58.14 91.465 58.38 ;
      RECT MASK 2 91.845 58.14 91.905 58.38 ;
      RECT MASK 2 92.285 58.14 92.345 58.38 ;
      RECT MASK 2 92.725 58.14 92.785 58.38 ;
      RECT MASK 2 93.165 58.14 93.225 58.38 ;
      RECT MASK 2 93.605 58.14 93.665 58.38 ;
      RECT MASK 2 94.045 58.14 94.105 58.38 ;
      RECT MASK 2 94.485 58.14 94.545 58.38 ;
      RECT MASK 2 94.925 58.14 94.985 58.38 ;
      RECT MASK 2 95.365 58.14 95.425 58.38 ;
      RECT MASK 2 95.805 58.14 95.865 58.38 ;
      RECT MASK 2 96.245 58.14 96.305 58.38 ;
      RECT MASK 2 96.685 58.14 96.745 58.38 ;
      RECT MASK 2 97.583 58.14 97.643 58.38 ;
      RECT MASK 2 98.023 58.14 98.083 58.38 ;
      RECT MASK 2 98.463 58.14 98.523 58.38 ;
      RECT MASK 2 98.903 58.14 98.963 58.38 ;
      RECT MASK 2 99.343 58.14 99.403 58.38 ;
      RECT MASK 2 99.783 58.14 99.843 58.38 ;
      RECT MASK 2 100.223 58.14 100.283 58.38 ;
      RECT MASK 2 100.663 58.14 100.723 58.38 ;
      RECT MASK 2 101.103 58.14 101.163 58.38 ;
      RECT MASK 2 101.543 58.14 101.603 58.38 ;
      RECT MASK 2 101.983 58.14 102.043 58.38 ;
      RECT MASK 2 102.423 58.14 102.483 58.38 ;
      RECT MASK 2 102.863 58.14 102.923 58.38 ;
      RECT MASK 2 103.303 58.14 103.363 58.38 ;
      RECT MASK 2 104.201 58.14 104.261 58.38 ;
      RECT MASK 2 104.641 58.14 104.701 58.38 ;
      RECT MASK 2 105.081 58.14 105.141 58.38 ;
      RECT MASK 2 105.521 58.14 105.581 58.38 ;
      RECT MASK 2 105.961 58.14 106.021 58.38 ;
      RECT MASK 2 106.401 58.14 106.461 58.38 ;
      RECT MASK 2 106.841 58.14 106.901 58.38 ;
      RECT MASK 2 107.281 58.14 107.341 58.38 ;
      RECT MASK 2 107.721 58.14 107.781 58.38 ;
      RECT MASK 2 108.161 58.14 108.221 58.38 ;
      RECT MASK 2 108.601 58.14 108.661 58.38 ;
      RECT MASK 2 109.041 58.14 109.101 58.38 ;
      RECT MASK 2 109.481 58.14 109.541 58.38 ;
      RECT MASK 2 109.921 58.14 109.981 58.38 ;
      RECT MASK 2 4.901 58.579 5.021 69.791 ;
      RECT MASK 2 5.341 58.579 5.461 69.791 ;
      RECT MASK 2 5.781 58.579 5.901 69.791 ;
      RECT MASK 2 6.221 58.579 6.341 69.791 ;
      RECT MASK 2 6.661 58.579 6.781 69.791 ;
      RECT MASK 2 7.101 58.579 7.221 69.791 ;
      RECT MASK 2 7.541 58.579 7.661 69.791 ;
      RECT MASK 2 7.981 58.579 8.101 69.791 ;
      RECT MASK 2 8.421 58.579 8.541 69.791 ;
      RECT MASK 2 8.861 58.579 8.981 69.791 ;
      RECT MASK 2 9.301 58.579 9.421 69.791 ;
      RECT MASK 2 9.741 58.579 9.861 69.791 ;
      RECT MASK 2 10.181 58.579 10.301 69.791 ;
      RECT MASK 2 10.621 58.579 10.741 69.791 ;
      RECT MASK 2 11.519 58.579 11.639 69.791 ;
      RECT MASK 2 11.959 58.579 12.079 69.791 ;
      RECT MASK 2 12.399 58.579 12.519 69.791 ;
      RECT MASK 2 12.839 58.579 12.959 69.791 ;
      RECT MASK 2 13.279 58.579 13.399 69.791 ;
      RECT MASK 2 13.719 58.579 13.839 69.791 ;
      RECT MASK 2 14.159 58.579 14.279 69.791 ;
      RECT MASK 2 14.599 58.579 14.719 69.791 ;
      RECT MASK 2 15.039 58.579 15.159 69.791 ;
      RECT MASK 2 15.479 58.579 15.599 69.791 ;
      RECT MASK 2 15.919 58.579 16.039 69.791 ;
      RECT MASK 2 16.359 58.579 16.479 69.791 ;
      RECT MASK 2 16.799 58.579 16.919 69.791 ;
      RECT MASK 2 17.239 58.579 17.359 69.791 ;
      RECT MASK 2 18.137 58.579 18.257 69.791 ;
      RECT MASK 2 18.577 58.579 18.697 69.791 ;
      RECT MASK 2 19.017 58.579 19.137 69.791 ;
      RECT MASK 2 19.457 58.579 19.577 69.791 ;
      RECT MASK 2 19.897 58.579 20.017 69.791 ;
      RECT MASK 2 20.337 58.579 20.457 69.791 ;
      RECT MASK 2 20.777 58.579 20.897 69.791 ;
      RECT MASK 2 21.217 58.579 21.337 69.791 ;
      RECT MASK 2 21.657 58.579 21.777 69.791 ;
      RECT MASK 2 22.097 58.579 22.217 69.791 ;
      RECT MASK 2 22.537 58.579 22.657 69.791 ;
      RECT MASK 2 22.977 58.579 23.097 69.791 ;
      RECT MASK 2 23.417 58.579 23.537 69.791 ;
      RECT MASK 2 23.857 58.579 23.977 69.791 ;
      RECT MASK 2 24.755 58.579 24.875 69.791 ;
      RECT MASK 2 25.195 58.579 25.315 69.791 ;
      RECT MASK 2 25.635 58.579 25.755 69.791 ;
      RECT MASK 2 26.075 58.579 26.195 69.791 ;
      RECT MASK 2 26.515 58.579 26.635 69.791 ;
      RECT MASK 2 26.955 58.579 27.075 69.791 ;
      RECT MASK 2 27.395 58.579 27.515 69.791 ;
      RECT MASK 2 27.835 58.579 27.955 69.791 ;
      RECT MASK 2 28.275 58.579 28.395 69.791 ;
      RECT MASK 2 28.715 58.579 28.835 69.791 ;
      RECT MASK 2 29.155 58.579 29.275 69.791 ;
      RECT MASK 2 29.595 58.579 29.715 69.791 ;
      RECT MASK 2 30.035 58.579 30.155 69.791 ;
      RECT MASK 2 30.475 58.579 30.595 69.791 ;
      RECT MASK 2 31.373 58.579 31.493 69.791 ;
      RECT MASK 2 31.813 58.579 31.933 69.791 ;
      RECT MASK 2 32.253 58.579 32.373 69.791 ;
      RECT MASK 2 32.693 58.579 32.813 69.791 ;
      RECT MASK 2 33.133 58.579 33.253 69.791 ;
      RECT MASK 2 33.573 58.579 33.693 69.791 ;
      RECT MASK 2 34.013 58.579 34.133 69.791 ;
      RECT MASK 2 34.453 58.579 34.573 69.791 ;
      RECT MASK 2 34.893 58.579 35.013 69.791 ;
      RECT MASK 2 35.333 58.579 35.453 69.791 ;
      RECT MASK 2 35.773 58.579 35.893 69.791 ;
      RECT MASK 2 36.213 58.579 36.333 69.791 ;
      RECT MASK 2 36.653 58.579 36.773 69.791 ;
      RECT MASK 2 37.093 58.579 37.213 69.791 ;
      RECT MASK 2 37.991 58.579 38.111 69.791 ;
      RECT MASK 2 38.431 58.579 38.551 69.791 ;
      RECT MASK 2 38.871 58.579 38.991 69.791 ;
      RECT MASK 2 39.311 58.579 39.431 69.791 ;
      RECT MASK 2 39.751 58.579 39.871 69.791 ;
      RECT MASK 2 40.191 58.579 40.311 69.791 ;
      RECT MASK 2 40.631 58.579 40.751 69.791 ;
      RECT MASK 2 41.071 58.579 41.191 69.791 ;
      RECT MASK 2 41.511 58.579 41.631 69.791 ;
      RECT MASK 2 41.951 58.579 42.071 69.791 ;
      RECT MASK 2 42.391 58.579 42.511 69.791 ;
      RECT MASK 2 42.831 58.579 42.951 69.791 ;
      RECT MASK 2 43.271 58.579 43.391 69.791 ;
      RECT MASK 2 43.711 58.579 43.831 69.791 ;
      RECT MASK 2 44.609 58.579 44.729 69.791 ;
      RECT MASK 2 45.049 58.579 45.169 69.791 ;
      RECT MASK 2 45.489 58.579 45.609 69.791 ;
      RECT MASK 2 45.929 58.579 46.049 69.791 ;
      RECT MASK 2 46.369 58.579 46.489 69.791 ;
      RECT MASK 2 46.809 58.579 46.929 69.791 ;
      RECT MASK 2 47.249 58.579 47.369 69.791 ;
      RECT MASK 2 47.689 58.579 47.809 69.791 ;
      RECT MASK 2 48.129 58.579 48.249 69.791 ;
      RECT MASK 2 48.569 58.579 48.689 69.791 ;
      RECT MASK 2 49.009 58.579 49.129 69.791 ;
      RECT MASK 2 49.449 58.579 49.569 69.791 ;
      RECT MASK 2 49.889 58.579 50.009 69.791 ;
      RECT MASK 2 50.329 58.579 50.449 69.791 ;
      RECT MASK 2 51.227 58.579 51.347 69.791 ;
      RECT MASK 2 51.667 58.579 51.787 69.791 ;
      RECT MASK 2 52.107 58.579 52.227 69.791 ;
      RECT MASK 2 52.547 58.579 52.667 69.791 ;
      RECT MASK 2 52.987 58.579 53.107 69.791 ;
      RECT MASK 2 53.427 58.579 53.547 69.791 ;
      RECT MASK 2 53.867 58.579 53.987 69.791 ;
      RECT MASK 2 54.307 58.579 54.427 69.791 ;
      RECT MASK 2 54.747 58.579 54.867 69.791 ;
      RECT MASK 2 55.187 58.579 55.307 69.791 ;
      RECT MASK 2 55.627 58.579 55.747 69.791 ;
      RECT MASK 2 56.067 58.579 56.187 69.791 ;
      RECT MASK 2 56.507 58.579 56.627 69.791 ;
      RECT MASK 2 56.947 58.579 57.067 69.791 ;
      RECT MASK 2 57.845 58.579 57.965 69.791 ;
      RECT MASK 2 58.285 58.579 58.405 69.791 ;
      RECT MASK 2 58.725 58.579 58.845 69.791 ;
      RECT MASK 2 59.165 58.579 59.285 69.791 ;
      RECT MASK 2 59.605 58.579 59.725 69.791 ;
      RECT MASK 2 60.045 58.579 60.165 69.791 ;
      RECT MASK 2 60.485 58.579 60.605 69.791 ;
      RECT MASK 2 60.925 58.579 61.045 69.791 ;
      RECT MASK 2 61.365 58.579 61.485 69.791 ;
      RECT MASK 2 61.805 58.579 61.925 69.791 ;
      RECT MASK 2 62.245 58.579 62.365 69.791 ;
      RECT MASK 2 62.685 58.579 62.805 69.791 ;
      RECT MASK 2 63.125 58.579 63.245 69.791 ;
      RECT MASK 2 63.565 58.579 63.685 69.791 ;
      RECT MASK 2 64.463 58.579 64.583 69.791 ;
      RECT MASK 2 64.903 58.579 65.023 69.791 ;
      RECT MASK 2 65.343 58.579 65.463 69.791 ;
      RECT MASK 2 65.783 58.579 65.903 69.791 ;
      RECT MASK 2 66.223 58.579 66.343 69.791 ;
      RECT MASK 2 66.663 58.579 66.783 69.791 ;
      RECT MASK 2 67.103 58.579 67.223 69.791 ;
      RECT MASK 2 67.543 58.579 67.663 69.791 ;
      RECT MASK 2 67.983 58.579 68.103 69.791 ;
      RECT MASK 2 68.423 58.579 68.543 69.791 ;
      RECT MASK 2 68.863 58.579 68.983 69.791 ;
      RECT MASK 2 69.303 58.579 69.423 69.791 ;
      RECT MASK 2 69.743 58.579 69.863 69.791 ;
      RECT MASK 2 70.183 58.579 70.303 69.791 ;
      RECT MASK 2 71.081 58.579 71.201 69.791 ;
      RECT MASK 2 71.521 58.579 71.641 69.791 ;
      RECT MASK 2 71.961 58.579 72.081 69.791 ;
      RECT MASK 2 72.401 58.579 72.521 69.791 ;
      RECT MASK 2 72.841 58.579 72.961 69.791 ;
      RECT MASK 2 73.281 58.579 73.401 69.791 ;
      RECT MASK 2 73.721 58.579 73.841 69.791 ;
      RECT MASK 2 74.161 58.579 74.281 69.791 ;
      RECT MASK 2 74.601 58.579 74.721 69.791 ;
      RECT MASK 2 75.041 58.579 75.161 69.791 ;
      RECT MASK 2 75.481 58.579 75.601 69.791 ;
      RECT MASK 2 75.921 58.579 76.041 69.791 ;
      RECT MASK 2 76.361 58.579 76.481 69.791 ;
      RECT MASK 2 76.801 58.579 76.921 69.791 ;
      RECT MASK 2 77.699 58.579 77.819 69.791 ;
      RECT MASK 2 78.139 58.579 78.259 69.791 ;
      RECT MASK 2 78.579 58.579 78.699 69.791 ;
      RECT MASK 2 79.019 58.579 79.139 69.791 ;
      RECT MASK 2 79.459 58.579 79.579 69.791 ;
      RECT MASK 2 79.899 58.579 80.019 69.791 ;
      RECT MASK 2 80.339 58.579 80.459 69.791 ;
      RECT MASK 2 80.779 58.579 80.899 69.791 ;
      RECT MASK 2 81.219 58.579 81.339 69.791 ;
      RECT MASK 2 81.659 58.579 81.779 69.791 ;
      RECT MASK 2 82.099 58.579 82.219 69.791 ;
      RECT MASK 2 82.539 58.579 82.659 69.791 ;
      RECT MASK 2 82.979 58.579 83.099 69.791 ;
      RECT MASK 2 83.419 58.579 83.539 69.791 ;
      RECT MASK 2 84.317 58.579 84.437 69.791 ;
      RECT MASK 2 84.757 58.579 84.877 69.791 ;
      RECT MASK 2 85.197 58.579 85.317 69.791 ;
      RECT MASK 2 85.637 58.579 85.757 69.791 ;
      RECT MASK 2 86.077 58.579 86.197 69.791 ;
      RECT MASK 2 86.517 58.579 86.637 69.791 ;
      RECT MASK 2 86.957 58.579 87.077 69.791 ;
      RECT MASK 2 87.397 58.579 87.517 69.791 ;
      RECT MASK 2 87.837 58.579 87.957 69.791 ;
      RECT MASK 2 88.277 58.579 88.397 69.791 ;
      RECT MASK 2 88.717 58.579 88.837 69.791 ;
      RECT MASK 2 89.157 58.579 89.277 69.791 ;
      RECT MASK 2 89.597 58.579 89.717 69.791 ;
      RECT MASK 2 90.037 58.579 90.157 69.791 ;
      RECT MASK 2 90.935 58.579 91.055 69.791 ;
      RECT MASK 2 91.375 58.579 91.495 69.791 ;
      RECT MASK 2 91.815 58.579 91.935 69.791 ;
      RECT MASK 2 92.255 58.579 92.375 69.791 ;
      RECT MASK 2 92.695 58.579 92.815 69.791 ;
      RECT MASK 2 93.135 58.579 93.255 69.791 ;
      RECT MASK 2 93.575 58.579 93.695 69.791 ;
      RECT MASK 2 94.015 58.579 94.135 69.791 ;
      RECT MASK 2 94.455 58.579 94.575 69.791 ;
      RECT MASK 2 94.895 58.579 95.015 69.791 ;
      RECT MASK 2 95.335 58.579 95.455 69.791 ;
      RECT MASK 2 95.775 58.579 95.895 69.791 ;
      RECT MASK 2 96.215 58.579 96.335 69.791 ;
      RECT MASK 2 96.655 58.579 96.775 69.791 ;
      RECT MASK 2 97.553 58.579 97.673 69.791 ;
      RECT MASK 2 97.993 58.579 98.113 69.791 ;
      RECT MASK 2 98.433 58.579 98.553 69.791 ;
      RECT MASK 2 98.873 58.579 98.993 69.791 ;
      RECT MASK 2 99.313 58.579 99.433 69.791 ;
      RECT MASK 2 99.753 58.579 99.873 69.791 ;
      RECT MASK 2 100.193 58.579 100.313 69.791 ;
      RECT MASK 2 100.633 58.579 100.753 69.791 ;
      RECT MASK 2 101.073 58.579 101.193 69.791 ;
      RECT MASK 2 101.513 58.579 101.633 69.791 ;
      RECT MASK 2 101.953 58.579 102.073 69.791 ;
      RECT MASK 2 102.393 58.579 102.513 69.791 ;
      RECT MASK 2 102.833 58.579 102.953 69.791 ;
      RECT MASK 2 103.273 58.579 103.393 69.791 ;
      RECT MASK 2 104.171 58.579 104.291 69.791 ;
      RECT MASK 2 104.611 58.579 104.731 69.791 ;
      RECT MASK 2 105.051 58.579 105.171 69.791 ;
      RECT MASK 2 105.491 58.579 105.611 69.791 ;
      RECT MASK 2 105.931 58.579 106.051 69.791 ;
      RECT MASK 2 106.371 58.579 106.491 69.791 ;
      RECT MASK 2 106.811 58.579 106.931 69.791 ;
      RECT MASK 2 107.251 58.579 107.371 69.791 ;
      RECT MASK 2 107.691 58.579 107.811 69.791 ;
      RECT MASK 2 108.131 58.579 108.251 69.791 ;
      RECT MASK 2 108.571 58.579 108.691 69.791 ;
      RECT MASK 2 109.011 58.579 109.131 69.791 ;
      RECT MASK 2 109.451 58.579 109.571 69.791 ;
      RECT MASK 2 109.891 58.579 110.011 69.791 ;
      RECT MASK 2 112.5865 59.209 112.7065 60.359 ;
      RECT MASK 2 113.0265 59.209 113.1465 60.359 ;
      RECT MASK 2 113.4665 59.209 113.5865 60.359 ;
      RECT MASK 2 113.9065 59.209 114.0265 60.359 ;
      RECT MASK 2 114.3465 59.209 114.4665 60.359 ;
      RECT MASK 2 114.7865 59.209 114.9065 60.359 ;
      RECT MASK 2 115.2265 59.209 115.3465 60.359 ;
      RECT MASK 2 115.6665 59.209 115.7865 60.359 ;
      RECT MASK 2 116.1065 59.209 116.2265 60.359 ;
      RECT MASK 2 116.5465 59.209 116.6665 60.359 ;
      RECT MASK 2 117.4265 59.209 117.5465 60.359 ;
      RECT MASK 2 117.8665 59.209 117.9865 60.359 ;
      RECT MASK 2 118.3065 59.209 118.4265 60.359 ;
      RECT MASK 2 118.7465 59.209 118.8665 60.359 ;
      RECT MASK 2 119.1865 59.209 119.3065 60.359 ;
      RECT MASK 2 119.6265 59.209 119.7465 60.359 ;
      RECT MASK 2 120.0665 59.209 120.1865 60.359 ;
      RECT MASK 2 120.5065 59.209 120.6265 60.359 ;
      RECT MASK 2 120.9465 59.209 121.0665 60.359 ;
      RECT MASK 2 121.3865 59.209 121.5065 60.359 ;
      RECT MASK 2 121.8265 59.209 121.9465 60.359 ;
      RECT MASK 2 122.2665 59.209 122.3865 60.359 ;
      RECT MASK 2 122.7065 59.209 122.8265 60.359 ;
      RECT MASK 2 123.1465 59.209 123.2665 60.359 ;
      RECT MASK 2 123.5865 59.209 123.7065 60.359 ;
      RECT MASK 2 112.5865 60.619 112.7065 61.649 ;
      RECT MASK 2 113.0265 60.619 113.1465 61.649 ;
      RECT MASK 2 113.4665 60.619 113.5865 61.649 ;
      RECT MASK 2 113.9065 60.619 114.0265 61.649 ;
      RECT MASK 2 114.3465 60.619 114.4665 61.649 ;
      RECT MASK 2 114.7865 60.619 114.9065 61.649 ;
      RECT MASK 2 115.2265 60.619 115.3465 61.649 ;
      RECT MASK 2 115.6665 60.619 115.7865 61.649 ;
      RECT MASK 2 116.1065 60.619 116.2265 61.649 ;
      RECT MASK 2 116.5465 60.619 116.6665 61.649 ;
      RECT MASK 2 117.4265 60.619 117.5465 61.649 ;
      RECT MASK 2 117.8665 60.619 117.9865 61.649 ;
      RECT MASK 2 118.3065 60.619 118.4265 61.649 ;
      RECT MASK 2 118.7465 60.619 118.8665 61.649 ;
      RECT MASK 2 119.1865 60.619 119.3065 61.649 ;
      RECT MASK 2 119.6265 60.619 119.7465 61.649 ;
      RECT MASK 2 120.0665 60.619 120.1865 61.649 ;
      RECT MASK 2 120.5065 60.619 120.6265 61.649 ;
      RECT MASK 2 120.9465 60.619 121.0665 61.649 ;
      RECT MASK 2 121.3865 60.619 121.5065 61.649 ;
      RECT MASK 2 121.8265 60.619 121.9465 61.649 ;
      RECT MASK 2 122.2665 60.619 122.3865 61.649 ;
      RECT MASK 2 122.7065 60.619 122.8265 61.649 ;
      RECT MASK 2 123.1465 60.619 123.2665 61.649 ;
      RECT MASK 2 123.5865 60.619 123.7065 61.649 ;
      RECT MASK 2 112.5865 61.909 112.7065 62.999 ;
      RECT MASK 2 113.0265 61.909 113.1465 62.999 ;
      RECT MASK 2 113.4665 61.909 113.5865 62.999 ;
      RECT MASK 2 113.9065 61.909 114.0265 62.999 ;
      RECT MASK 2 114.3465 61.909 114.4665 62.999 ;
      RECT MASK 2 114.7865 61.909 114.9065 62.999 ;
      RECT MASK 2 115.2265 61.909 115.3465 62.999 ;
      RECT MASK 2 115.6665 61.909 115.7865 62.999 ;
      RECT MASK 2 116.1065 61.909 116.2265 62.999 ;
      RECT MASK 2 116.5465 61.909 116.6665 62.999 ;
      RECT MASK 2 117.4265 61.909 117.5465 62.999 ;
      RECT MASK 2 117.8665 61.909 117.9865 62.999 ;
      RECT MASK 2 118.3065 61.909 118.4265 62.999 ;
      RECT MASK 2 118.7465 61.909 118.8665 62.999 ;
      RECT MASK 2 119.1865 61.909 119.3065 62.999 ;
      RECT MASK 2 119.6265 61.909 119.7465 62.999 ;
      RECT MASK 2 120.0665 61.909 120.1865 62.999 ;
      RECT MASK 2 120.5065 61.909 120.6265 62.999 ;
      RECT MASK 2 120.9465 61.909 121.0665 62.999 ;
      RECT MASK 2 121.3865 61.909 121.5065 62.999 ;
      RECT MASK 2 121.8265 61.909 121.9465 62.999 ;
      RECT MASK 2 122.2665 61.909 122.3865 62.999 ;
      RECT MASK 2 122.7065 61.909 122.8265 62.999 ;
      RECT MASK 2 123.1465 61.909 123.2665 62.999 ;
      RECT MASK 2 123.5865 61.909 123.7065 62.999 ;
      RECT MASK 2 112.5865 63.259 112.7065 65.069 ;
      RECT MASK 2 113.0265 63.259 113.1465 65.069 ;
      RECT MASK 2 113.4665 63.259 113.5865 65.069 ;
      RECT MASK 2 113.9065 63.259 114.0265 65.069 ;
      RECT MASK 2 114.3465 63.259 114.4665 65.069 ;
      RECT MASK 2 114.7865 63.259 114.9065 65.069 ;
      RECT MASK 2 115.2265 63.259 115.3465 65.069 ;
      RECT MASK 2 115.6665 63.259 115.7865 65.069 ;
      RECT MASK 2 116.1065 63.259 116.2265 65.069 ;
      RECT MASK 2 116.5465 63.259 116.6665 65.069 ;
      RECT MASK 2 117.4265 63.259 117.5465 65.069 ;
      RECT MASK 2 117.8665 63.259 117.9865 65.069 ;
      RECT MASK 2 118.3065 63.259 118.4265 65.069 ;
      RECT MASK 2 118.7465 63.259 118.8665 65.069 ;
      RECT MASK 2 119.1865 63.259 119.3065 65.069 ;
      RECT MASK 2 119.6265 63.259 119.7465 65.069 ;
      RECT MASK 2 120.0665 63.259 120.1865 65.069 ;
      RECT MASK 2 120.5065 63.259 120.6265 65.069 ;
      RECT MASK 2 120.9465 63.259 121.0665 65.069 ;
      RECT MASK 2 121.3865 63.259 121.5065 65.069 ;
      RECT MASK 2 121.8265 63.259 121.9465 65.069 ;
      RECT MASK 2 122.2665 63.259 122.3865 65.069 ;
      RECT MASK 2 122.7065 63.259 122.8265 65.069 ;
      RECT MASK 2 123.1465 63.259 123.2665 65.069 ;
      RECT MASK 2 123.5865 63.259 123.7065 65.069 ;
      RECT MASK 2 112.5865 65.329 112.7065 66.419 ;
      RECT MASK 2 113.0265 65.329 113.1465 66.419 ;
      RECT MASK 2 113.4665 65.329 113.5865 66.419 ;
      RECT MASK 2 113.9065 65.329 114.0265 66.419 ;
      RECT MASK 2 114.3465 65.329 114.4665 66.419 ;
      RECT MASK 2 114.7865 65.329 114.9065 66.419 ;
      RECT MASK 2 115.2265 65.329 115.3465 66.419 ;
      RECT MASK 2 115.6665 65.329 115.7865 66.419 ;
      RECT MASK 2 116.1065 65.329 116.2265 66.419 ;
      RECT MASK 2 116.5465 65.329 116.6665 66.419 ;
      RECT MASK 2 117.4265 65.329 117.5465 66.419 ;
      RECT MASK 2 117.8665 65.329 117.9865 66.419 ;
      RECT MASK 2 118.3065 65.329 118.4265 66.419 ;
      RECT MASK 2 118.7465 65.329 118.8665 66.419 ;
      RECT MASK 2 119.1865 65.329 119.3065 66.419 ;
      RECT MASK 2 119.6265 65.329 119.7465 66.419 ;
      RECT MASK 2 120.0665 65.329 120.1865 66.419 ;
      RECT MASK 2 120.5065 65.329 120.6265 66.419 ;
      RECT MASK 2 120.9465 65.329 121.0665 66.419 ;
      RECT MASK 2 121.3865 65.329 121.5065 66.419 ;
      RECT MASK 2 121.8265 65.329 121.9465 66.419 ;
      RECT MASK 2 122.2665 65.329 122.3865 66.419 ;
      RECT MASK 2 122.7065 65.329 122.8265 66.419 ;
      RECT MASK 2 123.1465 65.329 123.2665 66.419 ;
      RECT MASK 2 123.5865 65.329 123.7065 66.419 ;
      RECT MASK 2 112.5865 66.679 112.7065 67.769 ;
      RECT MASK 2 113.0265 66.679 113.1465 67.769 ;
      RECT MASK 2 113.4665 66.679 113.5865 67.769 ;
      RECT MASK 2 113.9065 66.679 114.0265 67.769 ;
      RECT MASK 2 114.3465 66.679 114.4665 67.769 ;
      RECT MASK 2 114.7865 66.679 114.9065 67.769 ;
      RECT MASK 2 115.2265 66.679 115.3465 67.769 ;
      RECT MASK 2 115.6665 66.679 115.7865 67.769 ;
      RECT MASK 2 116.1065 66.679 116.2265 67.769 ;
      RECT MASK 2 116.5465 66.679 116.6665 67.769 ;
      RECT MASK 2 117.4265 66.679 117.5465 67.769 ;
      RECT MASK 2 117.8665 66.679 117.9865 67.769 ;
      RECT MASK 2 118.3065 66.679 118.4265 67.769 ;
      RECT MASK 2 118.7465 66.679 118.8665 67.769 ;
      RECT MASK 2 119.1865 66.679 119.3065 67.769 ;
      RECT MASK 2 119.6265 66.679 119.7465 67.769 ;
      RECT MASK 2 120.0665 66.679 120.1865 67.769 ;
      RECT MASK 2 120.5065 66.679 120.6265 67.769 ;
      RECT MASK 2 120.9465 66.679 121.0665 67.769 ;
      RECT MASK 2 121.3865 66.679 121.5065 67.769 ;
      RECT MASK 2 121.8265 66.679 121.9465 67.769 ;
      RECT MASK 2 122.2665 66.679 122.3865 67.769 ;
      RECT MASK 2 122.7065 66.679 122.8265 67.769 ;
      RECT MASK 2 123.1465 66.679 123.2665 67.769 ;
      RECT MASK 2 123.5865 66.679 123.7065 67.769 ;
      RECT MASK 2 112.5865 68.029 112.7065 69.119 ;
      RECT MASK 2 113.0265 68.029 113.1465 69.119 ;
      RECT MASK 2 113.4665 68.029 113.5865 69.119 ;
      RECT MASK 2 113.9065 68.029 114.0265 69.119 ;
      RECT MASK 2 114.3465 68.029 114.4665 69.119 ;
      RECT MASK 2 114.7865 68.029 114.9065 69.119 ;
      RECT MASK 2 115.2265 68.029 115.3465 69.119 ;
      RECT MASK 2 115.6665 68.029 115.7865 69.119 ;
      RECT MASK 2 116.1065 68.029 116.2265 69.119 ;
      RECT MASK 2 116.5465 68.029 116.6665 69.119 ;
      RECT MASK 2 117.4265 68.029 117.5465 69.119 ;
      RECT MASK 2 117.8665 68.029 117.9865 69.119 ;
      RECT MASK 2 118.3065 68.029 118.4265 69.119 ;
      RECT MASK 2 118.7465 68.029 118.8665 69.119 ;
      RECT MASK 2 119.1865 68.029 119.3065 69.119 ;
      RECT MASK 2 119.6265 68.029 119.7465 69.119 ;
      RECT MASK 2 120.0665 68.029 120.1865 69.119 ;
      RECT MASK 2 120.5065 68.029 120.6265 69.119 ;
      RECT MASK 2 120.9465 68.029 121.0665 69.119 ;
      RECT MASK 2 121.3865 68.029 121.5065 69.119 ;
      RECT MASK 2 121.8265 68.029 121.9465 69.119 ;
      RECT MASK 2 122.2665 68.029 122.3865 69.119 ;
      RECT MASK 2 122.7065 68.029 122.8265 69.119 ;
      RECT MASK 2 123.1465 68.029 123.2665 69.119 ;
      RECT MASK 2 123.5865 68.029 123.7065 69.119 ;
      RECT MASK 2 112.5865 69.379 112.7065 71.189 ;
      RECT MASK 2 113.0265 69.379 113.1465 71.189 ;
      RECT MASK 2 113.4665 69.379 113.5865 71.189 ;
      RECT MASK 2 113.9065 69.379 114.0265 71.189 ;
      RECT MASK 2 114.3465 69.379 114.4665 71.189 ;
      RECT MASK 2 114.7865 69.379 114.9065 71.189 ;
      RECT MASK 2 115.2265 69.379 115.3465 71.189 ;
      RECT MASK 2 115.6665 69.379 115.7865 71.189 ;
      RECT MASK 2 116.1065 69.379 116.2265 71.189 ;
      RECT MASK 2 116.5465 69.379 116.6665 71.189 ;
      RECT MASK 2 117.4265 69.379 117.5465 71.189 ;
      RECT MASK 2 117.8665 69.379 117.9865 71.189 ;
      RECT MASK 2 118.3065 69.379 118.4265 71.189 ;
      RECT MASK 2 118.7465 69.379 118.8665 71.189 ;
      RECT MASK 2 119.1865 69.379 119.3065 71.189 ;
      RECT MASK 2 119.6265 69.379 119.7465 71.189 ;
      RECT MASK 2 120.0665 69.379 120.1865 71.189 ;
      RECT MASK 2 120.5065 69.379 120.6265 71.189 ;
      RECT MASK 2 120.9465 69.379 121.0665 71.189 ;
      RECT MASK 2 121.3865 69.379 121.5065 71.189 ;
      RECT MASK 2 121.8265 69.379 121.9465 71.189 ;
      RECT MASK 2 122.2665 69.379 122.3865 71.189 ;
      RECT MASK 2 122.7065 69.379 122.8265 71.189 ;
      RECT MASK 2 123.1465 69.379 123.2665 71.189 ;
      RECT MASK 2 123.5865 69.379 123.7065 71.189 ;
      RECT MASK 2 4.931 69.96 4.991 70.2 ;
      RECT MASK 2 5.371 69.96 5.431 70.2 ;
      RECT MASK 2 5.811 69.96 5.871 70.2 ;
      RECT MASK 2 6.251 69.96 6.311 70.2 ;
      RECT MASK 2 6.691 69.96 6.751 70.2 ;
      RECT MASK 2 7.131 69.96 7.191 70.2 ;
      RECT MASK 2 7.571 69.96 7.631 70.2 ;
      RECT MASK 2 8.011 69.96 8.071 70.2 ;
      RECT MASK 2 8.451 69.96 8.511 70.2 ;
      RECT MASK 2 8.891 69.96 8.951 70.2 ;
      RECT MASK 2 9.331 69.96 9.391 70.2 ;
      RECT MASK 2 9.771 69.96 9.831 70.2 ;
      RECT MASK 2 10.211 69.96 10.271 70.2 ;
      RECT MASK 2 10.651 69.96 10.711 70.2 ;
      RECT MASK 2 11.549 69.96 11.609 70.2 ;
      RECT MASK 2 11.989 69.96 12.049 70.2 ;
      RECT MASK 2 12.429 69.96 12.489 70.2 ;
      RECT MASK 2 12.869 69.96 12.929 70.2 ;
      RECT MASK 2 13.309 69.96 13.369 70.2 ;
      RECT MASK 2 13.749 69.96 13.809 70.2 ;
      RECT MASK 2 14.189 69.96 14.249 70.2 ;
      RECT MASK 2 14.629 69.96 14.689 70.2 ;
      RECT MASK 2 15.069 69.96 15.129 70.2 ;
      RECT MASK 2 15.509 69.96 15.569 70.2 ;
      RECT MASK 2 15.949 69.96 16.009 70.2 ;
      RECT MASK 2 16.389 69.96 16.449 70.2 ;
      RECT MASK 2 16.829 69.96 16.889 70.2 ;
      RECT MASK 2 17.269 69.96 17.329 70.2 ;
      RECT MASK 2 18.167 69.96 18.227 70.2 ;
      RECT MASK 2 18.607 69.96 18.667 70.2 ;
      RECT MASK 2 19.047 69.96 19.107 70.2 ;
      RECT MASK 2 19.487 69.96 19.547 70.2 ;
      RECT MASK 2 19.927 69.96 19.987 70.2 ;
      RECT MASK 2 20.367 69.96 20.427 70.2 ;
      RECT MASK 2 20.807 69.96 20.867 70.2 ;
      RECT MASK 2 21.247 69.96 21.307 70.2 ;
      RECT MASK 2 21.687 69.96 21.747 70.2 ;
      RECT MASK 2 22.127 69.96 22.187 70.2 ;
      RECT MASK 2 22.567 69.96 22.627 70.2 ;
      RECT MASK 2 23.007 69.96 23.067 70.2 ;
      RECT MASK 2 23.447 69.96 23.507 70.2 ;
      RECT MASK 2 23.887 69.96 23.947 70.2 ;
      RECT MASK 2 24.785 69.96 24.845 70.2 ;
      RECT MASK 2 25.225 69.96 25.285 70.2 ;
      RECT MASK 2 25.665 69.96 25.725 70.2 ;
      RECT MASK 2 26.105 69.96 26.165 70.2 ;
      RECT MASK 2 26.545 69.96 26.605 70.2 ;
      RECT MASK 2 26.985 69.96 27.045 70.2 ;
      RECT MASK 2 27.425 69.96 27.485 70.2 ;
      RECT MASK 2 27.865 69.96 27.925 70.2 ;
      RECT MASK 2 28.305 69.96 28.365 70.2 ;
      RECT MASK 2 28.745 69.96 28.805 70.2 ;
      RECT MASK 2 29.185 69.96 29.245 70.2 ;
      RECT MASK 2 29.625 69.96 29.685 70.2 ;
      RECT MASK 2 30.065 69.96 30.125 70.2 ;
      RECT MASK 2 30.505 69.96 30.565 70.2 ;
      RECT MASK 2 31.403 69.96 31.463 70.2 ;
      RECT MASK 2 31.843 69.96 31.903 70.2 ;
      RECT MASK 2 32.283 69.96 32.343 70.2 ;
      RECT MASK 2 32.723 69.96 32.783 70.2 ;
      RECT MASK 2 33.163 69.96 33.223 70.2 ;
      RECT MASK 2 33.603 69.96 33.663 70.2 ;
      RECT MASK 2 34.043 69.96 34.103 70.2 ;
      RECT MASK 2 34.483 69.96 34.543 70.2 ;
      RECT MASK 2 34.923 69.96 34.983 70.2 ;
      RECT MASK 2 35.363 69.96 35.423 70.2 ;
      RECT MASK 2 35.803 69.96 35.863 70.2 ;
      RECT MASK 2 36.243 69.96 36.303 70.2 ;
      RECT MASK 2 36.683 69.96 36.743 70.2 ;
      RECT MASK 2 37.123 69.96 37.183 70.2 ;
      RECT MASK 2 38.021 69.96 38.081 70.2 ;
      RECT MASK 2 38.461 69.96 38.521 70.2 ;
      RECT MASK 2 38.901 69.96 38.961 70.2 ;
      RECT MASK 2 39.341 69.96 39.401 70.2 ;
      RECT MASK 2 39.781 69.96 39.841 70.2 ;
      RECT MASK 2 40.221 69.96 40.281 70.2 ;
      RECT MASK 2 40.661 69.96 40.721 70.2 ;
      RECT MASK 2 41.101 69.96 41.161 70.2 ;
      RECT MASK 2 41.541 69.96 41.601 70.2 ;
      RECT MASK 2 42.861 69.96 42.921 70.2 ;
      RECT MASK 2 43.301 69.96 43.361 70.2 ;
      RECT MASK 2 43.741 69.96 43.801 70.2 ;
      RECT MASK 2 44.639 69.96 44.699 70.2 ;
      RECT MASK 2 45.079 69.96 45.139 70.2 ;
      RECT MASK 2 45.519 69.96 45.579 70.2 ;
      RECT MASK 2 45.959 69.96 46.019 70.2 ;
      RECT MASK 2 46.399 69.96 46.459 70.2 ;
      RECT MASK 2 46.839 69.96 46.899 70.2 ;
      RECT MASK 2 47.279 69.96 47.339 70.2 ;
      RECT MASK 2 47.719 69.96 47.779 70.2 ;
      RECT MASK 2 48.159 69.96 48.219 70.2 ;
      RECT MASK 2 48.599 69.96 48.659 70.2 ;
      RECT MASK 2 49.039 69.96 49.099 70.2 ;
      RECT MASK 2 49.479 69.96 49.539 70.2 ;
      RECT MASK 2 49.919 69.96 49.979 70.2 ;
      RECT MASK 2 50.359 69.96 50.419 70.2 ;
      RECT MASK 2 51.257 69.96 51.317 70.2 ;
      RECT MASK 2 51.697 69.96 51.757 70.2 ;
      RECT MASK 2 52.137 69.96 52.197 70.2 ;
      RECT MASK 2 52.577 69.96 52.637 70.2 ;
      RECT MASK 2 53.017 69.96 53.077 70.2 ;
      RECT MASK 2 53.457 69.96 53.517 70.2 ;
      RECT MASK 2 53.897 69.96 53.957 70.2 ;
      RECT MASK 2 54.337 69.96 54.397 70.2 ;
      RECT MASK 2 54.777 69.96 54.837 70.2 ;
      RECT MASK 2 55.217 69.96 55.277 70.2 ;
      RECT MASK 2 55.657 69.96 55.717 70.2 ;
      RECT MASK 2 56.097 69.96 56.157 70.2 ;
      RECT MASK 2 56.537 69.96 56.597 70.2 ;
      RECT MASK 2 56.977 69.96 57.037 70.2 ;
      RECT MASK 2 57.875 69.96 57.935 70.2 ;
      RECT MASK 2 58.315 69.96 58.375 70.2 ;
      RECT MASK 2 58.755 69.96 58.815 70.2 ;
      RECT MASK 2 59.195 69.96 59.255 70.2 ;
      RECT MASK 2 59.635 69.96 59.695 70.2 ;
      RECT MASK 2 60.075 69.96 60.135 70.2 ;
      RECT MASK 2 60.515 69.96 60.575 70.2 ;
      RECT MASK 2 60.955 69.96 61.015 70.2 ;
      RECT MASK 2 61.395 69.96 61.455 70.2 ;
      RECT MASK 2 61.835 69.96 61.895 70.2 ;
      RECT MASK 2 62.275 69.96 62.335 70.2 ;
      RECT MASK 2 62.715 69.96 62.775 70.2 ;
      RECT MASK 2 63.155 69.96 63.215 70.2 ;
      RECT MASK 2 63.595 69.96 63.655 70.2 ;
      RECT MASK 2 64.493 69.96 64.553 70.2 ;
      RECT MASK 2 64.933 69.96 64.993 70.2 ;
      RECT MASK 2 65.373 69.96 65.433 70.2 ;
      RECT MASK 2 65.813 69.96 65.873 70.2 ;
      RECT MASK 2 66.253 69.96 66.313 70.2 ;
      RECT MASK 2 66.693 69.96 66.753 70.2 ;
      RECT MASK 2 67.133 69.96 67.193 70.2 ;
      RECT MASK 2 67.573 69.96 67.633 70.2 ;
      RECT MASK 2 68.013 69.96 68.073 70.2 ;
      RECT MASK 2 68.453 69.96 68.513 70.2 ;
      RECT MASK 2 68.893 69.96 68.953 70.2 ;
      RECT MASK 2 69.333 69.96 69.393 70.2 ;
      RECT MASK 2 69.773 69.96 69.833 70.2 ;
      RECT MASK 2 70.213 69.96 70.273 70.2 ;
      RECT MASK 2 71.111 69.96 71.171 70.2 ;
      RECT MASK 2 71.551 69.96 71.611 70.2 ;
      RECT MASK 2 71.991 69.96 72.051 70.2 ;
      RECT MASK 2 72.431 69.96 72.491 70.2 ;
      RECT MASK 2 72.871 69.96 72.931 70.2 ;
      RECT MASK 2 73.311 69.96 73.371 70.2 ;
      RECT MASK 2 73.751 69.96 73.811 70.2 ;
      RECT MASK 2 74.191 69.96 74.251 70.2 ;
      RECT MASK 2 74.631 69.96 74.691 70.2 ;
      RECT MASK 2 75.071 69.96 75.131 70.2 ;
      RECT MASK 2 75.511 69.96 75.571 70.2 ;
      RECT MASK 2 75.951 69.96 76.011 70.2 ;
      RECT MASK 2 76.391 69.96 76.451 70.2 ;
      RECT MASK 2 76.831 69.96 76.891 70.2 ;
      RECT MASK 2 77.729 69.96 77.789 70.2 ;
      RECT MASK 2 78.169 69.96 78.229 70.2 ;
      RECT MASK 2 78.609 69.96 78.669 70.2 ;
      RECT MASK 2 79.049 69.96 79.109 70.2 ;
      RECT MASK 2 79.489 69.96 79.549 70.2 ;
      RECT MASK 2 79.929 69.96 79.989 70.2 ;
      RECT MASK 2 80.369 69.96 80.429 70.2 ;
      RECT MASK 2 80.809 69.96 80.869 70.2 ;
      RECT MASK 2 81.249 69.96 81.309 70.2 ;
      RECT MASK 2 81.689 69.96 81.749 70.2 ;
      RECT MASK 2 82.129 69.96 82.189 70.2 ;
      RECT MASK 2 83.449 69.96 83.509 70.2 ;
      RECT MASK 2 84.347 69.96 84.407 70.2 ;
      RECT MASK 2 84.787 69.96 84.847 70.2 ;
      RECT MASK 2 85.227 69.96 85.287 70.2 ;
      RECT MASK 2 85.667 69.96 85.727 70.2 ;
      RECT MASK 2 86.107 69.96 86.167 70.2 ;
      RECT MASK 2 86.547 69.96 86.607 70.2 ;
      RECT MASK 2 86.987 69.96 87.047 70.2 ;
      RECT MASK 2 87.427 69.96 87.487 70.2 ;
      RECT MASK 2 87.867 69.96 87.927 70.2 ;
      RECT MASK 2 88.307 69.96 88.367 70.2 ;
      RECT MASK 2 88.747 69.96 88.807 70.2 ;
      RECT MASK 2 89.187 69.96 89.247 70.2 ;
      RECT MASK 2 89.627 69.96 89.687 70.2 ;
      RECT MASK 2 90.067 69.96 90.127 70.2 ;
      RECT MASK 2 90.965 69.96 91.025 70.2 ;
      RECT MASK 2 91.405 69.96 91.465 70.2 ;
      RECT MASK 2 91.845 69.96 91.905 70.2 ;
      RECT MASK 2 92.285 69.96 92.345 70.2 ;
      RECT MASK 2 92.725 69.96 92.785 70.2 ;
      RECT MASK 2 93.165 69.96 93.225 70.2 ;
      RECT MASK 2 93.605 69.96 93.665 70.2 ;
      RECT MASK 2 94.045 69.96 94.105 70.2 ;
      RECT MASK 2 94.485 69.96 94.545 70.2 ;
      RECT MASK 2 94.925 69.96 94.985 70.2 ;
      RECT MASK 2 95.365 69.96 95.425 70.2 ;
      RECT MASK 2 95.805 69.96 95.865 70.2 ;
      RECT MASK 2 96.245 69.96 96.305 70.2 ;
      RECT MASK 2 96.685 69.96 96.745 70.2 ;
      RECT MASK 2 97.583 69.96 97.643 70.2 ;
      RECT MASK 2 98.023 69.96 98.083 70.2 ;
      RECT MASK 2 98.463 69.96 98.523 70.2 ;
      RECT MASK 2 98.903 69.96 98.963 70.2 ;
      RECT MASK 2 99.343 69.96 99.403 70.2 ;
      RECT MASK 2 99.783 69.96 99.843 70.2 ;
      RECT MASK 2 100.223 69.96 100.283 70.2 ;
      RECT MASK 2 100.663 69.96 100.723 70.2 ;
      RECT MASK 2 101.103 69.96 101.163 70.2 ;
      RECT MASK 2 101.543 69.96 101.603 70.2 ;
      RECT MASK 2 101.983 69.96 102.043 70.2 ;
      RECT MASK 2 102.423 69.96 102.483 70.2 ;
      RECT MASK 2 102.863 69.96 102.923 70.2 ;
      RECT MASK 2 103.303 69.96 103.363 70.2 ;
      RECT MASK 2 104.201 69.96 104.261 70.2 ;
      RECT MASK 2 104.641 69.96 104.701 70.2 ;
      RECT MASK 2 105.081 69.96 105.141 70.2 ;
      RECT MASK 2 105.521 69.96 105.581 70.2 ;
      RECT MASK 2 105.961 69.96 106.021 70.2 ;
      RECT MASK 2 106.401 69.96 106.461 70.2 ;
      RECT MASK 2 106.841 69.96 106.901 70.2 ;
      RECT MASK 2 107.281 69.96 107.341 70.2 ;
      RECT MASK 2 107.721 69.96 107.781 70.2 ;
      RECT MASK 2 108.161 69.96 108.221 70.2 ;
      RECT MASK 2 108.601 69.96 108.661 70.2 ;
      RECT MASK 2 109.041 69.96 109.101 70.2 ;
      RECT MASK 2 109.481 69.96 109.541 70.2 ;
      RECT MASK 2 109.921 69.96 109.981 70.2 ;
      RECT MASK 2 4.931 70.38 4.991 70.62 ;
      RECT MASK 2 5.371 70.38 5.431 70.62 ;
      RECT MASK 2 5.811 70.38 5.871 70.62 ;
      RECT MASK 2 6.251 70.38 6.311 70.62 ;
      RECT MASK 2 6.691 70.38 6.751 70.62 ;
      RECT MASK 2 7.131 70.38 7.191 70.62 ;
      RECT MASK 2 7.571 70.38 7.631 70.62 ;
      RECT MASK 2 8.011 70.38 8.071 70.62 ;
      RECT MASK 2 8.451 70.38 8.511 70.62 ;
      RECT MASK 2 8.891 70.38 8.951 70.62 ;
      RECT MASK 2 9.331 70.38 9.391 70.62 ;
      RECT MASK 2 9.771 70.38 9.831 70.62 ;
      RECT MASK 2 10.211 70.38 10.271 70.62 ;
      RECT MASK 2 10.651 70.38 10.711 70.62 ;
      RECT MASK 2 11.549 70.38 11.609 70.62 ;
      RECT MASK 2 11.989 70.38 12.049 70.62 ;
      RECT MASK 2 12.429 70.38 12.489 70.62 ;
      RECT MASK 2 12.869 70.38 12.929 70.62 ;
      RECT MASK 2 13.309 70.38 13.369 70.62 ;
      RECT MASK 2 13.749 70.38 13.809 70.62 ;
      RECT MASK 2 14.189 70.38 14.249 70.62 ;
      RECT MASK 2 14.629 70.38 14.689 70.62 ;
      RECT MASK 2 15.069 70.38 15.129 70.62 ;
      RECT MASK 2 15.509 70.38 15.569 70.62 ;
      RECT MASK 2 15.949 70.38 16.009 70.62 ;
      RECT MASK 2 16.389 70.38 16.449 70.62 ;
      RECT MASK 2 16.829 70.38 16.889 70.62 ;
      RECT MASK 2 17.269 70.38 17.329 70.62 ;
      RECT MASK 2 18.167 70.38 18.227 70.62 ;
      RECT MASK 2 18.607 70.38 18.667 70.62 ;
      RECT MASK 2 19.047 70.38 19.107 70.62 ;
      RECT MASK 2 19.487 70.38 19.547 70.62 ;
      RECT MASK 2 19.927 70.38 19.987 70.62 ;
      RECT MASK 2 20.367 70.38 20.427 70.62 ;
      RECT MASK 2 20.807 70.38 20.867 70.62 ;
      RECT MASK 2 21.247 70.38 21.307 70.62 ;
      RECT MASK 2 21.687 70.38 21.747 70.62 ;
      RECT MASK 2 22.127 70.38 22.187 70.62 ;
      RECT MASK 2 22.567 70.38 22.627 70.62 ;
      RECT MASK 2 23.007 70.38 23.067 70.62 ;
      RECT MASK 2 23.447 70.38 23.507 70.62 ;
      RECT MASK 2 23.887 70.38 23.947 70.62 ;
      RECT MASK 2 24.785 70.38 24.845 70.62 ;
      RECT MASK 2 25.225 70.38 25.285 70.62 ;
      RECT MASK 2 25.665 70.38 25.725 70.62 ;
      RECT MASK 2 26.105 70.38 26.165 70.62 ;
      RECT MASK 2 26.545 70.38 26.605 70.62 ;
      RECT MASK 2 26.985 70.38 27.045 70.62 ;
      RECT MASK 2 27.425 70.38 27.485 70.62 ;
      RECT MASK 2 27.865 70.38 27.925 70.62 ;
      RECT MASK 2 28.305 70.38 28.365 70.62 ;
      RECT MASK 2 28.745 70.38 28.805 70.62 ;
      RECT MASK 2 29.185 70.38 29.245 70.62 ;
      RECT MASK 2 29.625 70.38 29.685 70.62 ;
      RECT MASK 2 30.065 70.38 30.125 70.62 ;
      RECT MASK 2 30.505 70.38 30.565 70.62 ;
      RECT MASK 2 31.403 70.38 31.463 70.62 ;
      RECT MASK 2 31.843 70.38 31.903 70.62 ;
      RECT MASK 2 32.283 70.38 32.343 70.62 ;
      RECT MASK 2 32.723 70.38 32.783 70.62 ;
      RECT MASK 2 33.163 70.38 33.223 70.62 ;
      RECT MASK 2 33.603 70.38 33.663 70.62 ;
      RECT MASK 2 34.043 70.38 34.103 70.62 ;
      RECT MASK 2 34.483 70.38 34.543 70.62 ;
      RECT MASK 2 34.923 70.38 34.983 70.62 ;
      RECT MASK 2 35.363 70.38 35.423 70.62 ;
      RECT MASK 2 35.803 70.38 35.863 70.62 ;
      RECT MASK 2 36.243 70.38 36.303 70.62 ;
      RECT MASK 2 36.683 70.38 36.743 70.62 ;
      RECT MASK 2 37.123 70.38 37.183 70.62 ;
      RECT MASK 2 38.021 70.38 38.081 70.62 ;
      RECT MASK 2 38.461 70.38 38.521 70.62 ;
      RECT MASK 2 38.901 70.38 38.961 70.62 ;
      RECT MASK 2 39.341 70.38 39.401 70.62 ;
      RECT MASK 2 39.781 70.38 39.841 70.62 ;
      RECT MASK 2 40.221 70.38 40.281 70.62 ;
      RECT MASK 2 40.661 70.38 40.721 70.62 ;
      RECT MASK 2 41.101 70.38 41.161 70.62 ;
      RECT MASK 2 41.541 70.38 41.601 70.62 ;
      RECT MASK 2 42.861 70.38 42.921 70.62 ;
      RECT MASK 2 43.301 70.38 43.361 70.62 ;
      RECT MASK 2 43.741 70.38 43.801 70.62 ;
      RECT MASK 2 44.639 70.38 44.699 70.62 ;
      RECT MASK 2 45.079 70.38 45.139 70.62 ;
      RECT MASK 2 45.519 70.38 45.579 70.62 ;
      RECT MASK 2 45.959 70.38 46.019 70.62 ;
      RECT MASK 2 46.399 70.38 46.459 70.62 ;
      RECT MASK 2 46.839 70.38 46.899 70.62 ;
      RECT MASK 2 47.279 70.38 47.339 70.62 ;
      RECT MASK 2 47.719 70.38 47.779 70.62 ;
      RECT MASK 2 48.159 70.38 48.219 70.62 ;
      RECT MASK 2 48.599 70.38 48.659 70.62 ;
      RECT MASK 2 49.039 70.38 49.099 70.62 ;
      RECT MASK 2 49.479 70.38 49.539 70.62 ;
      RECT MASK 2 49.919 70.38 49.979 70.62 ;
      RECT MASK 2 50.359 70.38 50.419 70.62 ;
      RECT MASK 2 51.257 70.38 51.317 70.62 ;
      RECT MASK 2 51.697 70.38 51.757 70.62 ;
      RECT MASK 2 52.137 70.38 52.197 70.62 ;
      RECT MASK 2 52.577 70.38 52.637 70.62 ;
      RECT MASK 2 53.017 70.38 53.077 70.62 ;
      RECT MASK 2 53.457 70.38 53.517 70.62 ;
      RECT MASK 2 53.897 70.38 53.957 70.62 ;
      RECT MASK 2 54.337 70.38 54.397 70.62 ;
      RECT MASK 2 54.777 70.38 54.837 70.62 ;
      RECT MASK 2 55.217 70.38 55.277 70.62 ;
      RECT MASK 2 55.657 70.38 55.717 70.62 ;
      RECT MASK 2 56.097 70.38 56.157 70.62 ;
      RECT MASK 2 56.537 70.38 56.597 70.62 ;
      RECT MASK 2 56.977 70.38 57.037 70.62 ;
      RECT MASK 2 57.875 70.38 57.935 70.62 ;
      RECT MASK 2 58.315 70.38 58.375 70.62 ;
      RECT MASK 2 58.755 70.38 58.815 70.62 ;
      RECT MASK 2 59.195 70.38 59.255 70.62 ;
      RECT MASK 2 59.635 70.38 59.695 70.62 ;
      RECT MASK 2 60.075 70.38 60.135 70.62 ;
      RECT MASK 2 60.515 70.38 60.575 70.62 ;
      RECT MASK 2 60.955 70.38 61.015 70.62 ;
      RECT MASK 2 61.395 70.38 61.455 70.62 ;
      RECT MASK 2 61.835 70.38 61.895 70.62 ;
      RECT MASK 2 62.275 70.38 62.335 70.62 ;
      RECT MASK 2 62.715 70.38 62.775 70.62 ;
      RECT MASK 2 63.155 70.38 63.215 70.62 ;
      RECT MASK 2 63.595 70.38 63.655 70.62 ;
      RECT MASK 2 64.493 70.38 64.553 70.62 ;
      RECT MASK 2 64.933 70.38 64.993 70.62 ;
      RECT MASK 2 65.373 70.38 65.433 70.62 ;
      RECT MASK 2 65.813 70.38 65.873 70.62 ;
      RECT MASK 2 66.253 70.38 66.313 70.62 ;
      RECT MASK 2 66.693 70.38 66.753 70.62 ;
      RECT MASK 2 67.133 70.38 67.193 70.62 ;
      RECT MASK 2 67.573 70.38 67.633 70.62 ;
      RECT MASK 2 68.013 70.38 68.073 70.62 ;
      RECT MASK 2 68.453 70.38 68.513 70.62 ;
      RECT MASK 2 68.893 70.38 68.953 70.62 ;
      RECT MASK 2 69.333 70.38 69.393 70.62 ;
      RECT MASK 2 69.773 70.38 69.833 70.62 ;
      RECT MASK 2 70.213 70.38 70.273 70.62 ;
      RECT MASK 2 71.111 70.38 71.171 70.62 ;
      RECT MASK 2 71.551 70.38 71.611 70.62 ;
      RECT MASK 2 71.991 70.38 72.051 70.62 ;
      RECT MASK 2 72.431 70.38 72.491 70.62 ;
      RECT MASK 2 72.871 70.38 72.931 70.62 ;
      RECT MASK 2 73.311 70.38 73.371 70.62 ;
      RECT MASK 2 73.751 70.38 73.811 70.62 ;
      RECT MASK 2 74.191 70.38 74.251 70.62 ;
      RECT MASK 2 74.631 70.38 74.691 70.62 ;
      RECT MASK 2 75.071 70.38 75.131 70.62 ;
      RECT MASK 2 75.511 70.38 75.571 70.62 ;
      RECT MASK 2 75.951 70.38 76.011 70.62 ;
      RECT MASK 2 76.391 70.38 76.451 70.62 ;
      RECT MASK 2 76.831 70.38 76.891 70.62 ;
      RECT MASK 2 77.729 70.38 77.789 70.62 ;
      RECT MASK 2 78.169 70.38 78.229 70.62 ;
      RECT MASK 2 78.609 70.38 78.669 70.62 ;
      RECT MASK 2 79.049 70.38 79.109 70.62 ;
      RECT MASK 2 79.489 70.38 79.549 70.62 ;
      RECT MASK 2 79.929 70.38 79.989 70.62 ;
      RECT MASK 2 80.369 70.38 80.429 70.62 ;
      RECT MASK 2 80.809 70.38 80.869 70.62 ;
      RECT MASK 2 81.249 70.38 81.309 70.62 ;
      RECT MASK 2 81.689 70.38 81.749 70.62 ;
      RECT MASK 2 82.129 70.38 82.189 70.62 ;
      RECT MASK 2 83.449 70.38 83.509 70.62 ;
      RECT MASK 2 84.347 70.38 84.407 70.62 ;
      RECT MASK 2 84.787 70.38 84.847 70.62 ;
      RECT MASK 2 85.227 70.38 85.287 70.62 ;
      RECT MASK 2 85.667 70.38 85.727 70.62 ;
      RECT MASK 2 86.107 70.38 86.167 70.62 ;
      RECT MASK 2 86.547 70.38 86.607 70.62 ;
      RECT MASK 2 86.987 70.38 87.047 70.62 ;
      RECT MASK 2 87.427 70.38 87.487 70.62 ;
      RECT MASK 2 87.867 70.38 87.927 70.62 ;
      RECT MASK 2 88.307 70.38 88.367 70.62 ;
      RECT MASK 2 88.747 70.38 88.807 70.62 ;
      RECT MASK 2 89.187 70.38 89.247 70.62 ;
      RECT MASK 2 89.627 70.38 89.687 70.62 ;
      RECT MASK 2 90.067 70.38 90.127 70.62 ;
      RECT MASK 2 90.965 70.38 91.025 70.62 ;
      RECT MASK 2 91.405 70.38 91.465 70.62 ;
      RECT MASK 2 91.845 70.38 91.905 70.62 ;
      RECT MASK 2 92.285 70.38 92.345 70.62 ;
      RECT MASK 2 92.725 70.38 92.785 70.62 ;
      RECT MASK 2 93.165 70.38 93.225 70.62 ;
      RECT MASK 2 93.605 70.38 93.665 70.62 ;
      RECT MASK 2 94.045 70.38 94.105 70.62 ;
      RECT MASK 2 94.485 70.38 94.545 70.62 ;
      RECT MASK 2 94.925 70.38 94.985 70.62 ;
      RECT MASK 2 95.365 70.38 95.425 70.62 ;
      RECT MASK 2 95.805 70.38 95.865 70.62 ;
      RECT MASK 2 96.245 70.38 96.305 70.62 ;
      RECT MASK 2 96.685 70.38 96.745 70.62 ;
      RECT MASK 2 97.583 70.38 97.643 70.62 ;
      RECT MASK 2 98.023 70.38 98.083 70.62 ;
      RECT MASK 2 98.463 70.38 98.523 70.62 ;
      RECT MASK 2 98.903 70.38 98.963 70.62 ;
      RECT MASK 2 99.343 70.38 99.403 70.62 ;
      RECT MASK 2 99.783 70.38 99.843 70.62 ;
      RECT MASK 2 100.223 70.38 100.283 70.62 ;
      RECT MASK 2 100.663 70.38 100.723 70.62 ;
      RECT MASK 2 101.103 70.38 101.163 70.62 ;
      RECT MASK 2 101.543 70.38 101.603 70.62 ;
      RECT MASK 2 101.983 70.38 102.043 70.62 ;
      RECT MASK 2 102.423 70.38 102.483 70.62 ;
      RECT MASK 2 102.863 70.38 102.923 70.62 ;
      RECT MASK 2 103.303 70.38 103.363 70.62 ;
      RECT MASK 2 104.201 70.38 104.261 70.62 ;
      RECT MASK 2 104.641 70.38 104.701 70.62 ;
      RECT MASK 2 105.081 70.38 105.141 70.62 ;
      RECT MASK 2 105.521 70.38 105.581 70.62 ;
      RECT MASK 2 105.961 70.38 106.021 70.62 ;
      RECT MASK 2 106.401 70.38 106.461 70.62 ;
      RECT MASK 2 106.841 70.38 106.901 70.62 ;
      RECT MASK 2 107.281 70.38 107.341 70.62 ;
      RECT MASK 2 107.721 70.38 107.781 70.62 ;
      RECT MASK 2 108.161 70.38 108.221 70.62 ;
      RECT MASK 2 108.601 70.38 108.661 70.62 ;
      RECT MASK 2 109.041 70.38 109.101 70.62 ;
      RECT MASK 2 109.481 70.38 109.541 70.62 ;
      RECT MASK 2 109.921 70.38 109.981 70.62 ;
      RECT MASK 2 4.901 70.819 5.021 75.911 ;
      RECT MASK 2 5.341 70.819 5.461 75.911 ;
      RECT MASK 2 5.781 70.819 5.901 75.911 ;
      RECT MASK 2 6.221 70.819 6.341 75.911 ;
      RECT MASK 2 6.661 70.819 6.781 75.911 ;
      RECT MASK 2 7.101 70.819 7.221 75.911 ;
      RECT MASK 2 7.541 70.819 7.661 75.911 ;
      RECT MASK 2 7.981 70.819 8.101 75.911 ;
      RECT MASK 2 8.421 70.819 8.541 75.911 ;
      RECT MASK 2 8.861 70.819 8.981 75.911 ;
      RECT MASK 2 9.301 70.819 9.421 75.911 ;
      RECT MASK 2 9.741 70.819 9.861 75.911 ;
      RECT MASK 2 10.181 70.819 10.301 75.911 ;
      RECT MASK 2 10.621 70.819 10.741 75.911 ;
      RECT MASK 2 11.519 70.819 11.639 75.911 ;
      RECT MASK 2 11.959 70.819 12.079 75.911 ;
      RECT MASK 2 12.399 70.819 12.519 75.911 ;
      RECT MASK 2 12.839 70.819 12.959 75.911 ;
      RECT MASK 2 13.279 70.819 13.399 75.911 ;
      RECT MASK 2 13.719 70.819 13.839 75.911 ;
      RECT MASK 2 14.159 70.819 14.279 75.911 ;
      RECT MASK 2 14.599 70.819 14.719 75.911 ;
      RECT MASK 2 15.039 70.819 15.159 75.911 ;
      RECT MASK 2 15.479 70.819 15.599 75.911 ;
      RECT MASK 2 15.919 70.819 16.039 75.911 ;
      RECT MASK 2 16.359 70.819 16.479 75.911 ;
      RECT MASK 2 16.799 70.819 16.919 75.911 ;
      RECT MASK 2 17.239 70.819 17.359 75.911 ;
      RECT MASK 2 18.137 70.819 18.257 75.911 ;
      RECT MASK 2 18.577 70.819 18.697 75.911 ;
      RECT MASK 2 19.017 70.819 19.137 75.911 ;
      RECT MASK 2 19.457 70.819 19.577 75.911 ;
      RECT MASK 2 19.897 70.819 20.017 75.911 ;
      RECT MASK 2 20.337 70.819 20.457 75.911 ;
      RECT MASK 2 20.777 70.819 20.897 75.911 ;
      RECT MASK 2 21.217 70.819 21.337 75.911 ;
      RECT MASK 2 21.657 70.819 21.777 75.911 ;
      RECT MASK 2 22.097 70.819 22.217 75.911 ;
      RECT MASK 2 22.537 70.819 22.657 75.911 ;
      RECT MASK 2 22.977 70.819 23.097 75.911 ;
      RECT MASK 2 23.417 70.819 23.537 75.911 ;
      RECT MASK 2 23.857 70.819 23.977 75.911 ;
      RECT MASK 2 24.755 70.819 24.875 75.911 ;
      RECT MASK 2 25.195 70.819 25.315 75.911 ;
      RECT MASK 2 25.635 70.819 25.755 75.911 ;
      RECT MASK 2 26.075 70.819 26.195 75.911 ;
      RECT MASK 2 26.515 70.819 26.635 75.911 ;
      RECT MASK 2 26.955 70.819 27.075 75.911 ;
      RECT MASK 2 27.395 70.819 27.515 75.911 ;
      RECT MASK 2 27.835 70.819 27.955 75.911 ;
      RECT MASK 2 28.275 70.819 28.395 75.911 ;
      RECT MASK 2 28.715 70.819 28.835 75.911 ;
      RECT MASK 2 29.155 70.819 29.275 75.911 ;
      RECT MASK 2 29.595 70.819 29.715 75.911 ;
      RECT MASK 2 30.035 70.819 30.155 75.911 ;
      RECT MASK 2 30.475 70.819 30.595 75.911 ;
      RECT MASK 2 31.373 70.819 31.493 75.911 ;
      RECT MASK 2 31.813 70.819 31.933 75.911 ;
      RECT MASK 2 32.253 70.819 32.373 75.911 ;
      RECT MASK 2 32.693 70.819 32.813 75.911 ;
      RECT MASK 2 33.133 70.819 33.253 75.911 ;
      RECT MASK 2 33.573 70.819 33.693 75.911 ;
      RECT MASK 2 34.013 70.819 34.133 75.911 ;
      RECT MASK 2 34.453 70.819 34.573 75.911 ;
      RECT MASK 2 34.893 70.819 35.013 75.911 ;
      RECT MASK 2 35.333 70.819 35.453 75.911 ;
      RECT MASK 2 35.773 70.819 35.893 75.911 ;
      RECT MASK 2 36.213 70.819 36.333 75.911 ;
      RECT MASK 2 36.653 70.819 36.773 75.911 ;
      RECT MASK 2 37.093 70.819 37.213 75.911 ;
      RECT MASK 2 37.991 70.819 38.111 75.911 ;
      RECT MASK 2 38.431 70.819 38.551 75.911 ;
      RECT MASK 2 38.871 70.819 38.991 75.911 ;
      RECT MASK 2 39.311 70.819 39.431 75.911 ;
      RECT MASK 2 39.751 70.819 39.871 75.911 ;
      RECT MASK 2 40.191 70.819 40.311 75.911 ;
      RECT MASK 2 40.631 70.819 40.751 75.911 ;
      RECT MASK 2 41.071 70.819 41.191 75.911 ;
      RECT MASK 2 41.511 70.819 41.631 75.911 ;
      RECT MASK 2 41.951 70.819 42.071 75.911 ;
      RECT MASK 2 42.391 70.819 42.511 75.911 ;
      RECT MASK 2 42.831 70.819 42.951 75.911 ;
      RECT MASK 2 43.271 70.819 43.391 75.911 ;
      RECT MASK 2 43.711 70.819 43.831 75.911 ;
      RECT MASK 2 44.609 70.819 44.729 75.911 ;
      RECT MASK 2 45.049 70.819 45.169 75.911 ;
      RECT MASK 2 45.489 70.819 45.609 75.911 ;
      RECT MASK 2 45.929 70.819 46.049 75.911 ;
      RECT MASK 2 46.369 70.819 46.489 75.911 ;
      RECT MASK 2 46.809 70.819 46.929 75.911 ;
      RECT MASK 2 47.249 70.819 47.369 75.911 ;
      RECT MASK 2 47.689 70.819 47.809 75.911 ;
      RECT MASK 2 48.129 70.819 48.249 75.911 ;
      RECT MASK 2 48.569 70.819 48.689 75.911 ;
      RECT MASK 2 49.009 70.819 49.129 75.911 ;
      RECT MASK 2 49.449 70.819 49.569 75.911 ;
      RECT MASK 2 49.889 70.819 50.009 75.911 ;
      RECT MASK 2 50.329 70.819 50.449 75.911 ;
      RECT MASK 2 51.227 70.819 51.347 75.911 ;
      RECT MASK 2 51.667 70.819 51.787 75.911 ;
      RECT MASK 2 52.107 70.819 52.227 75.911 ;
      RECT MASK 2 52.547 70.819 52.667 75.911 ;
      RECT MASK 2 52.987 70.819 53.107 75.911 ;
      RECT MASK 2 53.427 70.819 53.547 75.911 ;
      RECT MASK 2 53.867 70.819 53.987 75.911 ;
      RECT MASK 2 54.307 70.819 54.427 75.911 ;
      RECT MASK 2 54.747 70.819 54.867 75.911 ;
      RECT MASK 2 55.187 70.819 55.307 75.911 ;
      RECT MASK 2 55.627 70.819 55.747 75.911 ;
      RECT MASK 2 56.067 70.819 56.187 75.911 ;
      RECT MASK 2 56.507 70.819 56.627 75.911 ;
      RECT MASK 2 56.947 70.819 57.067 75.911 ;
      RECT MASK 2 57.845 70.819 57.965 75.911 ;
      RECT MASK 2 58.285 70.819 58.405 75.911 ;
      RECT MASK 2 58.725 70.819 58.845 75.911 ;
      RECT MASK 2 59.165 70.819 59.285 75.911 ;
      RECT MASK 2 59.605 70.819 59.725 75.911 ;
      RECT MASK 2 60.045 70.819 60.165 75.911 ;
      RECT MASK 2 60.485 70.819 60.605 75.911 ;
      RECT MASK 2 60.925 70.819 61.045 75.911 ;
      RECT MASK 2 61.365 70.819 61.485 75.911 ;
      RECT MASK 2 61.805 70.819 61.925 75.911 ;
      RECT MASK 2 62.245 70.819 62.365 75.911 ;
      RECT MASK 2 62.685 70.819 62.805 75.911 ;
      RECT MASK 2 63.125 70.819 63.245 75.911 ;
      RECT MASK 2 63.565 70.819 63.685 75.911 ;
      RECT MASK 2 64.463 70.819 64.583 75.911 ;
      RECT MASK 2 64.903 70.819 65.023 75.911 ;
      RECT MASK 2 65.343 70.819 65.463 75.911 ;
      RECT MASK 2 65.783 70.819 65.903 75.911 ;
      RECT MASK 2 66.223 70.819 66.343 75.911 ;
      RECT MASK 2 66.663 70.819 66.783 75.911 ;
      RECT MASK 2 67.103 70.819 67.223 75.911 ;
      RECT MASK 2 67.543 70.819 67.663 75.911 ;
      RECT MASK 2 67.983 70.819 68.103 75.911 ;
      RECT MASK 2 68.423 70.819 68.543 75.911 ;
      RECT MASK 2 68.863 70.819 68.983 75.911 ;
      RECT MASK 2 69.303 70.819 69.423 75.911 ;
      RECT MASK 2 69.743 70.819 69.863 75.911 ;
      RECT MASK 2 70.183 70.819 70.303 75.911 ;
      RECT MASK 2 71.081 70.819 71.201 75.911 ;
      RECT MASK 2 71.521 70.819 71.641 75.911 ;
      RECT MASK 2 71.961 70.819 72.081 75.911 ;
      RECT MASK 2 72.401 70.819 72.521 75.911 ;
      RECT MASK 2 72.841 70.819 72.961 75.911 ;
      RECT MASK 2 73.281 70.819 73.401 75.911 ;
      RECT MASK 2 73.721 70.819 73.841 75.911 ;
      RECT MASK 2 74.161 70.819 74.281 75.911 ;
      RECT MASK 2 74.601 70.819 74.721 75.911 ;
      RECT MASK 2 75.041 70.819 75.161 75.911 ;
      RECT MASK 2 75.481 70.819 75.601 75.911 ;
      RECT MASK 2 75.921 70.819 76.041 75.911 ;
      RECT MASK 2 76.361 70.819 76.481 75.911 ;
      RECT MASK 2 76.801 70.819 76.921 75.911 ;
      RECT MASK 2 77.699 70.819 77.819 75.911 ;
      RECT MASK 2 78.139 70.819 78.259 75.911 ;
      RECT MASK 2 78.579 70.819 78.699 75.911 ;
      RECT MASK 2 79.019 70.819 79.139 75.911 ;
      RECT MASK 2 79.459 70.819 79.579 75.911 ;
      RECT MASK 2 79.899 70.819 80.019 75.911 ;
      RECT MASK 2 80.339 70.819 80.459 75.911 ;
      RECT MASK 2 80.779 70.819 80.899 75.911 ;
      RECT MASK 2 81.219 70.819 81.339 75.911 ;
      RECT MASK 2 81.659 70.819 81.779 75.911 ;
      RECT MASK 2 82.099 70.819 82.219 75.911 ;
      RECT MASK 2 82.539 70.819 82.659 75.911 ;
      RECT MASK 2 82.979 70.819 83.099 75.911 ;
      RECT MASK 2 83.419 70.819 83.539 75.911 ;
      RECT MASK 2 84.317 70.819 84.437 75.911 ;
      RECT MASK 2 84.757 70.819 84.877 75.911 ;
      RECT MASK 2 85.197 70.819 85.317 75.911 ;
      RECT MASK 2 85.637 70.819 85.757 75.911 ;
      RECT MASK 2 86.077 70.819 86.197 75.911 ;
      RECT MASK 2 86.517 70.819 86.637 75.911 ;
      RECT MASK 2 86.957 70.819 87.077 75.911 ;
      RECT MASK 2 87.397 70.819 87.517 75.911 ;
      RECT MASK 2 87.837 70.819 87.957 75.911 ;
      RECT MASK 2 88.277 70.819 88.397 75.911 ;
      RECT MASK 2 88.717 70.819 88.837 75.911 ;
      RECT MASK 2 89.157 70.819 89.277 75.911 ;
      RECT MASK 2 89.597 70.819 89.717 75.911 ;
      RECT MASK 2 90.037 70.819 90.157 75.911 ;
      RECT MASK 2 90.935 70.819 91.055 75.911 ;
      RECT MASK 2 91.375 70.819 91.495 75.911 ;
      RECT MASK 2 91.815 70.819 91.935 75.911 ;
      RECT MASK 2 92.255 70.819 92.375 75.911 ;
      RECT MASK 2 92.695 70.819 92.815 75.911 ;
      RECT MASK 2 93.135 70.819 93.255 75.911 ;
      RECT MASK 2 93.575 70.819 93.695 75.911 ;
      RECT MASK 2 94.015 70.819 94.135 75.911 ;
      RECT MASK 2 94.455 70.819 94.575 75.911 ;
      RECT MASK 2 94.895 70.819 95.015 75.911 ;
      RECT MASK 2 95.335 70.819 95.455 75.911 ;
      RECT MASK 2 95.775 70.819 95.895 75.911 ;
      RECT MASK 2 96.215 70.819 96.335 75.911 ;
      RECT MASK 2 96.655 70.819 96.775 75.911 ;
      RECT MASK 2 97.553 70.819 97.673 75.911 ;
      RECT MASK 2 97.993 70.819 98.113 75.911 ;
      RECT MASK 2 98.433 70.819 98.553 75.911 ;
      RECT MASK 2 98.873 70.819 98.993 75.911 ;
      RECT MASK 2 99.313 70.819 99.433 75.911 ;
      RECT MASK 2 99.753 70.819 99.873 75.911 ;
      RECT MASK 2 100.193 70.819 100.313 75.911 ;
      RECT MASK 2 100.633 70.819 100.753 75.911 ;
      RECT MASK 2 101.073 70.819 101.193 75.911 ;
      RECT MASK 2 101.513 70.819 101.633 75.911 ;
      RECT MASK 2 101.953 70.819 102.073 75.911 ;
      RECT MASK 2 102.393 70.819 102.513 75.911 ;
      RECT MASK 2 102.833 70.819 102.953 75.911 ;
      RECT MASK 2 103.273 70.819 103.393 75.911 ;
      RECT MASK 2 104.171 70.819 104.291 75.911 ;
      RECT MASK 2 104.611 70.819 104.731 75.911 ;
      RECT MASK 2 105.051 70.819 105.171 75.911 ;
      RECT MASK 2 105.491 70.819 105.611 75.911 ;
      RECT MASK 2 105.931 70.819 106.051 75.911 ;
      RECT MASK 2 106.371 70.819 106.491 75.911 ;
      RECT MASK 2 106.811 70.819 106.931 75.911 ;
      RECT MASK 2 107.251 70.819 107.371 75.911 ;
      RECT MASK 2 107.691 70.819 107.811 75.911 ;
      RECT MASK 2 108.131 70.819 108.251 75.911 ;
      RECT MASK 2 108.571 70.819 108.691 75.911 ;
      RECT MASK 2 109.011 70.819 109.131 75.911 ;
      RECT MASK 2 109.451 70.819 109.571 75.911 ;
      RECT MASK 2 109.891 70.819 110.011 75.911 ;
      RECT MASK 2 114.553 72.236 114.633 72.544 ;
      RECT MASK 2 114.885 72.236 114.965 72.932 ;
      RECT MASK 2 115.217 72.236 115.297 72.932 ;
      RECT MASK 2 115.549 72.236 115.629 72.932 ;
      RECT MASK 2 115.881 72.236 115.961 72.932 ;
      RECT MASK 2 116.213 72.236 116.293 72.544 ;
      RECT MASK 2 116.545 72.236 116.625 72.544 ;
      RECT MASK 2 116.877 72.236 116.957 72.544 ;
      RECT MASK 2 117.209 72.236 117.289 72.544 ;
      RECT MASK 2 117.541 72.236 117.621 72.544 ;
      RECT MASK 2 117.873 72.236 117.953 72.544 ;
      RECT MASK 2 118.205 72.236 118.285 72.544 ;
      RECT MASK 2 118.537 72.236 118.617 72.544 ;
      RECT MASK 2 118.869 72.236 118.949 72.544 ;
      RECT MASK 2 119.201 72.236 119.281 72.544 ;
      RECT MASK 2 119.533 72.236 119.613 72.544 ;
      RECT MASK 2 119.865 72.236 119.945 72.544 ;
      RECT MASK 2 120.197 72.236 120.277 72.544 ;
      RECT MASK 2 120.529 72.236 120.609 72.544 ;
      RECT MASK 2 120.861 72.236 120.941 72.544 ;
      RECT MASK 2 121.193 72.236 121.273 72.544 ;
      RECT MASK 2 121.525 72.236 121.605 72.544 ;
      RECT MASK 2 121.857 72.236 121.937 72.544 ;
      RECT MASK 2 122.189 72.236 122.269 72.544 ;
      RECT MASK 2 122.521 72.236 122.601 72.544 ;
      RECT MASK 2 122.853 72.236 122.933 72.544 ;
      RECT MASK 2 123.185 72.236 123.265 72.544 ;
      RECT MASK 2 123.517 72.236 123.597 72.544 ;
      RECT MASK 2 123.849 72.236 123.929 72.544 ;
      RECT MASK 2 125.509 72.236 125.589 72.544 ;
      RECT MASK 2 125.841 72.236 125.921 72.544 ;
      RECT MASK 2 126.173 72.236 126.253 72.544 ;
      RECT MASK 2 126.837 72.236 126.917 72.544 ;
      RECT MASK 2 127.501 72.236 127.581 72.544 ;
      RECT MASK 2 127.833 72.236 127.913 72.544 ;
      RECT MASK 2 128.165 72.236 128.245 72.544 ;
      RECT MASK 2 128.497 72.236 128.577 72.544 ;
      RECT MASK 2 115.539 73.196 115.659 80.458 ;
      RECT MASK 2 116.427 73.196 116.507 73.528 ;
      RECT MASK 2 116.759 73.196 116.839 73.528 ;
      RECT MASK 2 117.091 73.196 117.171 73.528 ;
      RECT MASK 2 117.423 73.196 117.503 73.528 ;
      RECT MASK 2 117.755 73.196 117.835 73.528 ;
      RECT MASK 2 118.087 73.196 118.167 73.528 ;
      RECT MASK 2 118.419 73.196 118.499 73.528 ;
      RECT MASK 2 118.751 73.196 118.831 73.528 ;
      RECT MASK 2 119.083 73.196 119.163 73.528 ;
      RECT MASK 2 119.415 73.196 119.495 73.528 ;
      RECT MASK 2 119.747 73.196 119.827 73.528 ;
      RECT MASK 2 120.079 73.196 120.159 73.528 ;
      RECT MASK 2 120.411 73.196 120.491 73.528 ;
      RECT MASK 2 120.743 73.196 120.823 73.528 ;
      RECT MASK 2 121.075 73.196 121.155 73.528 ;
      RECT MASK 2 121.407 73.196 121.487 73.528 ;
      RECT MASK 2 121.739 73.196 121.819 73.528 ;
      RECT MASK 2 122.071 73.196 122.151 73.528 ;
      RECT MASK 2 122.403 73.196 122.483 73.528 ;
      RECT MASK 2 122.735 73.196 122.815 73.528 ;
      RECT MASK 2 123.067 73.196 123.147 73.528 ;
      RECT MASK 2 123.399 73.196 123.479 73.528 ;
      RECT MASK 2 123.731 73.196 123.811 73.528 ;
      RECT MASK 2 124.063 73.196 124.143 73.528 ;
      RECT MASK 2 124.727 73.196 124.807 73.528 ;
      RECT MASK 2 125.391 73.196 125.471 73.528 ;
      RECT MASK 2 125.723 73.196 125.803 73.528 ;
      RECT MASK 2 126.055 73.196 126.135 73.528 ;
      RECT MASK 2 126.827 73.196 126.947 80.4615 ;
      RECT MASK 2 116.427 73.74 116.507 79.672 ;
      RECT MASK 2 116.759 73.74 116.839 79.672 ;
      RECT MASK 2 117.091 73.74 117.171 79.672 ;
      RECT MASK 2 117.423 73.74 117.503 79.672 ;
      RECT MASK 2 117.755 73.74 117.835 79.672 ;
      RECT MASK 2 118.087 73.74 118.167 79.672 ;
      RECT MASK 2 118.419 73.74 118.499 79.672 ;
      RECT MASK 2 118.751 73.74 118.831 79.672 ;
      RECT MASK 2 119.083 73.74 119.163 79.672 ;
      RECT MASK 2 119.415 73.74 119.495 79.672 ;
      RECT MASK 2 119.747 73.74 119.827 79.672 ;
      RECT MASK 2 120.079 73.74 120.159 79.672 ;
      RECT MASK 2 120.411 73.74 120.491 79.672 ;
      RECT MASK 2 120.743 73.74 120.823 79.672 ;
      RECT MASK 2 121.075 73.74 121.155 79.672 ;
      RECT MASK 2 121.407 73.74 121.487 79.672 ;
      RECT MASK 2 121.739 73.74 121.819 79.672 ;
      RECT MASK 2 122.071 73.74 122.151 79.672 ;
      RECT MASK 2 122.403 73.74 122.483 79.672 ;
      RECT MASK 2 122.735 73.74 122.815 79.672 ;
      RECT MASK 2 123.067 73.74 123.147 79.672 ;
      RECT MASK 2 123.399 73.74 123.479 79.672 ;
      RECT MASK 2 123.731 73.74 123.811 79.672 ;
      RECT MASK 2 124.063 73.74 124.143 79.672 ;
      RECT MASK 2 124.395 73.74 124.475 79.672 ;
      RECT MASK 2 124.727 73.74 124.807 79.672 ;
      RECT MASK 2 125.059 73.74 125.139 79.672 ;
      RECT MASK 2 125.391 73.74 125.471 79.672 ;
      RECT MASK 2 125.723 73.74 125.803 79.672 ;
      RECT MASK 2 126.055 73.74 126.135 79.672 ;
      RECT MASK 2 1.839 77.486 1.919 77.818 ;
      RECT MASK 2 2.171 77.486 2.251 77.818 ;
      RECT MASK 2 2.503 77.486 2.583 77.818 ;
      RECT MASK 2 4.163 77.486 4.243 77.818 ;
      RECT MASK 2 4.495 77.486 4.575 77.818 ;
      RECT MASK 2 4.827 77.486 4.907 77.818 ;
      RECT MASK 2 5.159 77.486 5.239 77.818 ;
      RECT MASK 2 5.491 77.486 5.571 77.818 ;
      RECT MASK 2 5.823 77.486 5.903 77.818 ;
      RECT MASK 2 6.155 77.486 6.235 77.818 ;
      RECT MASK 2 6.487 77.486 6.567 77.818 ;
      RECT MASK 2 6.819 77.486 6.899 77.818 ;
      RECT MASK 2 7.151 77.486 7.231 77.818 ;
      RECT MASK 2 7.483 77.486 7.563 77.818 ;
      RECT MASK 2 7.815 77.486 7.895 77.818 ;
      RECT MASK 2 8.147 77.486 8.227 77.818 ;
      RECT MASK 2 8.479 77.486 8.559 77.818 ;
      RECT MASK 2 8.811 77.486 8.891 77.818 ;
      RECT MASK 2 9.143 77.486 9.223 77.818 ;
      RECT MASK 2 9.475 77.486 9.555 77.818 ;
      RECT MASK 2 9.807 77.486 9.887 77.818 ;
      RECT MASK 2 10.139 77.486 10.219 77.818 ;
      RECT MASK 2 10.471 77.486 10.551 77.818 ;
      RECT MASK 2 10.803 77.486 10.883 77.818 ;
      RECT MASK 2 11.135 77.486 11.215 77.818 ;
      RECT MASK 2 11.467 77.486 11.547 77.818 ;
      RECT MASK 2 11.799 77.486 11.879 77.818 ;
      RECT MASK 2 12.131 77.486 12.211 77.818 ;
      RECT MASK 2 12.463 77.486 12.543 77.818 ;
      RECT MASK 2 12.795 77.486 12.875 77.818 ;
      RECT MASK 2 13.127 77.486 13.207 77.818 ;
      RECT MASK 2 13.459 77.486 13.539 77.818 ;
      RECT MASK 2 13.791 77.486 13.871 77.818 ;
      RECT MASK 2 14.123 77.486 14.203 77.818 ;
      RECT MASK 2 14.455 77.486 14.535 77.818 ;
      RECT MASK 2 14.787 77.486 14.867 77.818 ;
      RECT MASK 2 15.119 77.486 15.199 77.818 ;
      RECT MASK 2 15.451 77.486 15.531 77.818 ;
      RECT MASK 2 15.783 77.486 15.863 77.818 ;
      RECT MASK 2 16.115 77.486 16.195 77.818 ;
      RECT MASK 2 16.447 77.486 16.527 77.818 ;
      RECT MASK 2 16.779 77.486 16.859 77.818 ;
      RECT MASK 2 17.111 77.486 17.191 77.818 ;
      RECT MASK 2 17.443 77.486 17.523 77.818 ;
      RECT MASK 2 17.775 77.486 17.855 77.818 ;
      RECT MASK 2 18.107 77.486 18.187 77.818 ;
      RECT MASK 2 18.439 77.486 18.519 77.818 ;
      RECT MASK 2 18.771 77.486 18.851 77.818 ;
      RECT MASK 2 19.103 77.486 19.183 77.818 ;
      RECT MASK 2 19.435 77.486 19.515 77.818 ;
      RECT MASK 2 19.767 77.486 19.847 77.818 ;
      RECT MASK 2 20.099 77.486 20.179 77.818 ;
      RECT MASK 2 20.431 77.486 20.511 77.818 ;
      RECT MASK 2 20.763 77.486 20.843 77.818 ;
      RECT MASK 2 21.095 77.486 21.175 77.818 ;
      RECT MASK 2 21.427 77.486 21.507 77.818 ;
      RECT MASK 2 21.759 77.486 21.839 77.818 ;
      RECT MASK 2 22.091 77.486 22.171 77.818 ;
      RECT MASK 2 22.423 77.486 22.503 77.818 ;
      RECT MASK 2 22.755 77.486 22.835 77.818 ;
      RECT MASK 2 23.087 77.486 23.167 77.818 ;
      RECT MASK 2 23.419 77.486 23.499 77.818 ;
      RECT MASK 2 23.751 77.486 23.831 77.818 ;
      RECT MASK 2 24.083 77.486 24.163 77.818 ;
      RECT MASK 2 24.415 77.486 24.495 77.818 ;
      RECT MASK 2 24.747 77.486 24.827 77.818 ;
      RECT MASK 2 25.079 77.486 25.159 77.818 ;
      RECT MASK 2 25.411 77.486 25.491 77.818 ;
      RECT MASK 2 25.743 77.486 25.823 77.818 ;
      RECT MASK 2 26.075 77.486 26.155 77.818 ;
      RECT MASK 2 26.407 77.486 26.487 77.818 ;
      RECT MASK 2 26.739 77.486 26.819 77.818 ;
      RECT MASK 2 27.071 77.486 27.151 77.818 ;
      RECT MASK 2 27.403 77.486 27.483 77.818 ;
      RECT MASK 2 27.735 77.486 27.815 77.818 ;
      RECT MASK 2 28.067 77.486 28.147 77.818 ;
      RECT MASK 2 28.399 77.486 28.479 77.818 ;
      RECT MASK 2 28.731 77.486 28.811 77.818 ;
      RECT MASK 2 29.063 77.486 29.143 77.818 ;
      RECT MASK 2 29.395 77.486 29.475 77.818 ;
      RECT MASK 2 29.727 77.486 29.807 77.818 ;
      RECT MASK 2 30.059 77.486 30.139 77.818 ;
      RECT MASK 2 30.391 77.486 30.471 77.818 ;
      RECT MASK 2 30.723 77.486 30.803 77.818 ;
      RECT MASK 2 31.055 77.486 31.135 77.818 ;
      RECT MASK 2 31.387 77.486 31.467 77.818 ;
      RECT MASK 2 31.719 77.486 31.799 77.818 ;
      RECT MASK 2 32.051 77.486 32.131 77.818 ;
      RECT MASK 2 32.383 77.486 32.463 77.818 ;
      RECT MASK 2 32.715 77.486 32.795 77.818 ;
      RECT MASK 2 33.047 77.486 33.127 77.818 ;
      RECT MASK 2 33.379 77.486 33.459 77.818 ;
      RECT MASK 2 33.711 77.486 33.791 77.818 ;
      RECT MASK 2 34.043 77.486 34.123 77.818 ;
      RECT MASK 2 34.375 77.486 34.455 77.818 ;
      RECT MASK 2 34.707 77.486 34.787 77.818 ;
      RECT MASK 2 35.039 77.486 35.119 77.818 ;
      RECT MASK 2 35.371 77.486 35.451 77.818 ;
      RECT MASK 2 35.703 77.486 35.783 77.818 ;
      RECT MASK 2 36.035 77.486 36.115 77.818 ;
      RECT MASK 2 36.367 77.486 36.447 77.818 ;
      RECT MASK 2 36.699 77.486 36.779 77.818 ;
      RECT MASK 2 37.031 77.486 37.111 77.818 ;
      RECT MASK 2 37.363 77.486 37.443 77.818 ;
      RECT MASK 2 37.695 77.486 37.775 77.818 ;
      RECT MASK 2 38.027 77.486 38.107 77.818 ;
      RECT MASK 2 38.359 77.486 38.439 77.818 ;
      RECT MASK 2 38.691 77.486 38.771 77.818 ;
      RECT MASK 2 39.023 77.486 39.103 77.818 ;
      RECT MASK 2 39.355 77.486 39.435 77.818 ;
      RECT MASK 2 39.687 77.486 39.767 77.818 ;
      RECT MASK 2 40.019 77.486 40.099 77.818 ;
      RECT MASK 2 40.351 77.486 40.431 77.818 ;
      RECT MASK 2 40.683 77.486 40.763 77.818 ;
      RECT MASK 2 41.015 77.486 41.095 77.818 ;
      RECT MASK 2 41.347 77.486 41.427 77.818 ;
      RECT MASK 2 41.679 77.486 41.759 77.818 ;
      RECT MASK 2 42.011 77.486 42.091 77.818 ;
      RECT MASK 2 42.343 77.486 42.423 77.818 ;
      RECT MASK 2 42.675 77.486 42.755 77.818 ;
      RECT MASK 2 43.007 77.486 43.087 77.818 ;
      RECT MASK 2 43.339 77.486 43.419 77.818 ;
      RECT MASK 2 43.671 77.486 43.751 77.818 ;
      RECT MASK 2 44.003 77.486 44.083 77.818 ;
      RECT MASK 2 44.335 77.486 44.415 77.818 ;
      RECT MASK 2 44.667 77.486 44.747 77.818 ;
      RECT MASK 2 44.999 77.486 45.079 77.818 ;
      RECT MASK 2 45.331 77.486 45.411 77.818 ;
      RECT MASK 2 45.663 77.486 45.743 77.818 ;
      RECT MASK 2 45.995 77.486 46.075 77.818 ;
      RECT MASK 2 46.327 77.486 46.407 77.818 ;
      RECT MASK 2 46.659 77.486 46.739 77.818 ;
      RECT MASK 2 46.991 77.486 47.071 77.818 ;
      RECT MASK 2 47.323 77.486 47.403 77.818 ;
      RECT MASK 2 47.655 77.486 47.735 77.818 ;
      RECT MASK 2 47.987 77.486 48.067 77.818 ;
      RECT MASK 2 48.319 77.486 48.399 77.818 ;
      RECT MASK 2 48.651 77.486 48.731 77.818 ;
      RECT MASK 2 48.983 77.486 49.063 77.818 ;
      RECT MASK 2 49.315 77.486 49.395 77.818 ;
      RECT MASK 2 49.647 77.486 49.727 77.818 ;
      RECT MASK 2 49.979 77.486 50.059 77.818 ;
      RECT MASK 2 50.311 77.486 50.391 77.818 ;
      RECT MASK 2 50.643 77.486 50.723 77.818 ;
      RECT MASK 2 50.975 77.486 51.055 77.818 ;
      RECT MASK 2 51.307 77.486 51.387 77.818 ;
      RECT MASK 2 51.639 77.486 51.719 77.818 ;
      RECT MASK 2 51.971 77.486 52.051 77.818 ;
      RECT MASK 2 52.303 77.486 52.383 77.818 ;
      RECT MASK 2 52.635 77.486 52.715 77.818 ;
      RECT MASK 2 52.967 77.486 53.047 77.818 ;
      RECT MASK 2 53.299 77.486 53.379 77.818 ;
      RECT MASK 2 53.631 77.486 53.711 77.818 ;
      RECT MASK 2 53.963 77.486 54.043 77.818 ;
      RECT MASK 2 54.295 77.486 54.375 77.818 ;
      RECT MASK 2 54.627 77.486 54.707 77.818 ;
      RECT MASK 2 54.959 77.486 55.039 77.818 ;
      RECT MASK 2 55.291 77.486 55.371 77.818 ;
      RECT MASK 2 55.623 77.486 55.703 77.818 ;
      RECT MASK 2 55.955 77.486 56.035 77.818 ;
      RECT MASK 2 56.287 77.486 56.367 77.818 ;
      RECT MASK 2 56.619 77.486 56.699 77.818 ;
      RECT MASK 2 56.951 77.486 57.031 77.818 ;
      RECT MASK 2 57.283 77.486 57.363 77.818 ;
      RECT MASK 2 57.615 77.486 57.695 77.818 ;
      RECT MASK 2 57.947 77.486 58.027 77.818 ;
      RECT MASK 2 58.279 77.486 58.359 77.818 ;
      RECT MASK 2 58.611 77.486 58.691 77.818 ;
      RECT MASK 2 58.943 77.486 59.023 77.818 ;
      RECT MASK 2 59.275 77.486 59.355 77.818 ;
      RECT MASK 2 59.607 77.486 59.687 77.818 ;
      RECT MASK 2 59.939 77.486 60.019 77.818 ;
      RECT MASK 2 60.271 77.486 60.351 77.818 ;
      RECT MASK 2 60.603 77.486 60.683 77.818 ;
      RECT MASK 2 60.935 77.486 61.015 77.818 ;
      RECT MASK 2 61.267 77.486 61.347 77.818 ;
      RECT MASK 2 61.599 77.486 61.679 77.818 ;
      RECT MASK 2 61.931 77.486 62.011 77.818 ;
      RECT MASK 2 62.263 77.486 62.343 77.818 ;
      RECT MASK 2 62.595 77.486 62.675 77.818 ;
      RECT MASK 2 62.927 77.486 63.007 77.818 ;
      RECT MASK 2 63.259 77.486 63.339 77.818 ;
      RECT MASK 2 63.591 77.486 63.671 77.818 ;
      RECT MASK 2 63.923 77.486 64.003 77.818 ;
      RECT MASK 2 64.255 77.486 64.335 77.818 ;
      RECT MASK 2 64.587 77.486 64.667 77.818 ;
      RECT MASK 2 64.919 77.486 64.999 77.818 ;
      RECT MASK 2 65.251 77.486 65.331 77.818 ;
      RECT MASK 2 65.583 77.486 65.663 77.818 ;
      RECT MASK 2 65.915 77.486 65.995 77.818 ;
      RECT MASK 2 66.247 77.486 66.327 77.818 ;
      RECT MASK 2 66.579 77.486 66.659 77.818 ;
      RECT MASK 2 66.911 77.486 66.991 77.818 ;
      RECT MASK 2 67.243 77.486 67.323 77.818 ;
      RECT MASK 2 67.575 77.486 67.655 77.818 ;
      RECT MASK 2 67.907 77.486 67.987 77.818 ;
      RECT MASK 2 68.239 77.486 68.319 77.818 ;
      RECT MASK 2 68.571 77.486 68.651 77.818 ;
      RECT MASK 2 68.903 77.486 68.983 77.818 ;
      RECT MASK 2 69.235 77.486 69.315 77.818 ;
      RECT MASK 2 69.567 77.486 69.647 77.818 ;
      RECT MASK 2 69.899 77.486 69.979 77.818 ;
      RECT MASK 2 70.231 77.486 70.311 77.818 ;
      RECT MASK 2 70.563 77.486 70.643 77.818 ;
      RECT MASK 2 70.895 77.486 70.975 77.818 ;
      RECT MASK 2 71.227 77.486 71.307 77.818 ;
      RECT MASK 2 71.559 77.486 71.639 77.818 ;
      RECT MASK 2 71.891 77.486 71.971 77.818 ;
      RECT MASK 2 72.223 77.486 72.303 77.818 ;
      RECT MASK 2 72.555 77.486 72.635 77.818 ;
      RECT MASK 2 72.887 77.486 72.967 77.818 ;
      RECT MASK 2 73.219 77.486 73.299 77.818 ;
      RECT MASK 2 73.551 77.486 73.631 77.818 ;
      RECT MASK 2 73.883 77.486 73.963 77.818 ;
      RECT MASK 2 74.215 77.486 74.295 77.818 ;
      RECT MASK 2 74.547 77.486 74.627 77.818 ;
      RECT MASK 2 74.879 77.486 74.959 77.818 ;
      RECT MASK 2 75.211 77.486 75.291 77.818 ;
      RECT MASK 2 75.543 77.486 75.623 77.818 ;
      RECT MASK 2 75.875 77.486 75.955 77.818 ;
      RECT MASK 2 76.207 77.486 76.287 77.818 ;
      RECT MASK 2 76.539 77.486 76.619 77.818 ;
      RECT MASK 2 76.871 77.486 76.951 77.818 ;
      RECT MASK 2 77.203 77.486 77.283 77.818 ;
      RECT MASK 2 77.535 77.486 77.615 77.818 ;
      RECT MASK 2 77.867 77.486 77.947 77.818 ;
      RECT MASK 2 78.199 77.486 78.279 77.818 ;
      RECT MASK 2 78.531 77.486 78.611 77.818 ;
      RECT MASK 2 78.863 77.486 78.943 77.818 ;
      RECT MASK 2 79.195 77.486 79.275 77.818 ;
      RECT MASK 2 79.527 77.486 79.607 77.818 ;
      RECT MASK 2 79.859 77.486 79.939 77.818 ;
      RECT MASK 2 80.191 77.486 80.271 77.818 ;
      RECT MASK 2 80.523 77.486 80.603 77.818 ;
      RECT MASK 2 80.855 77.486 80.935 77.818 ;
      RECT MASK 2 81.187 77.486 81.267 77.818 ;
      RECT MASK 2 81.519 77.486 81.599 77.818 ;
      RECT MASK 2 81.851 77.486 81.931 77.818 ;
      RECT MASK 2 82.183 77.486 82.263 77.818 ;
      RECT MASK 2 82.515 77.486 82.595 77.818 ;
      RECT MASK 2 82.847 77.486 82.927 77.818 ;
      RECT MASK 2 83.179 77.486 83.259 77.818 ;
      RECT MASK 2 83.511 77.486 83.591 77.818 ;
      RECT MASK 2 83.843 77.486 83.923 77.818 ;
      RECT MASK 2 84.175 77.486 84.255 77.818 ;
      RECT MASK 2 84.507 77.486 84.587 77.818 ;
      RECT MASK 2 84.839 77.486 84.919 77.818 ;
      RECT MASK 2 85.171 77.486 85.251 77.818 ;
      RECT MASK 2 85.503 77.486 85.583 77.818 ;
      RECT MASK 2 85.835 77.486 85.915 77.818 ;
      RECT MASK 2 86.167 77.486 86.247 77.818 ;
      RECT MASK 2 86.499 77.486 86.579 77.818 ;
      RECT MASK 2 86.831 77.486 86.911 77.818 ;
      RECT MASK 2 87.163 77.486 87.243 77.818 ;
      RECT MASK 2 87.495 77.486 87.575 77.818 ;
      RECT MASK 2 87.827 77.486 87.907 77.818 ;
      RECT MASK 2 88.159 77.486 88.239 77.818 ;
      RECT MASK 2 88.491 77.486 88.571 77.818 ;
      RECT MASK 2 88.823 77.486 88.903 77.818 ;
      RECT MASK 2 89.155 77.486 89.235 77.818 ;
      RECT MASK 2 89.487 77.486 89.567 77.818 ;
      RECT MASK 2 89.819 77.486 89.899 77.818 ;
      RECT MASK 2 90.151 77.486 90.231 77.818 ;
      RECT MASK 2 90.483 77.486 90.563 77.818 ;
      RECT MASK 2 90.815 77.486 90.895 77.818 ;
      RECT MASK 2 91.147 77.486 91.227 77.818 ;
      RECT MASK 2 91.479 77.486 91.559 77.818 ;
      RECT MASK 2 91.811 77.486 91.891 77.818 ;
      RECT MASK 2 92.143 77.486 92.223 77.818 ;
      RECT MASK 2 92.475 77.486 92.555 77.818 ;
      RECT MASK 2 92.807 77.486 92.887 77.818 ;
      RECT MASK 2 93.139 77.486 93.219 77.818 ;
      RECT MASK 2 93.471 77.486 93.551 77.818 ;
      RECT MASK 2 93.803 77.486 93.883 77.818 ;
      RECT MASK 2 94.135 77.486 94.215 77.818 ;
      RECT MASK 2 94.467 77.486 94.547 77.818 ;
      RECT MASK 2 94.799 77.486 94.879 77.818 ;
      RECT MASK 2 95.131 77.486 95.211 77.818 ;
      RECT MASK 2 95.463 77.486 95.543 77.818 ;
      RECT MASK 2 95.795 77.486 95.875 77.818 ;
      RECT MASK 2 96.127 77.486 96.207 77.818 ;
      RECT MASK 2 96.459 77.486 96.539 77.818 ;
      RECT MASK 2 96.791 77.486 96.871 77.818 ;
      RECT MASK 2 97.123 77.486 97.203 77.818 ;
      RECT MASK 2 97.455 77.486 97.535 77.818 ;
      RECT MASK 2 97.787 77.486 97.867 77.818 ;
      RECT MASK 2 98.119 77.486 98.199 77.818 ;
      RECT MASK 2 98.451 77.486 98.531 77.818 ;
      RECT MASK 2 98.783 77.486 98.863 77.818 ;
      RECT MASK 2 99.115 77.486 99.195 77.818 ;
      RECT MASK 2 99.447 77.486 99.527 77.818 ;
      RECT MASK 2 99.779 77.486 99.859 77.818 ;
      RECT MASK 2 100.111 77.486 100.191 77.818 ;
      RECT MASK 2 100.443 77.486 100.523 77.818 ;
      RECT MASK 2 100.775 77.486 100.855 77.818 ;
      RECT MASK 2 101.107 77.486 101.187 77.818 ;
      RECT MASK 2 101.439 77.486 101.519 77.818 ;
      RECT MASK 2 101.771 77.486 101.851 77.818 ;
      RECT MASK 2 102.103 77.486 102.183 77.818 ;
      RECT MASK 2 102.435 77.486 102.515 77.818 ;
      RECT MASK 2 102.767 77.486 102.847 77.818 ;
      RECT MASK 2 103.099 77.486 103.179 77.818 ;
      RECT MASK 2 103.431 77.486 103.511 77.818 ;
      RECT MASK 2 103.763 77.486 103.843 77.818 ;
      RECT MASK 2 104.095 77.486 104.175 77.818 ;
      RECT MASK 2 104.427 77.486 104.507 77.818 ;
      RECT MASK 2 104.759 77.486 104.839 77.818 ;
      RECT MASK 2 105.091 77.486 105.171 77.818 ;
      RECT MASK 2 105.423 77.486 105.503 77.818 ;
      RECT MASK 2 105.755 77.486 105.835 77.818 ;
      RECT MASK 2 106.087 77.486 106.167 77.818 ;
      RECT MASK 2 106.419 77.486 106.499 77.818 ;
      RECT MASK 2 106.751 77.486 106.831 77.818 ;
      RECT MASK 2 107.083 77.486 107.163 77.818 ;
      RECT MASK 2 107.415 77.486 107.495 77.818 ;
      RECT MASK 2 107.747 77.486 107.827 77.818 ;
      RECT MASK 2 108.079 77.486 108.159 77.818 ;
      RECT MASK 2 108.411 77.486 108.491 77.818 ;
      RECT MASK 2 108.743 77.486 108.823 77.818 ;
      RECT MASK 2 109.075 77.486 109.155 77.818 ;
      RECT MASK 2 109.407 77.486 109.487 77.818 ;
      RECT MASK 2 109.739 77.486 109.819 77.818 ;
      RECT MASK 2 110.071 77.486 110.151 77.818 ;
      RECT MASK 2 110.403 77.486 110.483 77.818 ;
      RECT MASK 2 110.735 77.486 110.815 77.818 ;
      RECT MASK 2 112.395 77.486 112.475 77.818 ;
      RECT MASK 2 112.727 77.486 112.807 77.818 ;
      RECT MASK 2 113.059 77.486 113.139 77.818 ;
      RECT MASK 2 113.391 77.486 113.471 77.818 ;
      RECT MASK 2 6.661 78.03 6.721 78.3 ;
      RECT MASK 2 7.159 78.03 7.219 78.3 ;
      RECT MASK 2 7.491 78.03 7.551 78.3 ;
      RECT MASK 2 7.823 78.03 7.883 78.3 ;
      RECT MASK 2 8.321 78.03 8.381 78.3 ;
      RECT MASK 2 8.653 78.03 8.713 78.3 ;
      RECT MASK 2 8.985 78.03 9.045 78.3 ;
      RECT MASK 2 9.483 78.03 9.543 78.3 ;
      RECT MASK 2 9.815 78.03 9.875 78.3 ;
      RECT MASK 2 10.147 78.03 10.207 78.3 ;
      RECT MASK 2 12.117 78.03 12.177 78.3 ;
      RECT MASK 2 12.615 78.03 12.675 78.3 ;
      RECT MASK 2 12.947 78.03 13.007 78.3 ;
      RECT MASK 2 13.279 78.03 13.339 78.3 ;
      RECT MASK 2 13.777 78.03 13.837 78.3 ;
      RECT MASK 2 14.109 78.03 14.169 78.3 ;
      RECT MASK 2 14.441 78.03 14.501 78.3 ;
      RECT MASK 2 14.939 78.03 14.999 78.3 ;
      RECT MASK 2 15.271 78.03 15.331 78.3 ;
      RECT MASK 2 15.603 78.03 15.663 78.3 ;
      RECT MASK 2 16.101 78.03 16.161 78.3 ;
      RECT MASK 2 16.433 78.03 16.493 78.3 ;
      RECT MASK 2 16.765 78.03 16.825 79.402 ;
      RECT MASK 2 17.501 78.03 17.561 80.25 ;
      RECT MASK 2 17.833 78.03 17.893 80.25 ;
      RECT MASK 2 18.735 78.03 18.795 78.3 ;
      RECT MASK 2 19.233 78.03 19.293 78.3 ;
      RECT MASK 2 19.565 78.03 19.625 78.3 ;
      RECT MASK 2 19.897 78.03 19.957 78.3 ;
      RECT MASK 2 20.395 78.03 20.455 78.3 ;
      RECT MASK 2 20.727 78.03 20.787 78.3 ;
      RECT MASK 2 21.059 78.03 21.119 78.3 ;
      RECT MASK 2 21.557 78.03 21.617 78.3 ;
      RECT MASK 2 21.889 78.03 21.949 78.3 ;
      RECT MASK 2 22.221 78.03 22.281 78.3 ;
      RECT MASK 2 22.719 78.03 22.779 78.3 ;
      RECT MASK 2 23.051 78.03 23.111 78.3 ;
      RECT MASK 2 23.383 78.03 23.443 79.402 ;
      RECT MASK 2 25.353 78.03 25.413 78.3 ;
      RECT MASK 2 25.851 78.03 25.911 78.3 ;
      RECT MASK 2 26.183 78.03 26.243 78.3 ;
      RECT MASK 2 26.515 78.03 26.575 78.3 ;
      RECT MASK 2 27.013 78.03 27.073 78.3 ;
      RECT MASK 2 27.345 78.03 27.405 78.3 ;
      RECT MASK 2 27.677 78.03 27.737 78.3 ;
      RECT MASK 2 28.175 78.03 28.235 78.3 ;
      RECT MASK 2 28.507 78.03 28.567 78.3 ;
      RECT MASK 2 28.839 78.03 28.899 78.3 ;
      RECT MASK 2 29.337 78.03 29.397 78.3 ;
      RECT MASK 2 29.669 78.03 29.729 78.3 ;
      RECT MASK 2 30.001 78.03 30.061 79.402 ;
      RECT MASK 2 31.971 78.03 32.031 78.3 ;
      RECT MASK 2 32.469 78.03 32.529 78.3 ;
      RECT MASK 2 32.801 78.03 32.861 78.3 ;
      RECT MASK 2 33.133 78.03 33.193 78.3 ;
      RECT MASK 2 33.631 78.03 33.691 78.3 ;
      RECT MASK 2 33.963 78.03 34.023 78.3 ;
      RECT MASK 2 34.295 78.03 34.355 78.3 ;
      RECT MASK 2 34.793 78.03 34.853 78.3 ;
      RECT MASK 2 35.125 78.03 35.185 78.3 ;
      RECT MASK 2 35.457 78.03 35.517 78.3 ;
      RECT MASK 2 35.955 78.03 36.015 78.3 ;
      RECT MASK 2 36.287 78.03 36.347 78.3 ;
      RECT MASK 2 36.619 78.03 36.679 79.402 ;
      RECT MASK 2 38.589 78.03 38.649 78.3 ;
      RECT MASK 2 39.087 78.03 39.147 78.3 ;
      RECT MASK 2 39.419 78.03 39.479 78.3 ;
      RECT MASK 2 39.751 78.03 39.811 78.3 ;
      RECT MASK 2 40.249 78.03 40.309 78.3 ;
      RECT MASK 2 40.581 78.03 40.641 78.3 ;
      RECT MASK 2 40.913 78.03 40.973 78.3 ;
      RECT MASK 2 41.411 78.03 41.471 78.3 ;
      RECT MASK 2 41.743 78.03 41.803 78.3 ;
      RECT MASK 2 42.075 78.03 42.135 78.3 ;
      RECT MASK 2 42.573 78.03 42.633 78.3 ;
      RECT MASK 2 42.905 78.03 42.965 78.3 ;
      RECT MASK 2 43.237 78.03 43.297 79.402 ;
      RECT MASK 2 45.207 78.03 45.267 78.3 ;
      RECT MASK 2 45.705 78.03 45.765 78.3 ;
      RECT MASK 2 46.037 78.03 46.097 78.3 ;
      RECT MASK 2 46.369 78.03 46.429 78.3 ;
      RECT MASK 2 46.867 78.03 46.927 78.3 ;
      RECT MASK 2 47.199 78.03 47.259 78.3 ;
      RECT MASK 2 47.531 78.03 47.591 78.3 ;
      RECT MASK 2 48.029 78.03 48.089 78.3 ;
      RECT MASK 2 48.361 78.03 48.421 78.3 ;
      RECT MASK 2 48.693 78.03 48.753 78.3 ;
      RECT MASK 2 49.191 78.03 49.251 78.3 ;
      RECT MASK 2 49.523 78.03 49.583 78.3 ;
      RECT MASK 2 49.855 78.03 49.915 79.402 ;
      RECT MASK 2 51.825 78.03 51.885 78.3 ;
      RECT MASK 2 52.323 78.03 52.383 78.3 ;
      RECT MASK 2 52.655 78.03 52.715 78.3 ;
      RECT MASK 2 52.987 78.03 53.047 78.3 ;
      RECT MASK 2 53.485 78.03 53.545 78.3 ;
      RECT MASK 2 53.817 78.03 53.877 78.3 ;
      RECT MASK 2 54.149 78.03 54.209 78.3 ;
      RECT MASK 2 54.647 78.03 54.707 78.3 ;
      RECT MASK 2 54.979 78.03 55.039 78.3 ;
      RECT MASK 2 55.311 78.03 55.371 78.3 ;
      RECT MASK 2 55.809 78.03 55.869 78.3 ;
      RECT MASK 2 56.141 78.03 56.201 78.3 ;
      RECT MASK 2 56.473 78.03 56.533 79.402 ;
      RECT MASK 2 58.443 78.03 58.503 78.3 ;
      RECT MASK 2 58.941 78.03 59.001 78.3 ;
      RECT MASK 2 59.273 78.03 59.333 78.3 ;
      RECT MASK 2 59.605 78.03 59.665 78.3 ;
      RECT MASK 2 60.103 78.03 60.163 78.3 ;
      RECT MASK 2 60.435 78.03 60.495 78.3 ;
      RECT MASK 2 60.767 78.03 60.827 78.3 ;
      RECT MASK 2 61.265 78.03 61.325 78.3 ;
      RECT MASK 2 61.597 78.03 61.657 78.3 ;
      RECT MASK 2 61.929 78.03 61.989 78.3 ;
      RECT MASK 2 62.427 78.03 62.487 78.3 ;
      RECT MASK 2 62.759 78.03 62.819 78.3 ;
      RECT MASK 2 63.091 78.03 63.151 79.402 ;
      RECT MASK 2 65.061 78.03 65.121 78.3 ;
      RECT MASK 2 65.559 78.03 65.619 78.3 ;
      RECT MASK 2 65.891 78.03 65.951 78.3 ;
      RECT MASK 2 66.223 78.03 66.283 78.3 ;
      RECT MASK 2 66.721 78.03 66.781 78.3 ;
      RECT MASK 2 67.053 78.03 67.113 78.3 ;
      RECT MASK 2 67.385 78.03 67.445 78.3 ;
      RECT MASK 2 67.883 78.03 67.943 78.3 ;
      RECT MASK 2 68.215 78.03 68.275 78.3 ;
      RECT MASK 2 68.547 78.03 68.607 78.3 ;
      RECT MASK 2 69.045 78.03 69.105 78.3 ;
      RECT MASK 2 69.377 78.03 69.437 78.3 ;
      RECT MASK 2 69.709 78.03 69.769 79.402 ;
      RECT MASK 2 71.679 78.03 71.739 78.3 ;
      RECT MASK 2 72.177 78.03 72.237 78.3 ;
      RECT MASK 2 72.509 78.03 72.569 78.3 ;
      RECT MASK 2 72.841 78.03 72.901 78.3 ;
      RECT MASK 2 73.339 78.03 73.399 78.3 ;
      RECT MASK 2 73.671 78.03 73.731 78.3 ;
      RECT MASK 2 74.003 78.03 74.063 78.3 ;
      RECT MASK 2 74.501 78.03 74.561 78.3 ;
      RECT MASK 2 74.833 78.03 74.893 78.3 ;
      RECT MASK 2 75.165 78.03 75.225 78.3 ;
      RECT MASK 2 75.663 78.03 75.723 78.3 ;
      RECT MASK 2 75.995 78.03 76.055 78.3 ;
      RECT MASK 2 76.327 78.03 76.387 79.402 ;
      RECT MASK 2 78.297 78.03 78.357 78.3 ;
      RECT MASK 2 78.795 78.03 78.855 78.3 ;
      RECT MASK 2 79.127 78.03 79.187 78.3 ;
      RECT MASK 2 79.459 78.03 79.519 78.3 ;
      RECT MASK 2 79.957 78.03 80.017 78.3 ;
      RECT MASK 2 80.289 78.03 80.349 78.3 ;
      RECT MASK 2 80.621 78.03 80.681 78.3 ;
      RECT MASK 2 81.119 78.03 81.179 78.3 ;
      RECT MASK 2 81.451 78.03 81.511 78.3 ;
      RECT MASK 2 81.783 78.03 81.843 78.3 ;
      RECT MASK 2 82.281 78.03 82.341 78.3 ;
      RECT MASK 2 82.613 78.03 82.673 78.3 ;
      RECT MASK 2 82.945 78.03 83.005 79.402 ;
      RECT MASK 2 84.915 78.03 84.975 78.3 ;
      RECT MASK 2 85.413 78.03 85.473 78.3 ;
      RECT MASK 2 85.745 78.03 85.805 78.3 ;
      RECT MASK 2 86.077 78.03 86.137 78.3 ;
      RECT MASK 2 86.575 78.03 86.635 78.3 ;
      RECT MASK 2 86.907 78.03 86.967 78.3 ;
      RECT MASK 2 87.239 78.03 87.299 78.3 ;
      RECT MASK 2 87.737 78.03 87.797 78.3 ;
      RECT MASK 2 88.069 78.03 88.129 78.3 ;
      RECT MASK 2 88.401 78.03 88.461 78.3 ;
      RECT MASK 2 88.899 78.03 88.959 78.3 ;
      RECT MASK 2 89.231 78.03 89.291 78.3 ;
      RECT MASK 2 89.563 78.03 89.623 79.402 ;
      RECT MASK 2 91.533 78.03 91.593 78.3 ;
      RECT MASK 2 92.031 78.03 92.091 78.3 ;
      RECT MASK 2 92.363 78.03 92.423 78.3 ;
      RECT MASK 2 92.695 78.03 92.755 78.3 ;
      RECT MASK 2 93.193 78.03 93.253 78.3 ;
      RECT MASK 2 93.525 78.03 93.585 78.3 ;
      RECT MASK 2 93.857 78.03 93.917 78.3 ;
      RECT MASK 2 94.355 78.03 94.415 78.3 ;
      RECT MASK 2 94.687 78.03 94.747 78.3 ;
      RECT MASK 2 95.019 78.03 95.079 78.3 ;
      RECT MASK 2 95.517 78.03 95.577 78.3 ;
      RECT MASK 2 95.849 78.03 95.909 78.3 ;
      RECT MASK 2 96.181 78.03 96.241 79.402 ;
      RECT MASK 2 98.151 78.03 98.211 78.3 ;
      RECT MASK 2 98.649 78.03 98.709 78.3 ;
      RECT MASK 2 98.981 78.03 99.041 78.3 ;
      RECT MASK 2 99.313 78.03 99.373 78.3 ;
      RECT MASK 2 99.811 78.03 99.871 78.3 ;
      RECT MASK 2 100.143 78.03 100.203 78.3 ;
      RECT MASK 2 100.475 78.03 100.535 78.3 ;
      RECT MASK 2 100.973 78.03 101.033 78.3 ;
      RECT MASK 2 101.305 78.03 101.365 78.3 ;
      RECT MASK 2 101.637 78.03 101.697 78.3 ;
      RECT MASK 2 102.135 78.03 102.195 78.3 ;
      RECT MASK 2 102.467 78.03 102.527 78.3 ;
      RECT MASK 2 102.799 78.03 102.859 79.402 ;
      RECT MASK 2 104.769 78.03 104.829 78.3 ;
      RECT MASK 2 105.267 78.03 105.327 78.3 ;
      RECT MASK 2 105.599 78.03 105.659 78.3 ;
      RECT MASK 2 105.931 78.03 105.991 78.3 ;
      RECT MASK 2 106.429 78.03 106.489 78.3 ;
      RECT MASK 2 106.761 78.03 106.821 78.3 ;
      RECT MASK 2 107.093 78.03 107.153 78.3 ;
      RECT MASK 2 107.591 78.03 107.651 78.3 ;
      RECT MASK 2 107.923 78.03 107.983 78.3 ;
      RECT MASK 2 108.255 78.03 108.315 78.3 ;
      RECT MASK 2 108.753 78.03 108.813 78.3 ;
      RECT MASK 2 109.085 78.03 109.145 78.3 ;
      RECT MASK 2 109.417 78.03 109.477 79.402 ;
      RECT MASK 2 10.883 78.0305 10.943 80.25 ;
      RECT MASK 2 11.215 78.0305 11.275 80.25 ;
      RECT MASK 2 24.119 78.0305 24.179 80.25 ;
      RECT MASK 2 24.451 78.0305 24.511 80.25 ;
      RECT MASK 2 30.737 78.0305 30.797 80.25 ;
      RECT MASK 2 31.069 78.0305 31.129 80.25 ;
      RECT MASK 2 37.355 78.0305 37.415 80.25 ;
      RECT MASK 2 37.687 78.0305 37.747 80.25 ;
      RECT MASK 2 43.973 78.0305 44.033 80.25 ;
      RECT MASK 2 44.305 78.0305 44.365 80.25 ;
      RECT MASK 2 50.591 78.0305 50.651 80.25 ;
      RECT MASK 2 50.923 78.0305 50.983 80.25 ;
      RECT MASK 2 57.209 78.0305 57.269 80.25 ;
      RECT MASK 2 57.541 78.0305 57.601 80.25 ;
      RECT MASK 2 63.827 78.0305 63.887 80.25 ;
      RECT MASK 2 64.159 78.0305 64.219 80.25 ;
      RECT MASK 2 70.445 78.0305 70.505 80.25 ;
      RECT MASK 2 70.777 78.0305 70.837 80.25 ;
      RECT MASK 2 77.063 78.0305 77.123 80.25 ;
      RECT MASK 2 77.395 78.0305 77.455 80.25 ;
      RECT MASK 2 83.681 78.0305 83.741 80.25 ;
      RECT MASK 2 84.013 78.0305 84.073 80.25 ;
      RECT MASK 2 90.299 78.0305 90.359 80.25 ;
      RECT MASK 2 90.631 78.0305 90.691 80.25 ;
      RECT MASK 2 96.917 78.0305 96.977 80.25 ;
      RECT MASK 2 97.249 78.0305 97.309 80.25 ;
      RECT MASK 2 103.535 78.0305 103.595 80.25 ;
      RECT MASK 2 103.867 78.0305 103.927 80.25 ;
      RECT MASK 2 11.951 78.033 12.011 78.7115 ;
      RECT MASK 2 16.931 78.033 16.991 78.7115 ;
      RECT MASK 2 18.569 78.033 18.629 78.7115 ;
      RECT MASK 2 23.549 78.033 23.609 78.7115 ;
      RECT MASK 2 25.187 78.033 25.247 78.7115 ;
      RECT MASK 2 30.167 78.033 30.227 78.7115 ;
      RECT MASK 2 31.805 78.033 31.865 78.7115 ;
      RECT MASK 2 36.785 78.033 36.845 78.7115 ;
      RECT MASK 2 38.423 78.033 38.483 78.7115 ;
      RECT MASK 2 43.403 78.033 43.463 78.7115 ;
      RECT MASK 2 45.041 78.033 45.101 78.7115 ;
      RECT MASK 2 50.021 78.033 50.081 78.7115 ;
      RECT MASK 2 51.659 78.033 51.719 78.7115 ;
      RECT MASK 2 56.639 78.033 56.699 78.7115 ;
      RECT MASK 2 58.277 78.033 58.337 78.7115 ;
      RECT MASK 2 63.257 78.033 63.317 78.7115 ;
      RECT MASK 2 64.895 78.033 64.955 78.7115 ;
      RECT MASK 2 69.875 78.033 69.935 78.7115 ;
      RECT MASK 2 71.513 78.033 71.573 78.7115 ;
      RECT MASK 2 76.493 78.033 76.553 78.7115 ;
      RECT MASK 2 78.131 78.033 78.191 78.7115 ;
      RECT MASK 2 83.111 78.033 83.171 78.7115 ;
      RECT MASK 2 84.749 78.033 84.809 78.7115 ;
      RECT MASK 2 89.729 78.033 89.789 78.7115 ;
      RECT MASK 2 91.367 78.033 91.427 78.7115 ;
      RECT MASK 2 96.347 78.033 96.407 78.7115 ;
      RECT MASK 2 97.985 78.033 98.045 78.7115 ;
      RECT MASK 2 102.965 78.033 103.025 78.7115 ;
      RECT MASK 2 104.603 78.033 104.663 78.7115 ;
      RECT MASK 2 109.583 78.033 109.643 78.7115 ;
      RECT MASK 2 6.817 78.586 6.897 81.8885 ;
      RECT MASK 2 7.149 78.586 7.229 81.8885 ;
      RECT MASK 2 7.481 78.586 7.561 81.8885 ;
      RECT MASK 2 7.979 78.586 8.059 81.8885 ;
      RECT MASK 2 8.311 78.586 8.391 81.8885 ;
      RECT MASK 2 8.643 78.586 8.723 81.8885 ;
      RECT MASK 2 9.141 78.586 9.221 81.8885 ;
      RECT MASK 2 9.473 78.586 9.553 81.8885 ;
      RECT MASK 2 9.805 78.586 9.885 81.8885 ;
      RECT MASK 2 12.273 78.586 12.353 81.8885 ;
      RECT MASK 2 12.605 78.586 12.685 81.8885 ;
      RECT MASK 2 12.937 78.586 13.017 81.8885 ;
      RECT MASK 2 13.435 78.586 13.515 81.8885 ;
      RECT MASK 2 13.767 78.586 13.847 81.8885 ;
      RECT MASK 2 14.099 78.586 14.179 81.8885 ;
      RECT MASK 2 14.597 78.586 14.677 81.8885 ;
      RECT MASK 2 14.929 78.586 15.009 81.8885 ;
      RECT MASK 2 15.261 78.586 15.341 81.8885 ;
      RECT MASK 2 15.759 78.586 15.839 81.8885 ;
      RECT MASK 2 16.091 78.586 16.171 81.8885 ;
      RECT MASK 2 16.423 78.586 16.503 81.8885 ;
      RECT MASK 2 18.891 78.586 18.971 81.8885 ;
      RECT MASK 2 19.223 78.586 19.303 81.8885 ;
      RECT MASK 2 19.555 78.586 19.635 81.8885 ;
      RECT MASK 2 20.053 78.586 20.133 81.8885 ;
      RECT MASK 2 20.385 78.586 20.465 81.8885 ;
      RECT MASK 2 20.717 78.586 20.797 81.8885 ;
      RECT MASK 2 21.215 78.586 21.295 81.8885 ;
      RECT MASK 2 21.547 78.586 21.627 81.8885 ;
      RECT MASK 2 21.879 78.586 21.959 81.8885 ;
      RECT MASK 2 22.377 78.586 22.457 81.8885 ;
      RECT MASK 2 22.709 78.586 22.789 81.8885 ;
      RECT MASK 2 23.041 78.586 23.121 81.8885 ;
      RECT MASK 2 25.509 78.586 25.589 81.8885 ;
      RECT MASK 2 25.841 78.586 25.921 81.8885 ;
      RECT MASK 2 26.173 78.586 26.253 81.8885 ;
      RECT MASK 2 26.671 78.586 26.751 81.8885 ;
      RECT MASK 2 27.003 78.586 27.083 81.8885 ;
      RECT MASK 2 27.335 78.586 27.415 81.8885 ;
      RECT MASK 2 27.833 78.586 27.913 81.8885 ;
      RECT MASK 2 28.165 78.586 28.245 81.8885 ;
      RECT MASK 2 28.497 78.586 28.577 81.8885 ;
      RECT MASK 2 28.995 78.586 29.075 81.8885 ;
      RECT MASK 2 29.327 78.586 29.407 81.8885 ;
      RECT MASK 2 29.659 78.586 29.739 81.8885 ;
      RECT MASK 2 32.127 78.586 32.207 81.8885 ;
      RECT MASK 2 32.459 78.586 32.539 81.8885 ;
      RECT MASK 2 32.791 78.586 32.871 81.8885 ;
      RECT MASK 2 33.289 78.586 33.369 81.8885 ;
      RECT MASK 2 33.621 78.586 33.701 81.8885 ;
      RECT MASK 2 33.953 78.586 34.033 81.8885 ;
      RECT MASK 2 34.451 78.586 34.531 81.8885 ;
      RECT MASK 2 34.783 78.586 34.863 81.8885 ;
      RECT MASK 2 35.115 78.586 35.195 81.8885 ;
      RECT MASK 2 35.613 78.586 35.693 81.8885 ;
      RECT MASK 2 35.945 78.586 36.025 81.8885 ;
      RECT MASK 2 36.277 78.586 36.357 81.8885 ;
      RECT MASK 2 38.745 78.586 38.825 81.8885 ;
      RECT MASK 2 39.077 78.586 39.157 81.8885 ;
      RECT MASK 2 39.409 78.586 39.489 81.8885 ;
      RECT MASK 2 39.907 78.586 39.987 81.8885 ;
      RECT MASK 2 40.239 78.586 40.319 81.8885 ;
      RECT MASK 2 40.571 78.586 40.651 81.8885 ;
      RECT MASK 2 41.069 78.586 41.149 81.8885 ;
      RECT MASK 2 41.401 78.586 41.481 81.8885 ;
      RECT MASK 2 41.733 78.586 41.813 81.8885 ;
      RECT MASK 2 42.231 78.586 42.311 81.8885 ;
      RECT MASK 2 42.563 78.586 42.643 81.8885 ;
      RECT MASK 2 42.895 78.586 42.975 81.8885 ;
      RECT MASK 2 45.363 78.586 45.443 81.8885 ;
      RECT MASK 2 45.695 78.586 45.775 81.8885 ;
      RECT MASK 2 46.027 78.586 46.107 81.8885 ;
      RECT MASK 2 46.525 78.586 46.605 81.8885 ;
      RECT MASK 2 46.857 78.586 46.937 81.8885 ;
      RECT MASK 2 47.189 78.586 47.269 81.8885 ;
      RECT MASK 2 47.687 78.586 47.767 81.8885 ;
      RECT MASK 2 48.019 78.586 48.099 81.8885 ;
      RECT MASK 2 48.351 78.586 48.431 81.8885 ;
      RECT MASK 2 48.849 78.586 48.929 81.8885 ;
      RECT MASK 2 49.181 78.586 49.261 81.8885 ;
      RECT MASK 2 49.513 78.586 49.593 81.8885 ;
      RECT MASK 2 51.981 78.586 52.061 81.8885 ;
      RECT MASK 2 52.313 78.586 52.393 81.8885 ;
      RECT MASK 2 52.645 78.586 52.725 81.8885 ;
      RECT MASK 2 53.143 78.586 53.223 81.8885 ;
      RECT MASK 2 53.475 78.586 53.555 81.8885 ;
      RECT MASK 2 53.807 78.586 53.887 81.8885 ;
      RECT MASK 2 54.305 78.586 54.385 81.8885 ;
      RECT MASK 2 54.637 78.586 54.717 81.8885 ;
      RECT MASK 2 54.969 78.586 55.049 81.8885 ;
      RECT MASK 2 55.467 78.586 55.547 81.8885 ;
      RECT MASK 2 55.799 78.586 55.879 81.8885 ;
      RECT MASK 2 56.131 78.586 56.211 81.8885 ;
      RECT MASK 2 58.599 78.586 58.679 81.8885 ;
      RECT MASK 2 58.931 78.586 59.011 81.8885 ;
      RECT MASK 2 59.263 78.586 59.343 81.8885 ;
      RECT MASK 2 59.761 78.586 59.841 81.8885 ;
      RECT MASK 2 60.093 78.586 60.173 81.8885 ;
      RECT MASK 2 60.425 78.586 60.505 81.8885 ;
      RECT MASK 2 60.923 78.586 61.003 81.8885 ;
      RECT MASK 2 61.255 78.586 61.335 81.8885 ;
      RECT MASK 2 61.587 78.586 61.667 81.8885 ;
      RECT MASK 2 62.085 78.586 62.165 81.8885 ;
      RECT MASK 2 62.417 78.586 62.497 81.8885 ;
      RECT MASK 2 62.749 78.586 62.829 81.8885 ;
      RECT MASK 2 65.217 78.586 65.297 81.8885 ;
      RECT MASK 2 65.549 78.586 65.629 81.8885 ;
      RECT MASK 2 65.881 78.586 65.961 81.8885 ;
      RECT MASK 2 66.379 78.586 66.459 81.8885 ;
      RECT MASK 2 66.711 78.586 66.791 81.8885 ;
      RECT MASK 2 67.043 78.586 67.123 81.8885 ;
      RECT MASK 2 67.541 78.586 67.621 81.8885 ;
      RECT MASK 2 67.873 78.586 67.953 81.8885 ;
      RECT MASK 2 68.205 78.586 68.285 81.8885 ;
      RECT MASK 2 68.703 78.586 68.783 81.8885 ;
      RECT MASK 2 69.035 78.586 69.115 81.8885 ;
      RECT MASK 2 69.367 78.586 69.447 81.8885 ;
      RECT MASK 2 71.835 78.586 71.915 81.8885 ;
      RECT MASK 2 72.167 78.586 72.247 81.8885 ;
      RECT MASK 2 72.499 78.586 72.579 81.8885 ;
      RECT MASK 2 72.997 78.586 73.077 81.8885 ;
      RECT MASK 2 73.329 78.586 73.409 81.8885 ;
      RECT MASK 2 73.661 78.586 73.741 81.8885 ;
      RECT MASK 2 74.159 78.586 74.239 81.8885 ;
      RECT MASK 2 74.491 78.586 74.571 81.8885 ;
      RECT MASK 2 74.823 78.586 74.903 81.8885 ;
      RECT MASK 2 75.321 78.586 75.401 81.8885 ;
      RECT MASK 2 75.653 78.586 75.733 81.8885 ;
      RECT MASK 2 75.985 78.586 76.065 81.8885 ;
      RECT MASK 2 78.453 78.586 78.533 81.8885 ;
      RECT MASK 2 78.785 78.586 78.865 81.8885 ;
      RECT MASK 2 79.117 78.586 79.197 81.8885 ;
      RECT MASK 2 79.615 78.586 79.695 81.8885 ;
      RECT MASK 2 79.947 78.586 80.027 81.8885 ;
      RECT MASK 2 80.279 78.586 80.359 81.8885 ;
      RECT MASK 2 80.777 78.586 80.857 81.8885 ;
      RECT MASK 2 81.109 78.586 81.189 81.8885 ;
      RECT MASK 2 81.441 78.586 81.521 81.8885 ;
      RECT MASK 2 81.939 78.586 82.019 81.8885 ;
      RECT MASK 2 82.271 78.586 82.351 81.8885 ;
      RECT MASK 2 82.603 78.586 82.683 81.8885 ;
      RECT MASK 2 85.071 78.586 85.151 81.8885 ;
      RECT MASK 2 85.403 78.586 85.483 81.8885 ;
      RECT MASK 2 85.735 78.586 85.815 81.8885 ;
      RECT MASK 2 86.233 78.586 86.313 81.8885 ;
      RECT MASK 2 86.565 78.586 86.645 81.8885 ;
      RECT MASK 2 86.897 78.586 86.977 81.8885 ;
      RECT MASK 2 87.395 78.586 87.475 81.8885 ;
      RECT MASK 2 87.727 78.586 87.807 81.8885 ;
      RECT MASK 2 88.059 78.586 88.139 81.8885 ;
      RECT MASK 2 88.557 78.586 88.637 81.8885 ;
      RECT MASK 2 88.889 78.586 88.969 81.8885 ;
      RECT MASK 2 89.221 78.586 89.301 81.8885 ;
      RECT MASK 2 91.689 78.586 91.769 81.8885 ;
      RECT MASK 2 92.021 78.586 92.101 81.8885 ;
      RECT MASK 2 92.353 78.586 92.433 81.8885 ;
      RECT MASK 2 92.851 78.586 92.931 81.8885 ;
      RECT MASK 2 93.183 78.586 93.263 81.8885 ;
      RECT MASK 2 93.515 78.586 93.595 81.8885 ;
      RECT MASK 2 94.013 78.586 94.093 81.8885 ;
      RECT MASK 2 94.345 78.586 94.425 81.8885 ;
      RECT MASK 2 94.677 78.586 94.757 81.8885 ;
      RECT MASK 2 95.175 78.586 95.255 81.8885 ;
      RECT MASK 2 95.507 78.586 95.587 81.8885 ;
      RECT MASK 2 95.839 78.586 95.919 81.8885 ;
      RECT MASK 2 98.307 78.586 98.387 81.8885 ;
      RECT MASK 2 98.639 78.586 98.719 81.8885 ;
      RECT MASK 2 98.971 78.586 99.051 81.8885 ;
      RECT MASK 2 99.469 78.586 99.549 81.8885 ;
      RECT MASK 2 99.801 78.586 99.881 81.8885 ;
      RECT MASK 2 100.133 78.586 100.213 81.8885 ;
      RECT MASK 2 100.631 78.586 100.711 81.8885 ;
      RECT MASK 2 100.963 78.586 101.043 81.8885 ;
      RECT MASK 2 101.295 78.586 101.375 81.8885 ;
      RECT MASK 2 101.793 78.586 101.873 81.8885 ;
      RECT MASK 2 102.125 78.586 102.205 81.8885 ;
      RECT MASK 2 102.457 78.586 102.537 81.8885 ;
      RECT MASK 2 104.925 78.586 105.005 81.8885 ;
      RECT MASK 2 105.257 78.586 105.337 81.8885 ;
      RECT MASK 2 105.589 78.586 105.669 81.8885 ;
      RECT MASK 2 106.087 78.586 106.167 81.8885 ;
      RECT MASK 2 106.419 78.586 106.499 81.8885 ;
      RECT MASK 2 106.751 78.586 106.831 81.8885 ;
      RECT MASK 2 107.249 78.586 107.329 81.8885 ;
      RECT MASK 2 107.581 78.586 107.661 81.8885 ;
      RECT MASK 2 107.913 78.586 107.993 81.8885 ;
      RECT MASK 2 108.411 78.586 108.491 81.8885 ;
      RECT MASK 2 108.743 78.586 108.823 81.8885 ;
      RECT MASK 2 109.075 78.586 109.155 81.8885 ;
      RECT MASK 2 111.377 78.785 111.437 79.045 ;
      RECT MASK 2 111.709 78.785 111.769 79.045 ;
      RECT MASK 2 112.041 78.785 112.101 79.045 ;
      RECT MASK 2 112.373 78.785 112.433 79.045 ;
      RECT MASK 2 112.705 78.785 112.765 79.045 ;
      RECT MASK 2 113.037 78.785 113.097 79.045 ;
      RECT MASK 2 2.204 79.05 2.264 95.88 ;
      RECT MASK 2 2.478 79.05 2.538 95.88 ;
      RECT MASK 2 2.752 79.05 2.812 95.88 ;
      RECT MASK 2 3.026 79.05 3.086 95.88 ;
      RECT MASK 2 3.3 79.05 3.36 95.88 ;
      RECT MASK 2 3.574 79.05 3.634 95.88 ;
      RECT MASK 2 3.848 79.05 3.908 95.88 ;
      RECT MASK 2 4.122 79.05 4.182 95.88 ;
      RECT MASK 2 4.396 79.05 4.456 95.88 ;
      RECT MASK 2 111.792 79.211 111.852 81.511 ;
      RECT MASK 2 104.2115 79.661 104.2715 85.604 ;
      RECT MASK 2 112.622 79.679 112.682 81.979 ;
      RECT MASK 2 6.661 79.98 6.721 80.25 ;
      RECT MASK 2 7.823 79.98 7.883 80.25 ;
      RECT MASK 2 8.985 79.98 9.045 80.25 ;
      RECT MASK 2 10.147 79.98 10.207 80.25 ;
      RECT MASK 2 12.117 79.98 12.177 80.25 ;
      RECT MASK 2 13.279 79.98 13.339 80.25 ;
      RECT MASK 2 14.441 79.98 14.501 80.25 ;
      RECT MASK 2 15.603 79.98 15.663 80.25 ;
      RECT MASK 2 16.765 79.98 16.825 80.25 ;
      RECT MASK 2 18.735 79.98 18.795 80.25 ;
      RECT MASK 2 19.897 79.98 19.957 80.25 ;
      RECT MASK 2 21.059 79.98 21.119 80.25 ;
      RECT MASK 2 22.221 79.98 22.281 80.25 ;
      RECT MASK 2 23.383 79.98 23.443 80.25 ;
      RECT MASK 2 25.353 79.98 25.413 80.25 ;
      RECT MASK 2 26.515 79.98 26.575 80.25 ;
      RECT MASK 2 27.677 79.98 27.737 80.25 ;
      RECT MASK 2 28.839 79.98 28.899 80.25 ;
      RECT MASK 2 30.001 79.98 30.061 80.25 ;
      RECT MASK 2 31.971 79.98 32.031 80.25 ;
      RECT MASK 2 33.133 79.98 33.193 80.25 ;
      RECT MASK 2 34.295 79.98 34.355 80.25 ;
      RECT MASK 2 35.457 79.98 35.517 80.25 ;
      RECT MASK 2 36.619 79.98 36.679 80.25 ;
      RECT MASK 2 38.589 79.98 38.649 80.25 ;
      RECT MASK 2 39.751 79.98 39.811 80.25 ;
      RECT MASK 2 40.913 79.98 40.973 80.25 ;
      RECT MASK 2 42.075 79.98 42.135 80.25 ;
      RECT MASK 2 43.237 79.98 43.297 80.25 ;
      RECT MASK 2 45.207 79.98 45.267 80.25 ;
      RECT MASK 2 46.369 79.98 46.429 80.25 ;
      RECT MASK 2 47.531 79.98 47.591 80.25 ;
      RECT MASK 2 48.693 79.98 48.753 80.25 ;
      RECT MASK 2 49.855 79.98 49.915 80.25 ;
      RECT MASK 2 51.825 79.98 51.885 80.25 ;
      RECT MASK 2 52.987 79.98 53.047 80.25 ;
      RECT MASK 2 54.149 79.98 54.209 80.25 ;
      RECT MASK 2 55.311 79.98 55.371 80.25 ;
      RECT MASK 2 56.473 79.98 56.533 80.25 ;
      RECT MASK 2 58.443 79.98 58.503 80.25 ;
      RECT MASK 2 59.605 79.98 59.665 80.25 ;
      RECT MASK 2 60.767 79.98 60.827 80.25 ;
      RECT MASK 2 61.929 79.98 61.989 80.25 ;
      RECT MASK 2 63.091 79.98 63.151 80.25 ;
      RECT MASK 2 65.061 79.98 65.121 80.25 ;
      RECT MASK 2 66.223 79.98 66.283 80.25 ;
      RECT MASK 2 67.385 79.98 67.445 80.25 ;
      RECT MASK 2 68.547 79.98 68.607 80.25 ;
      RECT MASK 2 69.709 79.98 69.769 80.25 ;
      RECT MASK 2 71.679 79.98 71.739 80.25 ;
      RECT MASK 2 72.841 79.98 72.901 80.25 ;
      RECT MASK 2 74.003 79.98 74.063 80.25 ;
      RECT MASK 2 75.165 79.98 75.225 80.25 ;
      RECT MASK 2 76.327 79.98 76.387 80.25 ;
      RECT MASK 2 78.297 79.98 78.357 80.25 ;
      RECT MASK 2 79.459 79.98 79.519 80.25 ;
      RECT MASK 2 80.621 79.98 80.681 80.25 ;
      RECT MASK 2 81.783 79.98 81.843 80.25 ;
      RECT MASK 2 82.945 79.98 83.005 80.25 ;
      RECT MASK 2 84.915 79.98 84.975 80.25 ;
      RECT MASK 2 86.077 79.98 86.137 80.25 ;
      RECT MASK 2 87.239 79.98 87.299 80.25 ;
      RECT MASK 2 88.401 79.98 88.461 80.25 ;
      RECT MASK 2 89.563 79.98 89.623 80.25 ;
      RECT MASK 2 91.533 79.98 91.593 80.25 ;
      RECT MASK 2 92.695 79.98 92.755 80.25 ;
      RECT MASK 2 93.857 79.98 93.917 80.25 ;
      RECT MASK 2 95.019 79.98 95.079 80.25 ;
      RECT MASK 2 96.181 79.98 96.241 80.25 ;
      RECT MASK 2 98.151 79.98 98.211 80.25 ;
      RECT MASK 2 99.313 79.98 99.373 80.25 ;
      RECT MASK 2 100.475 79.98 100.535 80.25 ;
      RECT MASK 2 101.637 79.98 101.697 80.25 ;
      RECT MASK 2 102.799 79.98 102.859 80.25 ;
      RECT MASK 2 104.769 79.98 104.829 80.25 ;
      RECT MASK 2 105.931 79.98 105.991 80.25 ;
      RECT MASK 2 107.093 79.98 107.153 80.25 ;
      RECT MASK 2 108.255 79.98 108.315 80.25 ;
      RECT MASK 2 109.417 79.98 109.477 80.25 ;
      RECT MASK 2 116.427 80.126 116.507 80.458 ;
      RECT MASK 2 116.759 80.126 116.839 80.458 ;
      RECT MASK 2 117.091 80.126 117.171 80.458 ;
      RECT MASK 2 117.423 80.126 117.503 80.458 ;
      RECT MASK 2 117.755 80.126 117.835 80.458 ;
      RECT MASK 2 118.087 80.126 118.167 80.458 ;
      RECT MASK 2 118.419 80.126 118.499 80.458 ;
      RECT MASK 2 118.751 80.126 118.831 80.458 ;
      RECT MASK 2 119.083 80.126 119.163 80.458 ;
      RECT MASK 2 119.415 80.126 119.495 80.458 ;
      RECT MASK 2 119.747 80.126 119.827 80.458 ;
      RECT MASK 2 120.079 80.126 120.159 80.458 ;
      RECT MASK 2 120.411 80.126 120.491 80.458 ;
      RECT MASK 2 120.743 80.126 120.823 80.458 ;
      RECT MASK 2 121.075 80.126 121.155 80.458 ;
      RECT MASK 2 121.407 80.126 121.487 80.458 ;
      RECT MASK 2 121.739 80.126 121.819 80.458 ;
      RECT MASK 2 122.071 80.126 122.151 80.458 ;
      RECT MASK 2 122.403 80.126 122.483 80.458 ;
      RECT MASK 2 122.735 80.126 122.815 80.458 ;
      RECT MASK 2 123.067 80.126 123.147 80.458 ;
      RECT MASK 2 123.399 80.126 123.479 80.458 ;
      RECT MASK 2 123.731 80.126 123.811 80.458 ;
      RECT MASK 2 124.063 80.126 124.143 80.458 ;
      RECT MASK 2 124.395 80.126 124.475 80.458 ;
      RECT MASK 2 124.727 80.126 124.807 80.458 ;
      RECT MASK 2 125.059 80.126 125.139 80.458 ;
      RECT MASK 2 125.391 80.126 125.471 80.458 ;
      RECT MASK 2 125.723 80.126 125.803 80.458 ;
      RECT MASK 2 126.055 80.126 126.135 80.458 ;
      RECT MASK 2 6.661 80.43 6.721 80.7 ;
      RECT MASK 2 7.823 80.43 7.883 80.7 ;
      RECT MASK 2 8.985 80.43 9.045 80.7 ;
      RECT MASK 2 10.147 80.43 10.207 80.7 ;
      RECT MASK 2 12.117 80.43 12.177 80.7 ;
      RECT MASK 2 13.279 80.43 13.339 80.7 ;
      RECT MASK 2 14.441 80.43 14.501 80.7 ;
      RECT MASK 2 15.603 80.43 15.663 80.7 ;
      RECT MASK 2 16.765 80.43 16.825 80.7 ;
      RECT MASK 2 18.735 80.43 18.795 80.7 ;
      RECT MASK 2 19.897 80.43 19.957 80.7 ;
      RECT MASK 2 21.059 80.43 21.119 80.7 ;
      RECT MASK 2 22.221 80.43 22.281 80.7 ;
      RECT MASK 2 23.383 80.43 23.443 80.7 ;
      RECT MASK 2 25.353 80.43 25.413 80.7 ;
      RECT MASK 2 26.515 80.43 26.575 80.7 ;
      RECT MASK 2 27.677 80.43 27.737 80.7 ;
      RECT MASK 2 28.839 80.43 28.899 80.7 ;
      RECT MASK 2 30.001 80.43 30.061 80.7 ;
      RECT MASK 2 31.971 80.43 32.031 80.7 ;
      RECT MASK 2 33.133 80.43 33.193 80.7 ;
      RECT MASK 2 34.295 80.43 34.355 80.7 ;
      RECT MASK 2 35.457 80.43 35.517 80.7 ;
      RECT MASK 2 36.619 80.43 36.679 80.7 ;
      RECT MASK 2 38.589 80.43 38.649 80.7 ;
      RECT MASK 2 39.751 80.43 39.811 80.7 ;
      RECT MASK 2 40.913 80.43 40.973 80.7 ;
      RECT MASK 2 42.075 80.43 42.135 80.7 ;
      RECT MASK 2 43.237 80.43 43.297 80.7 ;
      RECT MASK 2 45.207 80.43 45.267 80.7 ;
      RECT MASK 2 46.369 80.43 46.429 80.7 ;
      RECT MASK 2 47.531 80.43 47.591 80.7 ;
      RECT MASK 2 48.693 80.43 48.753 80.7 ;
      RECT MASK 2 49.855 80.43 49.915 80.7 ;
      RECT MASK 2 51.825 80.43 51.885 80.7 ;
      RECT MASK 2 52.987 80.43 53.047 80.7 ;
      RECT MASK 2 54.149 80.43 54.209 80.7 ;
      RECT MASK 2 55.311 80.43 55.371 80.7 ;
      RECT MASK 2 56.473 80.43 56.533 80.7 ;
      RECT MASK 2 58.443 80.43 58.503 84.169 ;
      RECT MASK 2 59.605 80.43 59.665 84.157 ;
      RECT MASK 2 60.767 80.43 60.827 80.7 ;
      RECT MASK 2 61.929 80.43 61.989 80.7 ;
      RECT MASK 2 63.091 80.43 63.151 80.7 ;
      RECT MASK 2 63.544 80.43 63.694 84.157 ;
      RECT MASK 2 65.061 80.43 65.121 80.7 ;
      RECT MASK 2 66.223 80.43 66.283 80.7 ;
      RECT MASK 2 67.385 80.43 67.445 80.7 ;
      RECT MASK 2 68.547 80.43 68.607 80.7 ;
      RECT MASK 2 69.709 80.43 69.769 80.7 ;
      RECT MASK 2 71.679 80.43 71.739 80.7 ;
      RECT MASK 2 72.841 80.43 72.901 80.7 ;
      RECT MASK 2 74.003 80.43 74.063 80.7 ;
      RECT MASK 2 75.165 80.43 75.225 80.7 ;
      RECT MASK 2 76.327 80.43 76.387 80.7 ;
      RECT MASK 2 78.297 80.43 78.357 80.7 ;
      RECT MASK 2 79.459 80.43 79.519 80.7 ;
      RECT MASK 2 80.621 80.43 80.681 80.7 ;
      RECT MASK 2 81.783 80.43 81.843 80.7 ;
      RECT MASK 2 82.945 80.43 83.005 80.7 ;
      RECT MASK 2 84.915 80.43 84.975 80.7 ;
      RECT MASK 2 86.077 80.43 86.137 80.7 ;
      RECT MASK 2 87.239 80.43 87.299 80.7 ;
      RECT MASK 2 88.401 80.43 88.461 80.7 ;
      RECT MASK 2 89.563 80.43 89.623 80.7 ;
      RECT MASK 2 91.533 80.43 91.593 80.7 ;
      RECT MASK 2 92.695 80.43 92.755 80.7 ;
      RECT MASK 2 93.857 80.43 93.917 80.7 ;
      RECT MASK 2 95.019 80.43 95.079 80.7 ;
      RECT MASK 2 96.181 80.43 96.241 80.7 ;
      RECT MASK 2 98.151 80.43 98.211 80.7 ;
      RECT MASK 2 99.313 80.43 99.373 80.7 ;
      RECT MASK 2 100.475 80.43 100.535 80.7 ;
      RECT MASK 2 101.637 80.43 101.697 80.7 ;
      RECT MASK 2 102.799 80.43 102.859 80.7 ;
      RECT MASK 2 104.769 80.43 104.829 80.7 ;
      RECT MASK 2 105.931 80.43 105.991 80.7 ;
      RECT MASK 2 107.093 80.43 107.153 80.7 ;
      RECT MASK 2 108.255 80.43 108.315 80.7 ;
      RECT MASK 2 109.417 80.43 109.477 80.7 ;
      RECT MASK 2 18.403 80.4335 18.463 82.645 ;
      RECT MASK 2 23.715 80.4335 23.775 82.645 ;
      RECT MASK 2 25.021 80.4335 25.081 82.645 ;
      RECT MASK 2 30.333 80.4335 30.393 82.645 ;
      RECT MASK 2 31.639 80.4335 31.699 82.645 ;
      RECT MASK 2 36.951 80.4335 37.011 82.645 ;
      RECT MASK 2 38.257 80.4335 38.317 82.645 ;
      RECT MASK 2 43.569 80.4335 43.629 82.645 ;
      RECT MASK 2 44.875 80.4335 44.935 82.645 ;
      RECT MASK 2 50.187 80.4335 50.247 82.645 ;
      RECT MASK 2 51.493 80.4335 51.553 82.645 ;
      RECT MASK 2 56.805 80.4335 56.865 82.645 ;
      RECT MASK 2 57.9 80.4335 58.05 84.157 ;
      RECT MASK 2 64.729 80.4335 64.789 82.645 ;
      RECT MASK 2 70.041 80.4335 70.101 82.645 ;
      RECT MASK 2 71.347 80.4335 71.407 82.645 ;
      RECT MASK 2 76.659 80.4335 76.719 82.645 ;
      RECT MASK 2 77.965 80.4335 78.025 82.645 ;
      RECT MASK 2 83.277 80.4335 83.337 82.645 ;
      RECT MASK 2 84.583 80.4335 84.643 82.645 ;
      RECT MASK 2 89.895 80.4335 89.955 82.645 ;
      RECT MASK 2 91.201 80.4335 91.261 82.645 ;
      RECT MASK 2 96.513 80.4335 96.573 82.645 ;
      RECT MASK 2 97.819 80.4335 97.879 82.645 ;
      RECT MASK 2 104.437 80.4335 104.497 82.645 ;
      RECT MASK 2 10.883 80.4655 10.943 84.157 ;
      RECT MASK 2 11.215 80.4655 11.275 84.157 ;
      RECT MASK 2 17.501 80.4655 17.561 84.157 ;
      RECT MASK 2 17.833 80.4655 17.893 84.157 ;
      RECT MASK 2 24.119 80.4655 24.179 84.157 ;
      RECT MASK 2 24.451 80.4655 24.511 84.157 ;
      RECT MASK 2 30.737 80.4655 30.797 84.157 ;
      RECT MASK 2 31.069 80.4655 31.129 84.157 ;
      RECT MASK 2 37.355 80.4655 37.415 84.157 ;
      RECT MASK 2 37.687 80.4655 37.747 84.157 ;
      RECT MASK 2 43.973 80.4655 44.033 84.157 ;
      RECT MASK 2 44.305 80.4655 44.365 84.157 ;
      RECT MASK 2 50.591 80.4655 50.651 84.157 ;
      RECT MASK 2 50.923 80.4655 50.983 84.157 ;
      RECT MASK 2 57.209 80.4655 57.269 84.157 ;
      RECT MASK 2 57.541 80.4655 57.601 84.157 ;
      RECT MASK 2 63.827 80.4655 63.887 84.157 ;
      RECT MASK 2 64.159 80.4655 64.219 84.157 ;
      RECT MASK 2 70.445 80.4655 70.505 84.157 ;
      RECT MASK 2 70.777 80.4655 70.837 84.157 ;
      RECT MASK 2 77.063 80.4655 77.123 84.157 ;
      RECT MASK 2 77.395 80.4655 77.455 84.157 ;
      RECT MASK 2 83.681 80.4655 83.741 84.157 ;
      RECT MASK 2 84.013 80.4655 84.073 84.157 ;
      RECT MASK 2 90.299 80.4655 90.359 84.157 ;
      RECT MASK 2 90.631 80.4655 90.691 84.157 ;
      RECT MASK 2 96.917 80.4655 96.977 84.157 ;
      RECT MASK 2 97.249 80.4655 97.309 84.157 ;
      RECT MASK 2 103.535 80.4655 103.595 84.157 ;
      RECT MASK 2 103.867 80.4655 103.927 84.157 ;
      RECT MASK 2 111.792 81.631 111.852 81.925 ;
      RECT MASK 2 116.599 81.84 116.659 96.66 ;
      RECT MASK 2 116.873 81.84 116.933 96.66 ;
      RECT MASK 2 117.147 81.84 117.207 96.66 ;
      RECT MASK 2 117.421 81.84 117.481 96.66 ;
      RECT MASK 2 117.695 81.84 117.755 96.66 ;
      RECT MASK 2 117.969 81.84 118.029 96.66 ;
      RECT MASK 2 118.243 81.84 118.303 96.66 ;
      RECT MASK 2 118.517 81.84 118.577 96.66 ;
      RECT MASK 2 118.791 81.84 118.851 96.66 ;
      RECT MASK 2 119.065 81.84 119.125 96.66 ;
      RECT MASK 2 119.339 81.84 119.399 96.66 ;
      RECT MASK 2 119.613 81.84 119.673 96.66 ;
      RECT MASK 2 119.887 81.84 119.947 96.66 ;
      RECT MASK 2 120.161 81.84 120.221 96.66 ;
      RECT MASK 2 120.435 81.84 120.495 96.66 ;
      RECT MASK 2 120.709 81.84 120.769 96.66 ;
      RECT MASK 2 120.983 81.84 121.043 96.66 ;
      RECT MASK 2 121.257 81.84 121.317 96.66 ;
      RECT MASK 2 121.531 81.84 121.591 96.66 ;
      RECT MASK 2 121.805 81.84 121.865 96.66 ;
      RECT MASK 2 122.079 81.84 122.139 96.66 ;
      RECT MASK 2 122.353 81.84 122.413 96.66 ;
      RECT MASK 2 122.627 81.84 122.687 96.66 ;
      RECT MASK 2 122.901 81.84 122.961 96.66 ;
      RECT MASK 2 123.175 81.84 123.235 96.66 ;
      RECT MASK 2 123.449 81.84 123.509 96.66 ;
      RECT MASK 2 123.723 81.84 123.783 96.66 ;
      RECT MASK 2 123.997 81.84 124.057 96.66 ;
      RECT MASK 2 124.271 81.84 124.331 96.66 ;
      RECT MASK 2 124.545 81.84 124.605 96.66 ;
      RECT MASK 2 124.819 81.84 124.879 96.66 ;
      RECT MASK 2 125.093 81.84 125.153 96.66 ;
      RECT MASK 2 125.367 81.84 125.427 96.66 ;
      RECT MASK 2 125.641 81.84 125.701 96.66 ;
      RECT MASK 2 125.915 81.84 125.975 96.66 ;
      RECT MASK 2 126.189 81.84 126.249 96.66 ;
      RECT MASK 2 126.463 81.84 126.523 96.66 ;
      RECT MASK 2 126.737 81.84 126.797 96.66 ;
      RECT MASK 2 127.011 81.84 127.071 96.66 ;
      RECT MASK 2 127.285 81.84 127.345 96.66 ;
      RECT MASK 2 127.559 81.84 127.619 96.66 ;
      RECT MASK 2 63.046 81.893 63.196 84.157 ;
      RECT MASK 2 58.734 82.013 58.774 82.675 ;
      RECT MASK 2 59.896 82.013 59.936 82.675 ;
      RECT MASK 2 60.722 82.013 60.872 84.157 ;
      RECT MASK 2 61.058 82.013 61.098 82.675 ;
      RECT MASK 2 61.884 82.013 62.034 84.157 ;
      RECT MASK 2 62.22 82.013 62.26 82.675 ;
      RECT MASK 2 7.076 82.0405 7.136 85.241 ;
      RECT MASK 2 8.238 82.0405 8.298 85.241 ;
      RECT MASK 2 9.4 82.0405 9.46 85.241 ;
      RECT MASK 2 12.532 82.0405 12.592 85.241 ;
      RECT MASK 2 13.694 82.0405 13.754 85.241 ;
      RECT MASK 2 14.856 82.0405 14.916 85.241 ;
      RECT MASK 2 16.018 82.0405 16.078 85.241 ;
      RECT MASK 2 19.15 82.0405 19.21 85.241 ;
      RECT MASK 2 20.312 82.0405 20.372 85.241 ;
      RECT MASK 2 21.474 82.0405 21.534 85.241 ;
      RECT MASK 2 22.636 82.0405 22.696 85.241 ;
      RECT MASK 2 25.768 82.0405 25.828 85.241 ;
      RECT MASK 2 26.93 82.0405 26.99 85.241 ;
      RECT MASK 2 28.092 82.0405 28.152 85.241 ;
      RECT MASK 2 29.254 82.0405 29.314 85.241 ;
      RECT MASK 2 32.386 82.0405 32.446 85.241 ;
      RECT MASK 2 33.548 82.0405 33.608 85.241 ;
      RECT MASK 2 34.71 82.0405 34.77 85.241 ;
      RECT MASK 2 35.872 82.0405 35.932 85.241 ;
      RECT MASK 2 39.004 82.0405 39.064 85.241 ;
      RECT MASK 2 40.166 82.0405 40.226 85.241 ;
      RECT MASK 2 41.328 82.0405 41.388 85.241 ;
      RECT MASK 2 42.49 82.0405 42.55 85.241 ;
      RECT MASK 2 45.622 82.0405 45.682 85.241 ;
      RECT MASK 2 46.784 82.0405 46.844 85.241 ;
      RECT MASK 2 47.946 82.0405 48.006 85.241 ;
      RECT MASK 2 49.108 82.0405 49.168 85.241 ;
      RECT MASK 2 52.24 82.0405 52.3 85.241 ;
      RECT MASK 2 53.402 82.0405 53.462 85.241 ;
      RECT MASK 2 54.564 82.0405 54.624 85.241 ;
      RECT MASK 2 55.726 82.0405 55.786 85.241 ;
      RECT MASK 2 58.858 82.0405 58.918 85.241 ;
      RECT MASK 2 60.02 82.0405 60.08 85.241 ;
      RECT MASK 2 61.182 82.0405 61.242 85.241 ;
      RECT MASK 2 62.344 82.0405 62.404 85.241 ;
      RECT MASK 2 65.476 82.0405 65.536 85.241 ;
      RECT MASK 2 66.638 82.0405 66.698 85.241 ;
      RECT MASK 2 67.8 82.0405 67.86 85.241 ;
      RECT MASK 2 68.962 82.0405 69.022 85.241 ;
      RECT MASK 2 72.094 82.0405 72.154 85.241 ;
      RECT MASK 2 73.256 82.0405 73.316 85.241 ;
      RECT MASK 2 74.418 82.0405 74.478 85.241 ;
      RECT MASK 2 75.58 82.0405 75.64 85.241 ;
      RECT MASK 2 78.712 82.0405 78.772 85.241 ;
      RECT MASK 2 79.874 82.0405 79.934 85.241 ;
      RECT MASK 2 81.036 82.0405 81.096 85.241 ;
      RECT MASK 2 82.198 82.0405 82.258 85.241 ;
      RECT MASK 2 85.33 82.0405 85.39 85.241 ;
      RECT MASK 2 86.492 82.0405 86.552 85.241 ;
      RECT MASK 2 87.654 82.0405 87.714 85.241 ;
      RECT MASK 2 88.816 82.0405 88.876 85.241 ;
      RECT MASK 2 91.948 82.0405 92.008 85.241 ;
      RECT MASK 2 93.11 82.0405 93.17 85.241 ;
      RECT MASK 2 94.272 82.0405 94.332 85.241 ;
      RECT MASK 2 95.434 82.0405 95.494 85.241 ;
      RECT MASK 2 98.566 82.0405 98.626 85.241 ;
      RECT MASK 2 99.728 82.0405 99.788 85.241 ;
      RECT MASK 2 100.89 82.0405 100.95 85.241 ;
      RECT MASK 2 102.052 82.0405 102.112 85.241 ;
      RECT MASK 2 105.184 82.0405 105.244 85.241 ;
      RECT MASK 2 106.346 82.0405 106.406 85.241 ;
      RECT MASK 2 107.508 82.0405 107.568 85.241 ;
      RECT MASK 2 108.67 82.0405 108.73 85.241 ;
      RECT MASK 2 111.377 82.145 111.437 82.405 ;
      RECT MASK 2 111.709 82.145 111.769 82.405 ;
      RECT MASK 2 112.041 82.145 112.101 82.405 ;
      RECT MASK 2 112.373 82.145 112.433 82.405 ;
      RECT MASK 2 112.705 82.145 112.765 82.405 ;
      RECT MASK 2 113.037 82.145 113.097 82.405 ;
      RECT MASK 2 7.408 82.242 7.468 85.241 ;
      RECT MASK 2 8.57 82.242 8.63 85.241 ;
      RECT MASK 2 9.732 82.242 9.792 85.241 ;
      RECT MASK 2 12.864 82.242 12.924 85.241 ;
      RECT MASK 2 14.026 82.242 14.086 85.241 ;
      RECT MASK 2 15.188 82.242 15.248 85.241 ;
      RECT MASK 2 16.35 82.242 16.41 85.241 ;
      RECT MASK 2 19.482 82.242 19.542 85.241 ;
      RECT MASK 2 20.644 82.242 20.704 85.241 ;
      RECT MASK 2 21.806 82.242 21.866 85.241 ;
      RECT MASK 2 22.968 82.242 23.028 85.241 ;
      RECT MASK 2 26.1 82.242 26.16 85.241 ;
      RECT MASK 2 27.262 82.242 27.322 85.241 ;
      RECT MASK 2 28.424 82.242 28.484 85.241 ;
      RECT MASK 2 29.586 82.242 29.646 85.241 ;
      RECT MASK 2 32.718 82.242 32.778 85.241 ;
      RECT MASK 2 33.88 82.242 33.94 85.241 ;
      RECT MASK 2 35.042 82.242 35.102 85.241 ;
      RECT MASK 2 36.204 82.242 36.264 85.241 ;
      RECT MASK 2 39.336 82.242 39.396 85.241 ;
      RECT MASK 2 40.498 82.242 40.558 85.241 ;
      RECT MASK 2 41.66 82.242 41.72 85.241 ;
      RECT MASK 2 42.822 82.242 42.882 85.241 ;
      RECT MASK 2 45.954 82.242 46.014 85.241 ;
      RECT MASK 2 47.116 82.242 47.176 85.241 ;
      RECT MASK 2 48.278 82.242 48.338 85.241 ;
      RECT MASK 2 49.44 82.242 49.5 85.241 ;
      RECT MASK 2 52.572 82.242 52.632 85.241 ;
      RECT MASK 2 53.734 82.242 53.794 85.241 ;
      RECT MASK 2 54.896 82.242 54.956 85.241 ;
      RECT MASK 2 56.058 82.242 56.118 85.241 ;
      RECT MASK 2 59.19 82.242 59.25 85.241 ;
      RECT MASK 2 60.352 82.242 60.412 85.241 ;
      RECT MASK 2 61.514 82.242 61.574 85.241 ;
      RECT MASK 2 62.676 82.242 62.736 85.241 ;
      RECT MASK 2 65.808 82.242 65.868 85.241 ;
      RECT MASK 2 66.97 82.242 67.03 85.241 ;
      RECT MASK 2 68.132 82.242 68.192 85.241 ;
      RECT MASK 2 69.294 82.242 69.354 85.241 ;
      RECT MASK 2 72.426 82.242 72.486 85.241 ;
      RECT MASK 2 73.588 82.242 73.648 85.241 ;
      RECT MASK 2 74.75 82.242 74.81 85.241 ;
      RECT MASK 2 75.912 82.242 75.972 85.241 ;
      RECT MASK 2 79.044 82.242 79.104 85.241 ;
      RECT MASK 2 80.206 82.242 80.266 85.241 ;
      RECT MASK 2 81.368 82.242 81.428 85.241 ;
      RECT MASK 2 82.53 82.242 82.59 85.241 ;
      RECT MASK 2 85.662 82.242 85.722 85.241 ;
      RECT MASK 2 86.824 82.242 86.884 85.241 ;
      RECT MASK 2 87.986 82.242 88.046 85.241 ;
      RECT MASK 2 89.148 82.242 89.208 85.241 ;
      RECT MASK 2 92.28 82.242 92.34 85.241 ;
      RECT MASK 2 93.442 82.242 93.502 85.241 ;
      RECT MASK 2 94.604 82.242 94.664 85.241 ;
      RECT MASK 2 95.766 82.242 95.826 85.241 ;
      RECT MASK 2 98.898 82.242 98.958 85.241 ;
      RECT MASK 2 100.06 82.242 100.12 85.241 ;
      RECT MASK 2 101.222 82.242 101.282 85.241 ;
      RECT MASK 2 102.384 82.242 102.444 85.241 ;
      RECT MASK 2 105.516 82.242 105.576 85.241 ;
      RECT MASK 2 106.678 82.242 106.738 85.241 ;
      RECT MASK 2 107.84 82.242 107.9 85.241 ;
      RECT MASK 2 109.002 82.242 109.062 85.241 ;
      RECT MASK 2 6.661 82.38 6.721 82.65 ;
      RECT MASK 2 7.823 82.38 7.883 82.65 ;
      RECT MASK 2 8.985 82.38 9.045 82.65 ;
      RECT MASK 2 10.147 82.38 10.207 82.65 ;
      RECT MASK 2 12.117 82.38 12.177 82.65 ;
      RECT MASK 2 13.279 82.38 13.339 82.65 ;
      RECT MASK 2 14.441 82.38 14.501 82.65 ;
      RECT MASK 2 15.603 82.38 15.663 82.65 ;
      RECT MASK 2 16.765 82.38 16.825 82.65 ;
      RECT MASK 2 18.735 82.38 18.795 82.65 ;
      RECT MASK 2 19.897 82.38 19.957 82.65 ;
      RECT MASK 2 21.059 82.38 21.119 82.65 ;
      RECT MASK 2 22.221 82.38 22.281 82.65 ;
      RECT MASK 2 23.383 82.38 23.443 82.65 ;
      RECT MASK 2 25.353 82.38 25.413 82.65 ;
      RECT MASK 2 26.515 82.38 26.575 82.65 ;
      RECT MASK 2 27.677 82.38 27.737 82.65 ;
      RECT MASK 2 28.839 82.38 28.899 82.65 ;
      RECT MASK 2 30.001 82.38 30.061 82.65 ;
      RECT MASK 2 31.971 82.38 32.031 82.65 ;
      RECT MASK 2 33.133 82.38 33.193 82.65 ;
      RECT MASK 2 34.295 82.38 34.355 82.65 ;
      RECT MASK 2 35.457 82.38 35.517 82.65 ;
      RECT MASK 2 36.619 82.38 36.679 82.65 ;
      RECT MASK 2 38.589 82.38 38.649 82.65 ;
      RECT MASK 2 39.751 82.38 39.811 82.65 ;
      RECT MASK 2 40.913 82.38 40.973 82.65 ;
      RECT MASK 2 42.075 82.38 42.135 82.65 ;
      RECT MASK 2 43.237 82.38 43.297 82.65 ;
      RECT MASK 2 45.207 82.38 45.267 82.65 ;
      RECT MASK 2 46.369 82.38 46.429 82.65 ;
      RECT MASK 2 47.531 82.38 47.591 82.65 ;
      RECT MASK 2 48.693 82.38 48.753 82.65 ;
      RECT MASK 2 49.855 82.38 49.915 82.65 ;
      RECT MASK 2 51.825 82.38 51.885 82.65 ;
      RECT MASK 2 52.987 82.38 53.047 82.65 ;
      RECT MASK 2 54.149 82.38 54.209 82.65 ;
      RECT MASK 2 55.311 82.38 55.371 82.65 ;
      RECT MASK 2 56.473 82.38 56.533 82.65 ;
      RECT MASK 2 65.061 82.38 65.121 82.65 ;
      RECT MASK 2 66.223 82.38 66.283 82.65 ;
      RECT MASK 2 67.385 82.38 67.445 82.65 ;
      RECT MASK 2 68.547 82.38 68.607 82.65 ;
      RECT MASK 2 69.709 82.38 69.769 82.65 ;
      RECT MASK 2 71.679 82.38 71.739 82.65 ;
      RECT MASK 2 72.841 82.38 72.901 82.65 ;
      RECT MASK 2 74.003 82.38 74.063 82.65 ;
      RECT MASK 2 75.165 82.38 75.225 82.65 ;
      RECT MASK 2 76.327 82.38 76.387 82.65 ;
      RECT MASK 2 78.297 82.38 78.357 82.65 ;
      RECT MASK 2 79.459 82.38 79.519 82.65 ;
      RECT MASK 2 80.621 82.38 80.681 82.65 ;
      RECT MASK 2 81.783 82.38 81.843 82.65 ;
      RECT MASK 2 82.945 82.38 83.005 82.65 ;
      RECT MASK 2 84.915 82.38 84.975 82.65 ;
      RECT MASK 2 86.077 82.38 86.137 82.65 ;
      RECT MASK 2 87.239 82.38 87.299 82.65 ;
      RECT MASK 2 88.401 82.38 88.461 82.65 ;
      RECT MASK 2 89.563 82.38 89.623 82.65 ;
      RECT MASK 2 91.533 82.38 91.593 82.65 ;
      RECT MASK 2 92.695 82.38 92.755 82.65 ;
      RECT MASK 2 93.857 82.38 93.917 82.65 ;
      RECT MASK 2 95.019 82.38 95.079 82.65 ;
      RECT MASK 2 96.181 82.38 96.241 82.65 ;
      RECT MASK 2 98.151 82.38 98.211 82.65 ;
      RECT MASK 2 99.313 82.38 99.373 82.65 ;
      RECT MASK 2 100.475 82.38 100.535 82.65 ;
      RECT MASK 2 101.637 82.38 101.697 82.65 ;
      RECT MASK 2 102.799 82.38 102.859 82.65 ;
      RECT MASK 2 104.769 82.38 104.829 82.65 ;
      RECT MASK 2 105.931 82.38 105.991 82.65 ;
      RECT MASK 2 107.093 82.38 107.153 82.65 ;
      RECT MASK 2 108.255 82.38 108.315 82.65 ;
      RECT MASK 2 109.417 82.38 109.477 82.65 ;
      RECT MASK 2 10.883 84.308 10.943 86.0585 ;
      RECT MASK 2 11.215 84.308 11.275 86.0585 ;
      RECT MASK 2 17.501 84.308 17.561 86.0585 ;
      RECT MASK 2 17.833 84.308 17.893 86.0585 ;
      RECT MASK 2 24.119 84.308 24.179 86.0585 ;
      RECT MASK 2 24.451 84.308 24.511 86.0585 ;
      RECT MASK 2 30.737 84.308 30.797 86.0585 ;
      RECT MASK 2 31.069 84.308 31.129 86.0585 ;
      RECT MASK 2 37.355 84.308 37.415 86.0585 ;
      RECT MASK 2 37.687 84.308 37.747 86.0585 ;
      RECT MASK 2 43.973 84.308 44.033 86.0585 ;
      RECT MASK 2 44.305 84.308 44.365 86.0585 ;
      RECT MASK 2 50.591 84.308 50.651 86.0585 ;
      RECT MASK 2 50.923 84.308 50.983 86.0585 ;
      RECT MASK 2 57.209 84.308 57.269 86.0585 ;
      RECT MASK 2 57.541 84.308 57.601 86.0585 ;
      RECT MASK 2 63.827 84.308 63.887 86.0585 ;
      RECT MASK 2 64.159 84.308 64.219 86.0585 ;
      RECT MASK 2 70.445 84.308 70.505 86.0585 ;
      RECT MASK 2 70.777 84.308 70.837 86.0585 ;
      RECT MASK 2 77.063 84.308 77.123 86.0585 ;
      RECT MASK 2 77.395 84.308 77.455 86.0585 ;
      RECT MASK 2 83.681 84.308 83.741 86.0585 ;
      RECT MASK 2 84.013 84.308 84.073 86.0585 ;
      RECT MASK 2 90.299 84.308 90.359 86.0585 ;
      RECT MASK 2 90.631 84.308 90.691 86.0585 ;
      RECT MASK 2 96.917 84.308 96.977 86.0585 ;
      RECT MASK 2 97.249 84.308 97.309 86.0585 ;
      RECT MASK 2 103.535 84.308 103.595 86.0585 ;
      RECT MASK 2 103.867 84.308 103.927 86.0585 ;
      RECT MASK 2 8.982 85.4905 9.042 86.055 ;
      RECT MASK 2 15.6 85.4905 15.66 86.055 ;
      RECT MASK 2 7.242 85.4915 7.302 86.056 ;
      RECT MASK 2 7.82 85.4915 7.88 86.056 ;
      RECT MASK 2 8.404 85.4915 8.464 86.056 ;
      RECT MASK 2 9.566 85.4915 9.626 86.056 ;
      RECT MASK 2 10.198 85.4915 10.258 86.056 ;
      RECT MASK 2 13.86 85.4915 13.92 86.056 ;
      RECT MASK 2 14.438 85.4915 14.498 86.056 ;
      RECT MASK 2 15.022 85.4915 15.082 86.056 ;
      RECT MASK 2 16.184 85.4915 16.244 86.056 ;
      RECT MASK 2 16.816 85.4915 16.876 86.056 ;
      RECT MASK 2 12.0755 85.5 12.1355 86.056 ;
      RECT MASK 2 12.698 85.5 12.758 86.056 ;
      RECT MASK 2 6.6195 85.543 6.6795 86.056 ;
      RECT MASK 2 36.326 87.021 66.476 87.081 ;
      RECT MASK 2 72.716 87.021 102.866 87.081 ;
      RECT MASK 2 25.66 87.101 30.63 87.161 ;
      RECT MASK 2 13.243 87.188 13.343 94.372 ;
      RECT MASK 2 8.381 87.21 8.441 87.49 ;
      RECT MASK 2 8.713 87.21 8.773 87.49 ;
      RECT MASK 2 9.045 87.21 9.105 87.49 ;
      RECT MASK 2 9.377 87.21 9.437 87.49 ;
      RECT MASK 2 9.709 87.21 9.769 87.49 ;
      RECT MASK 2 10.041 87.21 10.101 87.49 ;
      RECT MASK 2 10.373 87.21 10.433 87.49 ;
      RECT MASK 2 10.705 87.21 10.765 87.49 ;
      RECT MASK 2 11.037 87.21 11.097 87.49 ;
      RECT MASK 2 11.369 87.21 11.429 87.49 ;
      RECT MASK 2 11.701 87.21 11.761 87.49 ;
      RECT MASK 2 12.033 87.21 12.093 87.49 ;
      RECT MASK 2 12.365 87.21 12.425 87.49 ;
      RECT MASK 2 13.761 87.21 13.821 87.49 ;
      RECT MASK 2 14.093 87.21 14.153 87.49 ;
      RECT MASK 2 14.425 87.21 14.485 87.49 ;
      RECT MASK 2 14.591 87.21 14.651 87.49 ;
      RECT MASK 2 14.923 87.21 14.983 87.49 ;
      RECT MASK 2 15.255 87.21 15.315 87.49 ;
      RECT MASK 2 15.587 87.21 15.647 87.49 ;
      RECT MASK 2 15.919 87.21 15.979 87.49 ;
      RECT MASK 2 16.251 87.21 16.311 87.49 ;
      RECT MASK 2 16.583 87.21 16.643 87.49 ;
      RECT MASK 2 16.915 87.21 16.975 87.49 ;
      RECT MASK 2 17.979 87.21 18.039 87.49 ;
      RECT MASK 2 18.311 87.21 18.371 87.49 ;
      RECT MASK 2 18.643 87.21 18.703 87.49 ;
      RECT MASK 2 18.975 87.21 19.035 87.49 ;
      RECT MASK 2 19.307 87.21 19.367 87.49 ;
      RECT MASK 2 19.639 87.21 19.699 87.49 ;
      RECT MASK 2 19.971 87.21 20.031 87.49 ;
      RECT MASK 2 20.303 87.21 20.363 87.49 ;
      RECT MASK 2 20.635 87.21 20.695 87.49 ;
      RECT MASK 2 20.967 87.21 21.027 87.49 ;
      RECT MASK 2 21.299 87.21 21.359 87.49 ;
      RECT MASK 2 21.631 87.21 21.691 87.49 ;
      RECT MASK 2 21.963 87.21 22.023 87.49 ;
      RECT MASK 2 36.326 87.273 66.476 87.333 ;
      RECT MASK 2 72.716 87.273 102.866 87.333 ;
      RECT MASK 2 22.627 87.285 22.687 94.77 ;
      RECT MASK 2 22.959 87.285 23.019 94.77 ;
      RECT MASK 2 23.291 87.285 23.351 94.77 ;
      RECT MASK 2 23.623 87.285 23.683 94.77 ;
      RECT MASK 2 23.955 87.285 24.015 94.77 ;
      RECT MASK 2 25.66 87.363 30.63 87.423 ;
      RECT MASK 2 6.59 87.641 6.65 89.941 ;
      RECT MASK 2 9.2965 87.66 9.3565 88.912 ;
      RECT MASK 2 11.6205 87.66 11.6805 88.912 ;
      RECT MASK 2 12.0985 87.66 12.1985 90.24 ;
      RECT MASK 2 13.9925 87.66 14.0925 88.07 ;
      RECT MASK 2 14.3245 87.66 14.4245 88.39 ;
      RECT MASK 2 14.6565 87.66 14.7565 88.39 ;
      RECT MASK 2 14.9885 87.66 15.0885 88.39 ;
      RECT MASK 2 15.3205 87.66 15.4205 88.39 ;
      RECT MASK 2 15.6525 87.66 15.7525 88.39 ;
      RECT MASK 2 15.9845 87.66 16.0845 88.39 ;
      RECT MASK 2 16.3165 87.66 16.4165 88.07 ;
      RECT MASK 2 18.5625 87.66 18.6225 88.912 ;
      RECT MASK 2 18.8945 87.66 18.9545 88.912 ;
      RECT MASK 2 19.2265 87.66 19.2865 88.912 ;
      RECT MASK 2 19.5585 87.66 19.6185 88.912 ;
      RECT MASK 2 19.8905 87.66 19.9505 88.912 ;
      RECT MASK 2 20.2225 87.66 20.2825 88.912 ;
      RECT MASK 2 20.5545 87.66 20.6145 88.912 ;
      RECT MASK 2 20.8865 87.66 20.9465 88.912 ;
      RECT MASK 2 21.2185 87.66 21.2785 88.912 ;
      RECT MASK 2 108.379 87.72 108.439 96.66 ;
      RECT MASK 2 108.653 87.72 108.713 96.66 ;
      RECT MASK 2 108.927 87.72 108.987 96.66 ;
      RECT MASK 2 109.201 87.72 109.261 96.66 ;
      RECT MASK 2 109.475 87.72 109.535 96.66 ;
      RECT MASK 2 109.749 87.72 109.809 96.66 ;
      RECT MASK 2 110.023 87.72 110.083 96.66 ;
      RECT MASK 2 110.297 87.72 110.357 96.66 ;
      RECT MASK 2 110.571 87.72 110.631 96.66 ;
      RECT MASK 2 110.845 87.72 110.905 96.66 ;
      RECT MASK 2 111.119 87.72 111.179 96.66 ;
      RECT MASK 2 111.393 87.72 111.453 96.66 ;
      RECT MASK 2 111.667 87.72 111.727 96.66 ;
      RECT MASK 2 111.941 87.72 112.001 96.66 ;
      RECT MASK 2 112.215 87.72 112.275 96.66 ;
      RECT MASK 2 112.489 87.72 112.549 96.66 ;
      RECT MASK 2 112.763 87.72 112.823 96.66 ;
      RECT MASK 2 113.037 87.72 113.097 96.66 ;
      RECT MASK 2 113.311 87.72 113.371 96.66 ;
      RECT MASK 2 113.585 87.72 113.645 96.66 ;
      RECT MASK 2 113.859 87.72 113.919 96.66 ;
      RECT MASK 2 114.133 87.72 114.193 96.66 ;
      RECT MASK 2 114.407 87.72 114.467 96.66 ;
      RECT MASK 2 114.681 87.72 114.741 96.66 ;
      RECT MASK 2 114.955 87.72 115.015 96.66 ;
      RECT MASK 2 115.229 87.72 115.289 96.66 ;
      RECT MASK 2 115.503 87.72 115.563 96.66 ;
      RECT MASK 2 115.777 87.72 115.837 96.66 ;
      RECT MASK 2 116.051 87.72 116.111 96.66 ;
      RECT MASK 2 116.325 87.72 116.385 96.66 ;
      RECT MASK 2 36.326 87.921 36.778 87.981 ;
      RECT MASK 2 37.048 87.921 65.754 87.981 ;
      RECT MASK 2 66.024 87.921 66.476 87.981 ;
      RECT MASK 2 72.716 87.921 73.168 87.981 ;
      RECT MASK 2 73.438 87.921 102.144 87.981 ;
      RECT MASK 2 102.414 87.921 102.866 87.981 ;
      RECT MASK 2 25.66 87.957 25.944 88.017 ;
      RECT MASK 2 26.205 87.957 30.085 88.017 ;
      RECT MASK 2 30.346 87.957 30.63 88.017 ;
      RECT MASK 2 36.326 88.173 36.778 88.233 ;
      RECT MASK 2 37.048 88.173 65.754 88.233 ;
      RECT MASK 2 66.024 88.173 66.476 88.233 ;
      RECT MASK 2 72.716 88.173 73.168 88.233 ;
      RECT MASK 2 73.438 88.173 102.144 88.233 ;
      RECT MASK 2 102.414 88.173 102.866 88.233 ;
      RECT MASK 2 9.6285 88.3795 9.6885 88.912 ;
      RECT MASK 2 9.9605 88.3795 10.0205 88.912 ;
      RECT MASK 2 10.2925 88.3795 10.3525 88.912 ;
      RECT MASK 2 10.6245 88.3795 10.6845 88.912 ;
      RECT MASK 2 10.9565 88.3795 11.0165 88.912 ;
      RECT MASK 2 11.2885 88.3795 11.3485 88.912 ;
      RECT MASK 2 25.66 88.541 30.63 88.601 ;
      RECT MASK 2 14.3445 88.595 14.4045 88.912 ;
      RECT MASK 2 14.6765 88.595 14.7365 88.912 ;
      RECT MASK 2 15.0085 88.595 15.0685 88.912 ;
      RECT MASK 2 15.3405 88.595 15.4005 88.912 ;
      RECT MASK 2 15.6725 88.595 15.7325 88.912 ;
      RECT MASK 2 16.0045 88.595 16.0645 88.912 ;
      RECT MASK 2 25.66 88.803 30.63 88.863 ;
      RECT MASK 2 36.326 88.821 66.476 88.881 ;
      RECT MASK 2 72.716 88.821 102.866 88.881 ;
      RECT MASK 2 9.0475 89.05 9.1075 89.33 ;
      RECT MASK 2 9.3795 89.05 9.4395 89.33 ;
      RECT MASK 2 11.7035 89.05 11.7635 89.33 ;
      RECT MASK 2 14.0955 89.05 14.1555 89.33 ;
      RECT MASK 2 14.4275 89.05 14.4875 89.33 ;
      RECT MASK 2 16.0875 89.05 16.1475 89.33 ;
      RECT MASK 2 18.6455 89.05 18.7055 89.33 ;
      RECT MASK 2 20.9695 89.05 21.0295 89.33 ;
      RECT MASK 2 21.3015 89.05 21.3615 89.33 ;
      RECT MASK 2 36.326 89.073 66.476 89.133 ;
      RECT MASK 2 72.716 89.073 102.866 89.133 ;
      RECT MASK 2 9.7115 89.0915 9.7715 89.2865 ;
      RECT MASK 2 10.0435 89.0915 10.1035 89.2865 ;
      RECT MASK 2 10.3755 89.0915 10.4355 89.2865 ;
      RECT MASK 2 10.7075 89.0915 10.7675 89.2865 ;
      RECT MASK 2 11.0395 89.0915 11.0995 89.2865 ;
      RECT MASK 2 14.7595 89.0915 14.8195 89.2865 ;
      RECT MASK 2 15.0915 89.0915 15.1515 89.2865 ;
      RECT MASK 2 15.4235 89.0915 15.4835 89.2865 ;
      RECT MASK 2 19.3095 89.0915 19.3695 89.2865 ;
      RECT MASK 2 19.6415 89.0915 19.7015 89.2865 ;
      RECT MASK 2 19.9735 89.0915 20.0335 89.2865 ;
      RECT MASK 2 20.3055 89.0915 20.3655 89.2865 ;
      RECT MASK 2 20.6375 89.0915 20.6975 89.2865 ;
      RECT MASK 2 25.66 89.441 30.63 89.501 ;
      RECT MASK 2 18.5625 89.455 18.6225 90.24 ;
      RECT MASK 2 18.8945 89.455 18.9545 90.24 ;
      RECT MASK 2 19.2265 89.455 19.2865 90.24 ;
      RECT MASK 2 19.5585 89.455 19.6185 90.24 ;
      RECT MASK 2 19.8905 89.455 19.9505 90.24 ;
      RECT MASK 2 20.2225 89.455 20.2825 90.24 ;
      RECT MASK 2 20.5545 89.455 20.6145 90.24 ;
      RECT MASK 2 20.8865 89.455 20.9465 90.24 ;
      RECT MASK 2 21.2185 89.455 21.2785 90.24 ;
      RECT MASK 2 9.2965 89.468 9.3565 90.24 ;
      RECT MASK 2 9.6285 89.468 9.6885 89.8075 ;
      RECT MASK 2 9.9605 89.468 10.0205 89.8075 ;
      RECT MASK 2 10.2925 89.468 10.3525 89.8075 ;
      RECT MASK 2 10.6245 89.468 10.6845 89.8075 ;
      RECT MASK 2 10.9565 89.468 11.0165 89.8075 ;
      RECT MASK 2 11.2885 89.468 11.3485 89.8075 ;
      RECT MASK 2 11.6205 89.468 11.6805 90.24 ;
      RECT MASK 2 14.3445 89.468 14.4045 89.692 ;
      RECT MASK 2 14.6765 89.468 14.7365 89.692 ;
      RECT MASK 2 15.0085 89.468 15.0685 89.692 ;
      RECT MASK 2 15.3405 89.468 15.4005 89.692 ;
      RECT MASK 2 15.6725 89.468 15.7325 89.692 ;
      RECT MASK 2 16.0045 89.468 16.0645 89.692 ;
      RECT MASK 2 25.66 89.703 30.63 89.763 ;
      RECT MASK 2 36.326 89.721 36.778 89.781 ;
      RECT MASK 2 37.048 89.721 65.754 89.781 ;
      RECT MASK 2 66.024 89.721 66.476 89.781 ;
      RECT MASK 2 72.716 89.721 73.168 89.781 ;
      RECT MASK 2 73.438 89.721 102.144 89.781 ;
      RECT MASK 2 102.414 89.721 102.866 89.781 ;
      RECT MASK 2 13.9925 89.905 14.0925 90.25 ;
      RECT MASK 2 14.3245 89.905 14.4245 90.25 ;
      RECT MASK 2 14.6565 89.905 14.7565 90.25 ;
      RECT MASK 2 14.9885 89.905 15.0885 90.25 ;
      RECT MASK 2 15.3205 89.905 15.4205 90.25 ;
      RECT MASK 2 15.6525 89.905 15.7525 90.25 ;
      RECT MASK 2 15.9845 89.905 16.0845 90.25 ;
      RECT MASK 2 16.3165 89.905 16.4165 90.25 ;
      RECT MASK 2 36.326 89.973 36.778 90.033 ;
      RECT MASK 2 37.048 89.973 65.754 90.033 ;
      RECT MASK 2 66.024 89.973 66.476 90.033 ;
      RECT MASK 2 72.716 89.973 73.168 90.033 ;
      RECT MASK 2 73.438 89.973 102.144 90.033 ;
      RECT MASK 2 102.414 89.973 102.866 90.033 ;
      RECT MASK 2 6.59 90.061 6.65 90.355 ;
      RECT MASK 2 25.66 90.297 25.944 90.357 ;
      RECT MASK 2 26.205 90.297 30.085 90.357 ;
      RECT MASK 2 30.346 90.297 30.63 90.357 ;
      RECT MASK 2 8.381 90.42 8.441 90.7 ;
      RECT MASK 2 8.713 90.42 8.773 90.7 ;
      RECT MASK 2 9.045 90.42 9.105 90.7 ;
      RECT MASK 2 9.377 90.42 9.437 90.7 ;
      RECT MASK 2 9.709 90.42 9.769 90.7 ;
      RECT MASK 2 10.041 90.42 10.101 90.7 ;
      RECT MASK 2 10.373 90.42 10.433 90.7 ;
      RECT MASK 2 10.705 90.42 10.765 90.7 ;
      RECT MASK 2 11.037 90.42 11.097 90.7 ;
      RECT MASK 2 11.369 90.42 11.429 90.7 ;
      RECT MASK 2 11.701 90.42 11.761 90.7 ;
      RECT MASK 2 12.033 90.42 12.093 90.7 ;
      RECT MASK 2 12.365 90.42 12.425 90.7 ;
      RECT MASK 2 13.761 90.42 13.821 90.7 ;
      RECT MASK 2 14.093 90.42 14.153 90.7 ;
      RECT MASK 2 14.425 90.42 14.485 90.7 ;
      RECT MASK 2 14.591 90.42 14.651 90.7 ;
      RECT MASK 2 14.923 90.42 14.983 90.7 ;
      RECT MASK 2 15.255 90.42 15.315 90.7 ;
      RECT MASK 2 15.587 90.42 15.647 90.7 ;
      RECT MASK 2 15.919 90.42 15.979 90.7 ;
      RECT MASK 2 16.251 90.42 16.311 90.7 ;
      RECT MASK 2 16.583 90.42 16.643 90.7 ;
      RECT MASK 2 16.915 90.42 16.975 90.7 ;
      RECT MASK 2 17.979 90.42 18.039 90.7 ;
      RECT MASK 2 18.311 90.42 18.371 90.7 ;
      RECT MASK 2 18.643 90.42 18.703 90.7 ;
      RECT MASK 2 18.975 90.42 19.035 90.7 ;
      RECT MASK 2 19.307 90.42 19.367 90.7 ;
      RECT MASK 2 19.639 90.42 19.699 90.7 ;
      RECT MASK 2 19.971 90.42 20.031 90.7 ;
      RECT MASK 2 20.303 90.42 20.363 90.7 ;
      RECT MASK 2 20.635 90.42 20.695 90.7 ;
      RECT MASK 2 20.967 90.42 21.027 90.7 ;
      RECT MASK 2 21.299 90.42 21.359 90.7 ;
      RECT MASK 2 21.631 90.42 21.691 90.7 ;
      RECT MASK 2 21.963 90.42 22.023 90.7 ;
      RECT MASK 2 36.326 90.621 66.476 90.681 ;
      RECT MASK 2 72.716 90.621 102.866 90.681 ;
      RECT MASK 2 6.59 90.73 6.65 93.451 ;
      RECT MASK 2 8.381 90.86 8.441 91.14 ;
      RECT MASK 2 8.713 90.86 8.773 91.14 ;
      RECT MASK 2 9.045 90.86 9.105 91.14 ;
      RECT MASK 2 9.377 90.86 9.437 91.14 ;
      RECT MASK 2 9.709 90.86 9.769 91.14 ;
      RECT MASK 2 10.041 90.86 10.101 91.14 ;
      RECT MASK 2 10.373 90.86 10.433 91.14 ;
      RECT MASK 2 10.705 90.86 10.765 91.14 ;
      RECT MASK 2 11.037 90.86 11.097 91.14 ;
      RECT MASK 2 11.369 90.86 11.429 91.14 ;
      RECT MASK 2 11.701 90.86 11.761 91.14 ;
      RECT MASK 2 12.033 90.86 12.093 91.14 ;
      RECT MASK 2 12.365 90.86 12.425 91.14 ;
      RECT MASK 2 13.761 90.86 13.821 91.14 ;
      RECT MASK 2 14.093 90.86 14.153 91.14 ;
      RECT MASK 2 14.425 90.86 14.485 91.14 ;
      RECT MASK 2 14.591 90.86 14.651 91.14 ;
      RECT MASK 2 14.923 90.86 14.983 91.14 ;
      RECT MASK 2 15.255 90.86 15.315 91.14 ;
      RECT MASK 2 15.587 90.86 15.647 91.14 ;
      RECT MASK 2 15.919 90.86 15.979 91.14 ;
      RECT MASK 2 16.251 90.86 16.311 91.14 ;
      RECT MASK 2 16.583 90.86 16.643 91.14 ;
      RECT MASK 2 16.915 90.86 16.975 91.14 ;
      RECT MASK 2 17.979 90.86 18.039 91.14 ;
      RECT MASK 2 18.311 90.86 18.371 91.14 ;
      RECT MASK 2 18.643 90.86 18.703 91.14 ;
      RECT MASK 2 18.975 90.86 19.035 91.14 ;
      RECT MASK 2 19.307 90.86 19.367 91.14 ;
      RECT MASK 2 19.639 90.86 19.699 91.14 ;
      RECT MASK 2 19.971 90.86 20.031 91.14 ;
      RECT MASK 2 20.303 90.86 20.363 91.14 ;
      RECT MASK 2 20.635 90.86 20.695 91.14 ;
      RECT MASK 2 20.967 90.86 21.027 91.14 ;
      RECT MASK 2 21.299 90.86 21.359 91.14 ;
      RECT MASK 2 21.631 90.86 21.691 91.14 ;
      RECT MASK 2 21.963 90.86 22.023 91.14 ;
      RECT MASK 2 36.326 90.873 66.476 90.933 ;
      RECT MASK 2 72.716 90.873 102.866 90.933 ;
      RECT MASK 2 25.66 90.881 30.63 90.941 ;
      RECT MASK 2 25.66 91.143 30.63 91.203 ;
      RECT MASK 2 13.9925 91.31 14.0925 91.655 ;
      RECT MASK 2 14.3245 91.31 14.4245 91.655 ;
      RECT MASK 2 14.6565 91.31 14.7565 91.655 ;
      RECT MASK 2 14.9885 91.31 15.0885 91.655 ;
      RECT MASK 2 15.3205 91.31 15.4205 91.655 ;
      RECT MASK 2 15.6525 91.31 15.7525 91.655 ;
      RECT MASK 2 15.9845 91.31 16.0845 91.655 ;
      RECT MASK 2 16.3165 91.31 16.4165 91.655 ;
      RECT MASK 2 8.969 91.32 9.029 92.092 ;
      RECT MASK 2 11.293 91.32 11.353 92.092 ;
      RECT MASK 2 11.771 91.32 11.871 93.9 ;
      RECT MASK 2 18.5625 91.32 18.6225 92.105 ;
      RECT MASK 2 18.8945 91.32 18.9545 92.105 ;
      RECT MASK 2 19.2265 91.32 19.2865 92.105 ;
      RECT MASK 2 19.5585 91.32 19.6185 92.105 ;
      RECT MASK 2 19.8905 91.32 19.9505 92.105 ;
      RECT MASK 2 20.2225 91.32 20.2825 92.105 ;
      RECT MASK 2 20.5545 91.32 20.6145 92.105 ;
      RECT MASK 2 20.8865 91.32 20.9465 92.105 ;
      RECT MASK 2 21.2185 91.32 21.2785 92.105 ;
      RECT MASK 2 36.326 91.521 36.778 91.581 ;
      RECT MASK 2 37.048 91.521 65.754 91.581 ;
      RECT MASK 2 66.024 91.521 66.476 91.581 ;
      RECT MASK 2 72.716 91.521 73.168 91.581 ;
      RECT MASK 2 73.438 91.521 102.144 91.581 ;
      RECT MASK 2 102.414 91.521 102.866 91.581 ;
      RECT MASK 2 25.1675 91.5285 31.1545 91.7685 ;
      RECT MASK 2 9.301 91.7525 9.361 92.092 ;
      RECT MASK 2 9.633 91.7525 9.693 92.092 ;
      RECT MASK 2 9.965 91.7525 10.025 92.092 ;
      RECT MASK 2 10.297 91.7525 10.357 92.092 ;
      RECT MASK 2 10.629 91.7525 10.689 92.092 ;
      RECT MASK 2 10.961 91.7525 11.021 92.092 ;
      RECT MASK 2 36.326 91.773 36.778 91.833 ;
      RECT MASK 2 37.048 91.773 65.754 91.833 ;
      RECT MASK 2 66.024 91.773 66.476 91.833 ;
      RECT MASK 2 72.716 91.773 73.168 91.833 ;
      RECT MASK 2 73.438 91.773 102.144 91.833 ;
      RECT MASK 2 102.414 91.773 102.866 91.833 ;
      RECT MASK 2 14.3445 91.868 14.4045 92.092 ;
      RECT MASK 2 14.6765 91.868 14.7365 92.095 ;
      RECT MASK 2 15.0085 91.868 15.0685 92.095 ;
      RECT MASK 2 15.3405 91.868 15.4005 92.095 ;
      RECT MASK 2 15.6725 91.868 15.7325 92.095 ;
      RECT MASK 2 16.0045 91.868 16.0645 92.092 ;
      RECT MASK 2 8.72 92.23 8.78 92.51 ;
      RECT MASK 2 9.052 92.23 9.112 92.51 ;
      RECT MASK 2 11.376 92.23 11.436 92.51 ;
      RECT MASK 2 14.0955 92.23 14.1555 92.51 ;
      RECT MASK 2 14.4275 92.23 14.4875 92.51 ;
      RECT MASK 2 16.0875 92.23 16.1475 92.51 ;
      RECT MASK 2 18.6455 92.23 18.7055 92.51 ;
      RECT MASK 2 20.9695 92.23 21.0295 92.51 ;
      RECT MASK 2 21.3015 92.23 21.3615 92.51 ;
      RECT MASK 2 9.716 92.2735 9.776 92.4685 ;
      RECT MASK 2 10.048 92.2735 10.108 92.4685 ;
      RECT MASK 2 10.38 92.2735 10.44 92.4685 ;
      RECT MASK 2 10.712 92.2735 10.772 92.4685 ;
      RECT MASK 2 14.7595 92.2735 14.8195 92.4685 ;
      RECT MASK 2 15.0915 92.2735 15.1515 92.4685 ;
      RECT MASK 2 15.4235 92.2735 15.4835 92.4685 ;
      RECT MASK 2 19.3095 92.2735 19.3695 92.4685 ;
      RECT MASK 2 19.6415 92.2735 19.7015 92.4685 ;
      RECT MASK 2 19.9735 92.2735 20.0335 92.4685 ;
      RECT MASK 2 20.3055 92.2735 20.3655 92.4685 ;
      RECT MASK 2 20.6375 92.2735 20.6975 92.4685 ;
      RECT MASK 2 36.326 92.421 66.476 92.481 ;
      RECT MASK 2 72.716 92.421 102.866 92.481 ;
      RECT MASK 2 8.969 92.648 9.029 93.9 ;
      RECT MASK 2 9.301 92.648 9.361 93.1805 ;
      RECT MASK 2 9.633 92.648 9.693 93.1805 ;
      RECT MASK 2 9.965 92.648 10.025 93.1805 ;
      RECT MASK 2 10.297 92.648 10.357 93.1805 ;
      RECT MASK 2 10.629 92.648 10.689 93.1805 ;
      RECT MASK 2 10.961 92.648 11.021 93.1805 ;
      RECT MASK 2 11.293 92.648 11.353 93.9 ;
      RECT MASK 2 14.3445 92.648 14.4045 92.965 ;
      RECT MASK 2 14.6765 92.648 14.7365 92.965 ;
      RECT MASK 2 15.0085 92.648 15.0685 92.965 ;
      RECT MASK 2 15.3405 92.648 15.4005 92.965 ;
      RECT MASK 2 15.6725 92.648 15.7325 92.965 ;
      RECT MASK 2 16.0045 92.648 16.0645 92.965 ;
      RECT MASK 2 18.5625 92.648 18.6225 93.9 ;
      RECT MASK 2 18.8945 92.648 18.9545 93.9 ;
      RECT MASK 2 19.2265 92.648 19.2865 93.9 ;
      RECT MASK 2 19.5585 92.648 19.6185 93.9 ;
      RECT MASK 2 19.8905 92.648 19.9505 93.9 ;
      RECT MASK 2 20.2225 92.648 20.2825 93.9 ;
      RECT MASK 2 20.5545 92.648 20.6145 93.9 ;
      RECT MASK 2 20.8865 92.648 20.9465 93.9 ;
      RECT MASK 2 21.2185 92.648 21.2785 93.9 ;
      RECT MASK 2 36.326 92.673 66.476 92.733 ;
      RECT MASK 2 72.716 92.673 102.866 92.733 ;
      RECT MASK 2 14.3245 93.17 14.4245 93.9 ;
      RECT MASK 2 14.6565 93.17 14.7565 93.9 ;
      RECT MASK 2 14.9885 93.17 15.0885 93.9 ;
      RECT MASK 2 15.3205 93.17 15.4205 93.9 ;
      RECT MASK 2 15.6525 93.17 15.7525 93.9 ;
      RECT MASK 2 15.9845 93.17 16.0845 93.9 ;
      RECT MASK 2 36.326 93.321 36.778 93.381 ;
      RECT MASK 2 37.048 93.321 65.754 93.381 ;
      RECT MASK 2 66.024 93.321 66.476 93.381 ;
      RECT MASK 2 72.716 93.321 73.168 93.381 ;
      RECT MASK 2 73.438 93.321 102.144 93.381 ;
      RECT MASK 2 102.414 93.321 102.866 93.381 ;
      RECT MASK 2 13.9925 93.49 14.0925 93.9 ;
      RECT MASK 2 16.3165 93.49 16.4165 93.9 ;
      RECT MASK 2 36.326 93.573 36.778 93.633 ;
      RECT MASK 2 37.048 93.573 65.754 93.633 ;
      RECT MASK 2 66.024 93.573 66.476 93.633 ;
      RECT MASK 2 72.716 93.573 73.168 93.633 ;
      RECT MASK 2 73.438 93.573 102.144 93.633 ;
      RECT MASK 2 102.414 93.573 102.866 93.633 ;
      RECT MASK 2 8.381 94.07 8.441 94.35 ;
      RECT MASK 2 8.713 94.07 8.773 94.35 ;
      RECT MASK 2 9.045 94.07 9.105 94.35 ;
      RECT MASK 2 9.377 94.07 9.437 94.35 ;
      RECT MASK 2 9.709 94.07 9.769 94.35 ;
      RECT MASK 2 10.041 94.07 10.101 94.35 ;
      RECT MASK 2 10.373 94.07 10.433 94.35 ;
      RECT MASK 2 10.705 94.07 10.765 94.35 ;
      RECT MASK 2 11.037 94.07 11.097 94.35 ;
      RECT MASK 2 11.369 94.07 11.429 94.35 ;
      RECT MASK 2 11.701 94.07 11.761 94.35 ;
      RECT MASK 2 12.033 94.07 12.093 94.35 ;
      RECT MASK 2 12.365 94.07 12.425 94.35 ;
      RECT MASK 2 13.761 94.07 13.821 94.35 ;
      RECT MASK 2 14.093 94.07 14.153 94.35 ;
      RECT MASK 2 14.425 94.07 14.485 94.35 ;
      RECT MASK 2 14.591 94.07 14.651 94.35 ;
      RECT MASK 2 14.923 94.07 14.983 94.35 ;
      RECT MASK 2 15.255 94.07 15.315 94.35 ;
      RECT MASK 2 15.587 94.07 15.647 94.35 ;
      RECT MASK 2 15.919 94.07 15.979 94.35 ;
      RECT MASK 2 16.251 94.07 16.311 94.35 ;
      RECT MASK 2 16.583 94.07 16.643 94.35 ;
      RECT MASK 2 16.915 94.07 16.975 94.35 ;
      RECT MASK 2 17.979 94.07 18.039 94.35 ;
      RECT MASK 2 18.311 94.07 18.371 94.35 ;
      RECT MASK 2 18.643 94.07 18.703 94.35 ;
      RECT MASK 2 18.975 94.07 19.035 94.35 ;
      RECT MASK 2 19.307 94.07 19.367 94.35 ;
      RECT MASK 2 19.639 94.07 19.699 94.35 ;
      RECT MASK 2 19.971 94.07 20.031 94.35 ;
      RECT MASK 2 20.303 94.07 20.363 94.35 ;
      RECT MASK 2 20.635 94.07 20.695 94.35 ;
      RECT MASK 2 20.967 94.07 21.027 94.35 ;
      RECT MASK 2 21.299 94.07 21.359 94.35 ;
      RECT MASK 2 21.631 94.07 21.691 94.35 ;
      RECT MASK 2 21.963 94.07 22.023 94.35 ;
      RECT MASK 2 36.326 94.221 66.476 94.281 ;
      RECT MASK 2 72.716 94.221 102.866 94.281 ;
      RECT MASK 2 36.326 94.473 66.476 94.533 ;
      RECT MASK 2 72.716 94.473 102.866 94.533 ;
      RECT MASK 2 24.287 94.53 24.347 94.77 ;
      RECT MASK 2 24.619 94.53 24.679 94.77 ;
      RECT MASK 2 24.951 94.53 25.011 94.77 ;
      RECT MASK 2 25.283 94.53 25.343 94.77 ;
      RECT MASK 2 25.615 94.53 25.675 94.77 ;
      RECT MASK 2 25.947 94.53 26.007 94.77 ;
      RECT MASK 2 26.279 94.53 26.339 94.77 ;
      RECT MASK 2 26.611 94.53 26.671 94.77 ;
      RECT MASK 2 26.943 94.53 27.003 94.77 ;
      RECT MASK 2 27.275 94.53 27.335 94.77 ;
      RECT MASK 2 27.607 94.53 27.667 94.77 ;
      RECT MASK 2 27.939 94.53 27.999 94.77 ;
      RECT MASK 2 28.271 94.53 28.331 94.77 ;
      RECT MASK 2 28.603 94.53 28.663 94.77 ;
      RECT MASK 2 28.935 94.53 28.995 94.77 ;
      RECT MASK 2 29.267 94.53 29.327 94.77 ;
      RECT MASK 2 29.599 94.53 29.659 94.77 ;
      RECT MASK 2 29.931 94.53 29.991 94.77 ;
      RECT MASK 2 30.263 94.53 30.323 94.77 ;
      RECT MASK 2 30.595 94.53 30.655 94.77 ;
      RECT MASK 2 30.927 94.53 30.987 94.77 ;
      RECT MASK 2 31.259 94.53 31.319 94.77 ;
      RECT MASK 2 22.627 94.95 22.687 95.19 ;
      RECT MASK 2 22.959 94.95 23.019 95.19 ;
      RECT MASK 2 23.291 94.95 23.351 95.19 ;
      RECT MASK 2 23.623 94.95 23.683 95.19 ;
      RECT MASK 2 23.955 94.95 24.015 95.19 ;
      RECT MASK 2 24.287 94.95 24.347 95.19 ;
      RECT MASK 2 24.619 94.95 24.679 95.19 ;
      RECT MASK 2 24.951 94.95 25.011 95.19 ;
      RECT MASK 2 25.283 94.95 25.343 95.19 ;
      RECT MASK 2 25.615 94.95 25.675 95.19 ;
      RECT MASK 2 25.947 94.95 26.007 95.19 ;
      RECT MASK 2 26.279 94.95 26.339 95.19 ;
      RECT MASK 2 26.611 94.95 26.671 95.19 ;
      RECT MASK 2 26.943 94.95 27.003 95.19 ;
      RECT MASK 2 27.275 94.95 27.335 95.19 ;
      RECT MASK 2 27.607 94.95 27.667 95.19 ;
      RECT MASK 2 27.939 94.95 27.999 95.19 ;
      RECT MASK 2 28.271 94.95 28.331 95.19 ;
      RECT MASK 2 28.603 94.95 28.663 95.19 ;
      RECT MASK 2 28.935 94.95 28.995 95.19 ;
      RECT MASK 2 29.267 94.95 29.327 95.19 ;
      RECT MASK 2 29.599 94.95 29.659 95.19 ;
      RECT MASK 2 29.931 94.95 29.991 95.19 ;
      RECT MASK 2 30.263 94.95 30.323 95.19 ;
      RECT MASK 2 30.595 94.95 30.655 95.19 ;
      RECT MASK 2 30.927 94.95 30.987 95.19 ;
      RECT MASK 2 31.259 94.95 31.319 95.19 ;
      RECT MASK 2 22.627 95.37 22.687 95.61 ;
      RECT MASK 2 22.959 95.37 23.019 95.61 ;
      RECT MASK 2 23.291 95.37 23.351 95.61 ;
      RECT MASK 2 23.623 95.37 23.683 95.61 ;
      RECT MASK 2 23.955 95.37 24.015 95.61 ;
      RECT MASK 2 24.287 95.37 24.347 95.61 ;
      RECT MASK 2 24.619 95.37 24.679 95.61 ;
      RECT MASK 2 24.951 95.37 25.011 95.61 ;
      RECT MASK 2 25.283 95.37 25.343 95.61 ;
      RECT MASK 2 25.615 95.37 25.675 95.61 ;
      RECT MASK 2 25.947 95.37 26.007 95.61 ;
      RECT MASK 2 26.279 95.37 26.339 95.61 ;
      RECT MASK 2 26.611 95.37 26.671 95.61 ;
      RECT MASK 2 26.943 95.37 27.003 95.61 ;
      RECT MASK 2 27.275 95.37 27.335 95.61 ;
      RECT MASK 2 27.607 95.37 27.667 95.61 ;
      RECT MASK 2 27.939 95.37 27.999 95.61 ;
      RECT MASK 2 28.271 95.37 28.331 95.61 ;
      RECT MASK 2 28.603 95.37 28.663 95.61 ;
      RECT MASK 2 28.935 95.37 28.995 95.61 ;
      RECT MASK 2 29.267 95.37 29.327 95.61 ;
      RECT MASK 2 29.599 95.37 29.659 95.61 ;
      RECT MASK 2 29.931 95.37 29.991 95.61 ;
      RECT MASK 2 30.263 95.37 30.323 95.61 ;
      RECT MASK 2 30.595 95.37 30.655 95.61 ;
      RECT MASK 2 30.927 95.37 30.987 95.61 ;
      RECT MASK 2 31.259 95.37 31.319 95.61 ;
      RECT MASK 2 22.627 95.79 22.687 96.03 ;
      RECT MASK 2 22.959 95.79 23.019 96.03 ;
      RECT MASK 2 23.291 95.79 23.351 96.03 ;
      RECT MASK 2 23.623 95.79 23.683 96.03 ;
      RECT MASK 2 23.955 95.79 24.015 96.03 ;
      RECT MASK 2 24.287 95.79 24.347 96.03 ;
      RECT MASK 2 24.619 95.79 24.679 96.03 ;
      RECT MASK 2 24.951 95.79 25.011 96.03 ;
      RECT MASK 2 25.283 95.79 25.343 96.03 ;
      RECT MASK 2 25.615 95.79 25.675 96.03 ;
      RECT MASK 2 25.947 95.79 26.007 96.03 ;
      RECT MASK 2 26.279 95.79 26.339 96.03 ;
      RECT MASK 2 26.611 95.79 26.671 96.03 ;
      RECT MASK 2 26.943 95.79 27.003 96.03 ;
      RECT MASK 2 27.275 95.79 27.335 96.03 ;
      RECT MASK 2 27.607 95.79 27.667 96.03 ;
      RECT MASK 2 27.939 95.79 27.999 96.03 ;
      RECT MASK 2 28.271 95.79 28.331 96.03 ;
      RECT MASK 2 28.603 95.79 28.663 96.03 ;
      RECT MASK 2 28.935 95.79 28.995 96.03 ;
      RECT MASK 2 29.267 95.79 29.327 96.03 ;
      RECT MASK 2 29.599 95.79 29.659 96.03 ;
      RECT MASK 2 29.931 95.79 29.991 96.03 ;
      RECT MASK 2 30.263 95.79 30.323 96.03 ;
      RECT MASK 2 30.595 95.79 30.655 96.03 ;
      RECT MASK 2 30.927 95.79 30.987 96.03 ;
      RECT MASK 2 31.259 95.79 31.319 96.03 ;
      RECT MASK 2 31.591 95.79 31.651 96.03 ;
      RECT MASK 2 31.923 95.79 31.983 96.03 ;
      RECT MASK 2 32.255 95.79 32.315 96.03 ;
      RECT MASK 2 32.587 95.79 32.647 96.03 ;
      RECT MASK 2 32.919 95.79 32.979 96.03 ;
      RECT MASK 2 33.251 95.79 33.311 96.03 ;
      RECT MASK 2 33.583 95.79 33.643 96.03 ;
      RECT MASK 2 33.915 95.79 33.975 96.03 ;
      RECT MASK 2 34.247 95.79 34.307 96.03 ;
      RECT MASK 2 34.579 95.79 34.639 96.03 ;
      RECT MASK 2 34.911 95.79 34.971 96.03 ;
      RECT MASK 2 35.243 95.79 35.303 96.03 ;
      RECT MASK 2 35.575 95.79 35.635 96.03 ;
      RECT MASK 2 35.907 95.79 35.967 96.03 ;
      RECT MASK 2 36.239 95.79 36.299 96.03 ;
      RECT MASK 2 36.571 95.79 36.631 96.03 ;
      RECT MASK 2 22.627 96.21 22.687 96.45 ;
      RECT MASK 2 22.959 96.21 23.019 96.45 ;
      RECT MASK 2 23.291 96.21 23.351 96.45 ;
      RECT MASK 2 23.623 96.21 23.683 96.45 ;
      RECT MASK 2 23.955 96.21 24.015 96.45 ;
      RECT MASK 2 24.287 96.21 24.347 96.45 ;
      RECT MASK 2 24.619 96.21 24.679 96.45 ;
      RECT MASK 2 24.951 96.21 25.011 96.45 ;
      RECT MASK 2 25.283 96.21 25.343 96.45 ;
      RECT MASK 2 25.615 96.21 25.675 96.45 ;
      RECT MASK 2 25.947 96.21 26.007 96.45 ;
      RECT MASK 2 26.279 96.21 26.339 96.45 ;
      RECT MASK 2 26.611 96.21 26.671 96.45 ;
      RECT MASK 2 26.943 96.21 27.003 96.45 ;
      RECT MASK 2 27.275 96.21 27.335 96.45 ;
      RECT MASK 2 27.607 96.21 27.667 96.45 ;
      RECT MASK 2 27.939 96.21 27.999 96.45 ;
      RECT MASK 2 28.271 96.21 28.331 96.45 ;
      RECT MASK 2 28.603 96.21 28.663 96.45 ;
      RECT MASK 2 28.935 96.21 28.995 96.45 ;
      RECT MASK 2 29.267 96.21 29.327 96.45 ;
      RECT MASK 2 29.599 96.21 29.659 96.45 ;
      RECT MASK 2 29.931 96.21 29.991 96.45 ;
      RECT MASK 2 30.263 96.21 30.323 96.45 ;
      RECT MASK 2 30.595 96.21 30.655 96.45 ;
      RECT MASK 2 30.927 96.21 30.987 96.45 ;
      RECT MASK 2 31.259 96.21 31.319 96.45 ;
      RECT MASK 2 31.591 96.21 31.651 96.45 ;
      RECT MASK 2 31.923 96.21 31.983 96.45 ;
      RECT MASK 2 32.255 96.21 32.315 96.45 ;
      RECT MASK 2 32.587 96.21 32.647 96.45 ;
      RECT MASK 2 32.919 96.21 32.979 96.45 ;
      RECT MASK 2 33.251 96.21 33.311 96.45 ;
      RECT MASK 2 33.583 96.21 33.643 96.45 ;
      RECT MASK 2 33.915 96.21 33.975 96.45 ;
      RECT MASK 2 34.247 96.21 34.307 96.45 ;
      RECT MASK 2 34.579 96.21 34.639 96.45 ;
      RECT MASK 2 34.911 96.21 34.971 96.45 ;
      RECT MASK 2 35.243 96.21 35.303 96.45 ;
      RECT MASK 2 35.575 96.21 35.635 96.45 ;
      RECT MASK 2 35.907 96.21 35.967 96.45 ;
      RECT MASK 2 36.239 96.21 36.299 96.45 ;
      RECT MASK 2 36.571 96.21 36.631 96.45 ;
      RECT MASK 2 2.338 97.238 2.398 107.61 ;
      RECT MASK 2 2.612 97.238 2.672 107.61 ;
      RECT MASK 2 2.886 97.238 2.946 107.61 ;
      RECT MASK 2 3.16 97.238 3.22 107.61 ;
      RECT MASK 2 3.434 97.238 3.494 107.61 ;
      RECT MASK 2 3.708 97.238 3.768 107.61 ;
      RECT MASK 2 3.982 97.238 4.042 107.61 ;
      RECT MASK 2 4.256 97.238 4.316 107.61 ;
      RECT MASK 2 4.53 97.238 4.59 107.61 ;
      RECT MASK 2 4.804 97.238 4.864 107.61 ;
      RECT MASK 2 5.078 97.238 5.138 107.61 ;
      RECT MASK 2 5.352 97.238 5.412 107.61 ;
      RECT MASK 2 5.626 97.238 5.686 107.61 ;
      RECT MASK 2 5.9 97.238 5.96 107.61 ;
      RECT MASK 2 6.174 97.238 6.234 107.61 ;
      RECT MASK 2 6.448 97.238 6.508 107.61 ;
      RECT MASK 2 6.722 97.238 6.782 107.61 ;
      RECT MASK 2 6.996 97.238 7.056 107.61 ;
      RECT MASK 2 7.27 97.238 7.33 107.61 ;
      RECT MASK 2 7.544 97.238 7.604 107.61 ;
      RECT MASK 2 7.818 97.238 7.878 107.61 ;
      RECT MASK 2 8.092 97.238 8.152 107.61 ;
      RECT MASK 2 8.366 97.238 8.426 107.61 ;
      RECT MASK 2 8.64 97.238 8.7 107.61 ;
      RECT MASK 2 8.914 97.238 8.974 107.61 ;
      RECT MASK 2 9.188 97.238 9.248 107.61 ;
      RECT MASK 2 9.462 97.238 9.522 107.61 ;
      RECT MASK 2 9.736 97.238 9.796 107.61 ;
      RECT MASK 2 10.01 97.238 10.07 107.61 ;
      RECT MASK 2 10.284 97.238 10.344 107.61 ;
      RECT MASK 2 10.558 97.238 10.618 107.61 ;
      RECT MASK 2 10.832 97.238 10.892 107.61 ;
      RECT MASK 2 11.106 97.238 11.166 107.61 ;
      RECT MASK 2 11.38 97.238 11.44 107.61 ;
      RECT MASK 2 11.654 97.238 11.714 107.61 ;
      RECT MASK 2 11.928 97.238 11.988 107.61 ;
      RECT MASK 2 12.202 97.238 12.262 107.61 ;
      RECT MASK 2 12.476 97.238 12.536 107.61 ;
      RECT MASK 2 12.75 97.238 12.81 107.61 ;
      RECT MASK 2 13.024 97.238 13.084 107.61 ;
      RECT MASK 2 13.298 97.238 13.358 107.61 ;
      RECT MASK 2 13.572 97.238 13.632 107.61 ;
      RECT MASK 2 13.846 97.238 13.906 107.61 ;
      RECT MASK 2 14.12 97.238 14.18 107.61 ;
      RECT MASK 2 14.394 97.238 14.454 107.61 ;
      RECT MASK 2 14.668 97.238 14.728 107.61 ;
      RECT MASK 2 14.942 97.238 15.002 107.61 ;
      RECT MASK 2 15.216 97.238 15.276 107.61 ;
      RECT MASK 2 15.49 97.238 15.55 107.61 ;
      RECT MASK 2 15.764 97.238 15.824 107.61 ;
      RECT MASK 2 16.038 97.238 16.098 107.61 ;
      RECT MASK 2 16.312 97.238 16.372 107.61 ;
      RECT MASK 2 16.586 97.238 16.646 107.61 ;
      RECT MASK 2 16.86 97.238 16.92 107.61 ;
      RECT MASK 2 17.134 97.238 17.194 107.61 ;
      RECT MASK 2 17.408 97.238 17.468 107.61 ;
      RECT MASK 2 17.682 97.238 17.742 107.61 ;
      RECT MASK 2 17.956 97.238 18.016 107.61 ;
      RECT MASK 2 18.23 97.238 18.29 107.61 ;
      RECT MASK 2 18.504 97.238 18.564 107.61 ;
      RECT MASK 2 18.778 97.238 18.838 107.61 ;
      RECT MASK 2 19.052 97.238 19.112 107.61 ;
      RECT MASK 2 19.326 97.238 19.386 107.61 ;
      RECT MASK 2 19.6 97.238 19.66 107.61 ;
      RECT MASK 2 19.874 97.238 19.934 107.61 ;
      RECT MASK 2 20.148 97.238 20.208 107.61 ;
      RECT MASK 2 20.422 97.238 20.482 107.61 ;
      RECT MASK 2 20.696 97.238 20.756 107.61 ;
      RECT MASK 2 20.97 97.238 21.03 107.61 ;
      RECT MASK 2 21.244 97.238 21.304 107.61 ;
      RECT MASK 2 21.518 97.238 21.578 107.61 ;
      RECT MASK 2 21.792 97.238 21.852 107.61 ;
      RECT MASK 2 22.066 97.238 22.126 107.61 ;
      RECT MASK 2 22.34 97.238 22.4 107.61 ;
      RECT MASK 2 22.614 97.238 22.674 107.61 ;
      RECT MASK 2 22.888 97.238 22.948 107.61 ;
      RECT MASK 2 23.162 97.238 23.222 107.61 ;
      RECT MASK 2 23.436 97.238 23.496 107.61 ;
      RECT MASK 2 23.71 97.238 23.77 107.61 ;
      RECT MASK 2 23.984 97.238 24.044 107.61 ;
      RECT MASK 2 24.258 97.238 24.318 107.61 ;
      RECT MASK 2 24.532 97.238 24.592 107.61 ;
      RECT MASK 2 24.806 97.238 24.866 107.61 ;
      RECT MASK 2 25.08 97.238 25.14 107.61 ;
      RECT MASK 2 25.354 97.238 25.414 107.61 ;
      RECT MASK 2 25.628 97.238 25.688 107.61 ;
      RECT MASK 2 25.902 97.238 25.962 107.61 ;
      RECT MASK 2 26.176 97.238 26.236 107.61 ;
      RECT MASK 2 26.45 97.238 26.51 107.61 ;
      RECT MASK 2 26.724 97.238 26.784 107.61 ;
      RECT MASK 2 26.998 97.238 27.058 107.61 ;
      RECT MASK 2 27.272 97.238 27.332 107.61 ;
      RECT MASK 2 27.546 97.238 27.606 107.61 ;
      RECT MASK 2 27.82 97.238 27.88 107.61 ;
      RECT MASK 2 28.094 97.238 28.154 107.61 ;
      RECT MASK 2 28.368 97.238 28.428 107.61 ;
      RECT MASK 2 28.642 97.238 28.702 107.61 ;
      RECT MASK 2 28.916 97.238 28.976 107.61 ;
      RECT MASK 2 29.19 97.238 29.25 107.61 ;
      RECT MASK 2 29.464 97.238 29.524 107.61 ;
      RECT MASK 2 29.738 97.238 29.798 107.61 ;
      RECT MASK 2 30.012 97.238 30.072 107.61 ;
      RECT MASK 2 30.286 97.238 30.346 107.61 ;
      RECT MASK 2 30.56 97.238 30.62 107.61 ;
      RECT MASK 2 30.834 97.238 30.894 107.61 ;
      RECT MASK 2 31.108 97.238 31.168 107.61 ;
      RECT MASK 2 31.382 97.238 31.442 107.61 ;
      RECT MASK 2 31.656 97.238 31.716 107.61 ;
      RECT MASK 2 31.93 97.238 31.99 107.61 ;
      RECT MASK 2 32.204 97.238 32.264 107.61 ;
      RECT MASK 2 32.478 97.238 32.538 107.61 ;
      RECT MASK 2 32.752 97.238 32.812 107.61 ;
      RECT MASK 2 33.026 97.238 33.086 107.61 ;
      RECT MASK 2 33.3 97.238 33.36 107.61 ;
      RECT MASK 2 33.574 97.238 33.634 107.61 ;
      RECT MASK 2 33.848 97.238 33.908 107.61 ;
      RECT MASK 2 34.122 97.238 34.182 107.61 ;
      RECT MASK 2 34.396 97.238 34.456 107.61 ;
      RECT MASK 2 34.67 97.238 34.73 107.61 ;
      RECT MASK 2 34.944 97.238 35.004 107.61 ;
      RECT MASK 2 35.218 97.238 35.278 107.61 ;
      RECT MASK 2 35.492 97.238 35.552 107.61 ;
      RECT MASK 2 35.766 97.238 35.826 107.61 ;
      RECT MASK 2 36.04 97.238 36.1 107.61 ;
      RECT MASK 2 36.314 97.238 36.374 107.61 ;
      RECT MASK 2 36.588 97.238 36.648 107.61 ;
      RECT MASK 2 36.862 97.238 36.922 107.61 ;
      RECT MASK 2 37.136 97.238 37.196 107.61 ;
      RECT MASK 2 37.41 97.238 37.47 107.61 ;
      RECT MASK 2 37.684 97.238 37.744 107.61 ;
      RECT MASK 2 37.958 97.238 38.018 107.61 ;
      RECT MASK 2 38.232 97.238 38.292 107.61 ;
      RECT MASK 2 38.506 97.238 38.566 107.61 ;
      RECT MASK 2 38.78 97.238 38.84 107.61 ;
      RECT MASK 2 39.054 97.238 39.114 107.61 ;
      RECT MASK 2 39.328 97.238 39.388 107.61 ;
      RECT MASK 2 39.602 97.238 39.662 107.61 ;
      RECT MASK 2 39.876 97.238 39.936 107.61 ;
      RECT MASK 2 40.15 97.238 40.21 107.61 ;
      RECT MASK 2 40.424 97.238 40.484 107.61 ;
      RECT MASK 2 40.698 97.238 40.758 107.61 ;
      RECT MASK 2 40.972 97.238 41.032 107.61 ;
      RECT MASK 2 41.246 97.238 41.306 107.61 ;
      RECT MASK 2 41.52 97.238 41.58 107.61 ;
      RECT MASK 2 41.794 97.238 41.854 107.61 ;
      RECT MASK 2 42.068 97.238 42.128 107.61 ;
      RECT MASK 2 42.342 97.238 42.402 107.61 ;
      RECT MASK 2 42.616 97.238 42.676 107.61 ;
      RECT MASK 2 42.89 97.238 42.95 107.61 ;
      RECT MASK 2 43.164 97.238 43.224 107.61 ;
      RECT MASK 2 43.438 97.238 43.498 107.61 ;
      RECT MASK 2 45.73 97.238 45.79 107.61 ;
      RECT MASK 2 46.004 97.238 46.064 107.61 ;
      RECT MASK 2 46.278 97.238 46.338 107.61 ;
      RECT MASK 2 46.552 97.238 46.612 107.61 ;
      RECT MASK 2 46.826 97.238 46.886 107.61 ;
      RECT MASK 2 47.1 97.238 47.16 107.61 ;
      RECT MASK 2 47.374 97.238 47.434 107.61 ;
      RECT MASK 2 47.648 97.238 47.708 107.61 ;
      RECT MASK 2 47.922 97.238 47.982 107.61 ;
      RECT MASK 2 48.196 97.238 48.256 107.61 ;
      RECT MASK 2 48.47 97.238 48.53 107.61 ;
      RECT MASK 2 48.744 97.238 48.804 107.61 ;
      RECT MASK 2 49.018 97.238 49.078 107.61 ;
      RECT MASK 2 49.292 97.238 49.352 107.61 ;
      RECT MASK 2 49.566 97.238 49.626 107.61 ;
      RECT MASK 2 49.84 97.238 49.9 107.61 ;
      RECT MASK 2 50.114 97.238 50.174 107.61 ;
      RECT MASK 2 50.388 97.238 50.448 107.61 ;
      RECT MASK 2 50.662 97.238 50.722 107.61 ;
      RECT MASK 2 50.936 97.238 50.996 107.61 ;
      RECT MASK 2 51.21 97.238 51.27 107.61 ;
      RECT MASK 2 51.484 97.238 51.544 107.61 ;
      RECT MASK 2 51.758 97.238 51.818 107.61 ;
      RECT MASK 2 52.032 97.238 52.092 107.61 ;
      RECT MASK 2 52.306 97.238 52.366 107.61 ;
      RECT MASK 2 52.58 97.238 52.64 107.61 ;
      RECT MASK 2 52.854 97.238 52.914 107.61 ;
      RECT MASK 2 53.128 97.238 53.188 107.61 ;
      RECT MASK 2 53.402 97.238 53.462 107.61 ;
      RECT MASK 2 53.676 97.238 53.736 107.61 ;
      RECT MASK 2 53.95 97.238 54.01 107.61 ;
      RECT MASK 2 54.224 97.238 54.284 107.61 ;
      RECT MASK 2 54.498 97.238 54.558 107.61 ;
      RECT MASK 2 54.772 97.238 54.832 107.61 ;
      RECT MASK 2 55.046 97.238 55.106 107.61 ;
      RECT MASK 2 55.32 97.238 55.38 107.61 ;
      RECT MASK 2 55.594 97.238 55.654 107.61 ;
      RECT MASK 2 55.868 97.238 55.928 107.61 ;
      RECT MASK 2 56.142 97.238 56.202 107.61 ;
      RECT MASK 2 56.416 97.238 56.476 107.61 ;
      RECT MASK 2 56.69 97.238 56.75 107.61 ;
      RECT MASK 2 56.964 97.238 57.024 107.61 ;
      RECT MASK 2 57.238 97.238 57.298 107.61 ;
      RECT MASK 2 57.512 97.238 57.572 107.61 ;
      RECT MASK 2 57.786 97.238 57.846 107.61 ;
      RECT MASK 2 58.06 97.238 58.12 107.61 ;
      RECT MASK 2 58.334 97.238 58.394 107.61 ;
      RECT MASK 2 58.608 97.238 58.668 107.61 ;
      RECT MASK 2 58.882 97.238 58.942 107.61 ;
      RECT MASK 2 59.156 97.238 59.216 107.61 ;
      RECT MASK 2 59.43 97.238 59.49 107.61 ;
      RECT MASK 2 59.704 97.238 59.764 107.61 ;
      RECT MASK 2 59.978 97.238 60.038 107.61 ;
      RECT MASK 2 60.252 97.238 60.312 107.61 ;
      RECT MASK 2 60.526 97.238 60.586 107.61 ;
      RECT MASK 2 60.8 97.238 60.86 107.61 ;
      RECT MASK 2 61.074 97.238 61.134 107.61 ;
      RECT MASK 2 61.348 97.238 61.408 107.61 ;
      RECT MASK 2 61.622 97.238 61.682 107.61 ;
      RECT MASK 2 61.896 97.238 61.956 107.61 ;
      RECT MASK 2 62.17 97.238 62.23 107.61 ;
      RECT MASK 2 62.444 97.238 62.504 107.61 ;
      RECT MASK 2 62.718 97.238 62.778 107.61 ;
      RECT MASK 2 62.992 97.238 63.052 107.61 ;
      RECT MASK 2 63.266 97.238 63.326 107.61 ;
      RECT MASK 2 63.54 97.238 63.6 107.61 ;
      RECT MASK 2 63.814 97.238 63.874 107.61 ;
      RECT MASK 2 64.088 97.238 64.148 107.61 ;
      RECT MASK 2 64.362 97.238 64.422 107.61 ;
      RECT MASK 2 64.636 97.238 64.696 107.61 ;
      RECT MASK 2 64.91 97.238 64.97 107.61 ;
      RECT MASK 2 65.184 97.238 65.244 107.61 ;
      RECT MASK 2 65.458 97.238 65.518 107.61 ;
      RECT MASK 2 65.732 97.238 65.792 107.61 ;
      RECT MASK 2 66.006 97.238 66.066 107.61 ;
      RECT MASK 2 66.28 97.238 66.34 107.61 ;
      RECT MASK 2 66.554 97.238 66.614 107.61 ;
      RECT MASK 2 66.828 97.238 66.888 107.61 ;
      RECT MASK 2 67.102 97.238 67.162 107.61 ;
      RECT MASK 2 67.376 97.238 67.436 107.61 ;
      RECT MASK 2 67.65 97.238 67.71 107.61 ;
      RECT MASK 2 67.924 97.238 67.984 107.61 ;
      RECT MASK 2 68.198 97.238 68.258 107.61 ;
      RECT MASK 2 68.472 97.238 68.532 107.61 ;
      RECT MASK 2 68.746 97.238 68.806 107.61 ;
      RECT MASK 2 69.02 97.238 69.08 107.61 ;
      RECT MASK 2 69.294 97.238 69.354 107.61 ;
      RECT MASK 2 69.568 97.238 69.628 107.61 ;
      RECT MASK 2 69.842 97.238 69.902 107.61 ;
      RECT MASK 2 70.116 97.238 70.176 107.61 ;
      RECT MASK 2 70.39 97.238 70.45 107.61 ;
      RECT MASK 2 70.664 97.238 70.724 107.61 ;
      RECT MASK 2 70.938 97.238 70.998 107.61 ;
      RECT MASK 2 71.212 97.238 71.272 107.61 ;
      RECT MASK 2 71.486 97.238 71.546 107.61 ;
      RECT MASK 2 71.76 97.238 71.82 107.61 ;
      RECT MASK 2 72.034 97.238 72.094 107.61 ;
      RECT MASK 2 72.308 97.238 72.368 107.61 ;
      RECT MASK 2 72.582 97.238 72.642 107.61 ;
      RECT MASK 2 72.856 97.238 72.916 107.61 ;
      RECT MASK 2 73.13 97.238 73.19 107.61 ;
      RECT MASK 2 73.404 97.238 73.464 107.61 ;
      RECT MASK 2 73.678 97.238 73.738 107.61 ;
      RECT MASK 2 73.952 97.238 74.012 107.61 ;
      RECT MASK 2 74.226 97.238 74.286 107.61 ;
      RECT MASK 2 74.5 97.238 74.56 107.61 ;
      RECT MASK 2 74.774 97.238 74.834 107.61 ;
      RECT MASK 2 75.048 97.238 75.108 107.61 ;
      RECT MASK 2 75.322 97.238 75.382 107.61 ;
      RECT MASK 2 75.596 97.238 75.656 107.61 ;
      RECT MASK 2 75.87 97.238 75.93 107.61 ;
      RECT MASK 2 76.144 97.238 76.204 107.61 ;
      RECT MASK 2 76.418 97.238 76.478 107.61 ;
      RECT MASK 2 76.692 97.238 76.752 107.61 ;
      RECT MASK 2 76.966 97.238 77.026 107.61 ;
      RECT MASK 2 77.24 97.238 77.3 107.61 ;
      RECT MASK 2 77.514 97.238 77.574 107.61 ;
      RECT MASK 2 77.788 97.238 77.848 107.61 ;
      RECT MASK 2 78.062 97.238 78.122 107.61 ;
      RECT MASK 2 78.336 97.238 78.396 107.61 ;
      RECT MASK 2 78.61 97.238 78.67 107.61 ;
      RECT MASK 2 78.884 97.238 78.944 107.61 ;
      RECT MASK 2 79.158 97.238 79.218 107.61 ;
      RECT MASK 2 79.432 97.238 79.492 107.61 ;
      RECT MASK 2 79.706 97.238 79.766 107.61 ;
      RECT MASK 2 79.98 97.238 80.04 107.61 ;
      RECT MASK 2 80.254 97.238 80.314 107.61 ;
      RECT MASK 2 80.528 97.238 80.588 107.61 ;
      RECT MASK 2 80.802 97.238 80.862 107.61 ;
      RECT MASK 2 81.076 97.238 81.136 107.61 ;
      RECT MASK 2 81.35 97.238 81.41 107.61 ;
      RECT MASK 2 81.624 97.238 81.684 107.61 ;
      RECT MASK 2 81.898 97.238 81.958 107.61 ;
      RECT MASK 2 82.172 97.238 82.232 107.61 ;
      RECT MASK 2 82.446 97.238 82.506 107.61 ;
      RECT MASK 2 82.72 97.238 82.78 107.61 ;
      RECT MASK 2 82.994 97.238 83.054 107.61 ;
      RECT MASK 2 83.268 97.238 83.328 107.61 ;
      RECT MASK 2 83.542 97.238 83.602 107.61 ;
      RECT MASK 2 83.816 97.238 83.876 107.61 ;
      RECT MASK 2 84.09 97.238 84.15 107.61 ;
      RECT MASK 2 84.364 97.238 84.424 107.61 ;
      RECT MASK 2 84.638 97.238 84.698 107.61 ;
      RECT MASK 2 84.912 97.238 84.972 107.61 ;
      RECT MASK 2 85.186 97.238 85.246 107.61 ;
      RECT MASK 2 85.46 97.238 85.52 107.61 ;
      RECT MASK 2 85.734 97.238 85.794 107.61 ;
      RECT MASK 2 86.008 97.238 86.068 107.61 ;
      RECT MASK 2 86.282 97.238 86.342 107.61 ;
      RECT MASK 2 86.556 97.238 86.616 107.61 ;
      RECT MASK 2 86.83 97.238 86.89 107.61 ;
      RECT MASK 2 89.089 97.238 89.149 107.61 ;
      RECT MASK 2 89.363 97.238 89.423 107.61 ;
      RECT MASK 2 89.637 97.238 89.697 107.61 ;
      RECT MASK 2 89.911 97.238 89.971 107.61 ;
      RECT MASK 2 90.185 97.238 90.245 107.61 ;
      RECT MASK 2 90.459 97.238 90.519 107.61 ;
      RECT MASK 2 90.733 97.238 90.793 107.61 ;
      RECT MASK 2 91.007 97.238 91.067 107.61 ;
      RECT MASK 2 91.281 97.238 91.341 107.61 ;
      RECT MASK 2 91.555 97.238 91.615 107.61 ;
      RECT MASK 2 91.829 97.238 91.889 107.61 ;
      RECT MASK 2 92.103 97.238 92.163 107.61 ;
      RECT MASK 2 92.377 97.238 92.437 107.61 ;
      RECT MASK 2 92.651 97.238 92.711 107.61 ;
      RECT MASK 2 92.925 97.238 92.985 107.61 ;
      RECT MASK 2 93.199 97.238 93.259 107.61 ;
      RECT MASK 2 93.473 97.238 93.533 107.61 ;
      RECT MASK 2 93.747 97.238 93.807 107.61 ;
      RECT MASK 2 94.021 97.238 94.081 107.61 ;
      RECT MASK 2 94.295 97.238 94.355 107.61 ;
      RECT MASK 2 94.569 97.238 94.629 107.61 ;
      RECT MASK 2 94.843 97.238 94.903 107.61 ;
      RECT MASK 2 95.117 97.238 95.177 107.61 ;
      RECT MASK 2 95.391 97.238 95.451 107.61 ;
      RECT MASK 2 95.665 97.238 95.725 107.61 ;
      RECT MASK 2 95.939 97.238 95.999 107.61 ;
      RECT MASK 2 96.213 97.238 96.273 107.61 ;
      RECT MASK 2 96.487 97.238 96.547 107.61 ;
      RECT MASK 2 96.761 97.238 96.821 107.61 ;
      RECT MASK 2 97.035 97.238 97.095 107.61 ;
      RECT MASK 2 97.309 97.238 97.369 107.61 ;
      RECT MASK 2 97.583 97.238 97.643 107.61 ;
      RECT MASK 2 97.857 97.238 97.917 107.61 ;
      RECT MASK 2 98.131 97.238 98.191 107.61 ;
      RECT MASK 2 98.405 97.238 98.465 107.61 ;
      RECT MASK 2 98.679 97.238 98.739 107.61 ;
      RECT MASK 2 98.953 97.238 99.013 107.61 ;
      RECT MASK 2 99.227 97.238 99.287 107.61 ;
      RECT MASK 2 99.501 97.238 99.561 107.61 ;
      RECT MASK 2 99.775 97.238 99.835 107.61 ;
      RECT MASK 2 100.049 97.238 100.109 107.61 ;
      RECT MASK 2 100.323 97.238 100.383 107.61 ;
      RECT MASK 2 100.597 97.238 100.657 107.61 ;
      RECT MASK 2 100.871 97.238 100.931 107.61 ;
      RECT MASK 2 101.145 97.238 101.205 107.61 ;
      RECT MASK 2 101.419 97.238 101.479 107.61 ;
      RECT MASK 2 101.693 97.238 101.753 107.61 ;
      RECT MASK 2 101.967 97.238 102.027 107.61 ;
      RECT MASK 2 102.241 97.238 102.301 107.61 ;
      RECT MASK 2 102.515 97.238 102.575 107.61 ;
      RECT MASK 2 102.789 97.238 102.849 107.61 ;
      RECT MASK 2 103.063 97.238 103.123 107.61 ;
      RECT MASK 2 103.337 97.238 103.397 107.61 ;
      RECT MASK 2 103.611 97.238 103.671 107.61 ;
      RECT MASK 2 103.885 97.238 103.945 107.61 ;
      RECT MASK 2 104.159 97.238 104.219 107.61 ;
      RECT MASK 2 104.433 97.238 104.493 107.61 ;
      RECT MASK 2 104.707 97.238 104.767 107.61 ;
      RECT MASK 2 104.981 97.238 105.041 107.61 ;
      RECT MASK 2 105.255 97.238 105.315 107.61 ;
      RECT MASK 2 105.529 97.238 105.589 107.61 ;
      RECT MASK 2 105.803 97.238 105.863 107.61 ;
      RECT MASK 2 106.077 97.238 106.137 107.61 ;
      RECT MASK 2 106.351 97.238 106.411 107.61 ;
      RECT MASK 2 106.625 97.238 106.685 107.61 ;
      RECT MASK 2 106.899 97.238 106.959 107.61 ;
      RECT MASK 2 107.173 97.238 107.233 107.61 ;
      RECT MASK 2 107.447 97.238 107.507 107.61 ;
      RECT MASK 2 107.721 97.238 107.781 107.61 ;
      RECT MASK 2 107.995 97.238 108.055 107.61 ;
      RECT MASK 2 108.269 97.238 108.329 107.61 ;
      RECT MASK 2 108.543 97.238 108.603 107.61 ;
      RECT MASK 2 108.817 97.238 108.877 107.61 ;
      RECT MASK 2 109.091 97.238 109.151 107.61 ;
      RECT MASK 2 109.365 97.238 109.425 107.61 ;
      RECT MASK 2 109.639 97.238 109.699 107.61 ;
      RECT MASK 2 109.913 97.238 109.973 107.61 ;
      RECT MASK 2 110.187 97.238 110.247 107.61 ;
      RECT MASK 2 110.461 97.238 110.521 107.61 ;
      RECT MASK 2 110.735 97.238 110.795 107.61 ;
      RECT MASK 2 111.009 97.238 111.069 107.61 ;
      RECT MASK 2 111.283 97.238 111.343 107.61 ;
      RECT MASK 2 111.557 97.238 111.617 107.61 ;
      RECT MASK 2 111.831 97.238 111.891 107.61 ;
      RECT MASK 2 112.105 97.238 112.165 107.61 ;
      RECT MASK 2 112.379 97.238 112.439 107.61 ;
      RECT MASK 2 112.653 97.238 112.713 107.61 ;
      RECT MASK 2 112.927 97.238 112.987 107.61 ;
      RECT MASK 2 113.201 97.238 113.261 107.61 ;
      RECT MASK 2 113.475 97.238 113.535 107.61 ;
      RECT MASK 2 113.749 97.238 113.809 107.61 ;
      RECT MASK 2 114.023 97.238 114.083 107.61 ;
      RECT MASK 2 114.297 97.238 114.357 107.61 ;
      RECT MASK 2 114.571 97.238 114.631 107.61 ;
      RECT MASK 2 114.845 97.238 114.905 107.61 ;
      RECT MASK 2 115.119 97.238 115.179 107.61 ;
      RECT MASK 2 115.393 97.238 115.453 107.61 ;
      RECT MASK 2 115.667 97.238 115.727 107.61 ;
      RECT MASK 2 115.941 97.238 116.001 107.61 ;
      RECT MASK 2 116.215 97.238 116.275 107.61 ;
      RECT MASK 2 116.489 97.238 116.549 107.61 ;
      RECT MASK 2 116.763 97.238 116.823 107.61 ;
      RECT MASK 2 117.037 97.238 117.097 107.61 ;
      RECT MASK 2 117.311 97.238 117.371 107.61 ;
      RECT MASK 2 117.585 97.238 117.645 107.61 ;
      RECT MASK 2 117.859 97.238 117.919 107.61 ;
      RECT MASK 2 118.133 97.238 118.193 107.61 ;
      RECT MASK 2 118.407 97.238 118.467 107.61 ;
      RECT MASK 2 118.681 97.238 118.741 107.61 ;
      RECT MASK 2 118.955 97.238 119.015 107.61 ;
      RECT MASK 2 119.229 97.238 119.289 107.61 ;
      RECT MASK 2 119.503 97.238 119.563 107.61 ;
      RECT MASK 2 119.777 97.238 119.837 107.61 ;
      RECT MASK 2 120.051 97.238 120.111 107.61 ;
      RECT MASK 2 120.325 97.238 120.385 107.61 ;
      RECT MASK 2 120.599 97.238 120.659 107.61 ;
      RECT MASK 2 120.873 97.238 120.933 107.61 ;
      RECT MASK 2 121.147 97.238 121.207 107.61 ;
      RECT MASK 2 121.421 97.238 121.481 107.61 ;
      RECT MASK 2 121.695 97.238 121.755 107.61 ;
      RECT MASK 2 121.969 97.238 122.029 107.61 ;
      RECT MASK 2 122.243 97.238 122.303 107.61 ;
      RECT MASK 2 122.517 97.238 122.577 107.61 ;
      RECT MASK 2 122.791 97.238 122.851 107.61 ;
      RECT MASK 2 123.065 97.238 123.125 107.61 ;
      RECT MASK 2 123.339 97.238 123.399 107.61 ;
      RECT MASK 2 123.613 97.238 123.673 107.61 ;
      RECT MASK 2 123.887 97.238 123.947 107.61 ;
      RECT MASK 2 124.161 97.238 124.221 107.61 ;
      RECT MASK 2 124.435 97.238 124.495 107.61 ;
      RECT MASK 2 124.709 97.238 124.769 107.61 ;
      RECT MASK 2 124.983 97.238 125.043 107.61 ;
      RECT MASK 2 125.257 97.238 125.317 107.61 ;
      RECT MASK 2 125.531 97.238 125.591 107.61 ;
      RECT MASK 2 125.805 97.238 125.865 107.61 ;
      RECT MASK 2 126.079 97.238 126.139 107.61 ;
      RECT MASK 2 126.353 97.238 126.413 107.61 ;
      RECT MASK 2 126.627 97.238 126.687 107.61 ;
      RECT MASK 2 126.901 97.238 126.961 107.61 ;
      RECT MASK 2 127.175 97.238 127.235 107.61 ;
      RECT MASK 2 127.449 97.238 127.509 107.61 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 1 22.6135 0.75 46.3385 0.79 ;
      RECT MASK 1 24.0135 0.95 48.496 0.99 ;
      RECT MASK 1 22.175 1.15 45.8385 1.19 ;
      RECT MASK 1 58.969 1.18 65.033 1.22 ;
      RECT MASK 1 61.03 1.42 63.793 1.46 ;
      RECT MASK 1 49.934 1.45 52.6425 1.49 ;
      RECT MASK 1 3.1975 1.5515 43.5385 1.5915 ;
      RECT MASK 1 58.74 1.66 59.766 1.7 ;
      RECT MASK 1 61.259 1.66 61.827 1.7 ;
      RECT MASK 1 62.175 1.66 62.743 1.7 ;
      RECT MASK 1 63.708 1.66 63.919 1.7 ;
      RECT MASK 1 64.599 1.66 64.842 1.7 ;
      RECT MASK 1 116.256 1.78 128.056 1.82 ;
      RECT MASK 1 49.9865 1.9 52.6425 1.94 ;
      RECT MASK 1 61.488 1.9 63.793 1.94 ;
      RECT MASK 1 46.106 1.97 49.1005 2.05 ;
      RECT MASK 1 116.256 2.02 128.056 2.06 ;
      RECT MASK 1 21.633 2.07 25.304 2.15 ;
      RECT MASK 1 6.2185 2.11 21.2995 2.15 ;
      RECT MASK 1 25.6375 2.11 40.7185 2.15 ;
      RECT MASK 1 57.536 2.14 60.453 2.18 ;
      RECT MASK 1 63.778 2.14 66.237 2.18 ;
      RECT MASK 1 116.256 2.26 128.056 2.3 ;
      RECT MASK 1 45.697 2.29 47.0605 2.33 ;
      RECT MASK 1 3.8695 2.35 7.1295 2.39 ;
      RECT MASK 1 8.4845 2.35 9.1875 2.39 ;
      RECT MASK 1 10.7775 2.35 11.7125 2.39 ;
      RECT MASK 1 35.2245 2.35 36.1595 2.39 ;
      RECT MASK 1 37.7495 2.35 38.4525 2.39 ;
      RECT MASK 1 39.8075 2.35 43.0675 2.39 ;
      RECT MASK 1 57.536 2.43 66.237 2.61 ;
      RECT MASK 1 49.9865 2.48 52.6425 2.52 ;
      RECT MASK 1 116.256 2.5 128.056 2.54 ;
      RECT MASK 1 3.1975 2.59 3.5085 2.63 ;
      RECT MASK 1 3.8695 2.59 9.8545 2.63 ;
      RECT MASK 1 10.0225 2.59 22.5235 2.63 ;
      RECT MASK 1 22.949 2.59 23.454 2.63 ;
      RECT MASK 1 23.7135 2.59 24.179 2.63 ;
      RECT MASK 1 24.4135 2.59 36.9145 2.63 ;
      RECT MASK 1 37.0825 2.59 43.0675 2.63 ;
      RECT MASK 1 43.3585 2.59 43.653 2.63 ;
      RECT MASK 1 116.256 2.74 128.056 2.78 ;
      RECT MASK 1 4.4395 2.83 5.0075 2.87 ;
      RECT MASK 1 7.1225 2.83 8.0295 2.87 ;
      RECT MASK 1 38.9075 2.83 39.8145 2.87 ;
      RECT MASK 1 41.9295 2.83 42.4975 2.87 ;
      RECT MASK 1 57.536 2.86 66.237 2.9 ;
      RECT MASK 1 116.256 2.98 128.056 3.02 ;
      RECT MASK 1 22.0175 3.03 24.8685 3.11 ;
      RECT MASK 1 47.543 3.03 48.2475 3.07 ;
      RECT MASK 1 1.3865 3.07 13.7315 3.11 ;
      RECT MASK 1 14.2605 3.07 21.7575 3.11 ;
      RECT MASK 1 25.1795 3.07 32.6765 3.11 ;
      RECT MASK 1 33.2055 3.07 45.5505 3.11 ;
      RECT MASK 1 60.029 3.1 65.491 3.14 ;
      RECT MASK 1 47.115 3.19 47.4605 3.23 ;
      RECT MASK 1 116.256 3.22 128.056 3.26 ;
      RECT MASK 1 62.2375 3.34 62.9075 3.38 ;
      RECT MASK 1 63.535 3.34 65.033 3.38 ;
      RECT MASK 1 56.3455 3.3585 59.444 3.3985 ;
      RECT MASK 1 1.3865 3.36 13.7315 3.54 ;
      RECT MASK 1 14.3195 3.36 21.7575 3.54 ;
      RECT MASK 1 22.0685 3.36 24.8685 3.54 ;
      RECT MASK 1 25.1795 3.36 32.6175 3.54 ;
      RECT MASK 1 33.2055 3.36 45.5505 3.54 ;
      RECT MASK 1 45.9035 3.41 49.1005 3.49 ;
      RECT MASK 1 116.256 3.46 128.056 3.5 ;
      RECT MASK 1 62.235 3.578 66.703 3.618 ;
      RECT MASK 1 47.9205 3.67 49.497 3.71 ;
      RECT MASK 1 116.256 3.7 128.056 3.74 ;
      RECT MASK 1 59.147 3.82 59.308 3.86 ;
      RECT MASK 1 59.656 3.82 60.139 3.86 ;
      RECT MASK 1 63.778 3.82 64.346 3.86 ;
      RECT MASK 1 64.694 3.82 65.262 3.86 ;
      RECT MASK 1 46.943 3.83 47.4155 3.87 ;
      RECT MASK 1 47.5755 3.83 48.2565 3.87 ;
      RECT MASK 1 1.3865 3.84 13.7315 4.02 ;
      RECT MASK 1 14.3195 3.84 21.7575 4.02 ;
      RECT MASK 1 22.0175 3.84 24.8685 4.02 ;
      RECT MASK 1 25.1795 3.84 32.6175 4.02 ;
      RECT MASK 1 33.2055 3.84 45.5505 4.02 ;
      RECT MASK 1 116.256 3.94 128.056 3.98 ;
      RECT MASK 1 116.256 4.18 128.056 4.22 ;
      RECT MASK 1 1.3865 4.27 13.7315 4.31 ;
      RECT MASK 1 14.2605 4.27 21.7575 4.31 ;
      RECT MASK 1 22.0175 4.27 24.8685 4.35 ;
      RECT MASK 1 25.1795 4.27 32.6765 4.31 ;
      RECT MASK 1 33.2055 4.27 45.5505 4.31 ;
      RECT MASK 1 59.147 4.3 59.308 4.34 ;
      RECT MASK 1 59.656 4.3 60.139 4.34 ;
      RECT MASK 1 63.778 4.3 64.346 4.34 ;
      RECT MASK 1 64.694 4.3 65.262 4.34 ;
      RECT MASK 1 116.256 4.42 128.056 4.46 ;
      RECT MASK 1 4.4395 4.51 5.6525 4.55 ;
      RECT MASK 1 7.1225 4.51 8.0295 4.55 ;
      RECT MASK 1 38.9075 4.51 39.8145 4.55 ;
      RECT MASK 1 41.9295 4.51 42.4975 4.55 ;
      RECT MASK 1 56.536 4.538 67.016 4.578 ;
      RECT MASK 1 116.256 4.66 128.056 4.7 ;
      RECT MASK 1 22.7685 4.738 23.0685 4.778 ;
      RECT MASK 1 3.1975 4.75 3.5085 4.79 ;
      RECT MASK 1 3.8695 4.75 9.8545 4.79 ;
      RECT MASK 1 10.0225 4.75 22.5235 4.79 ;
      RECT MASK 1 23.6775 4.75 24.1705 4.79 ;
      RECT MASK 1 24.4135 4.75 36.9145 4.79 ;
      RECT MASK 1 37.0825 4.75 43.0675 4.79 ;
      RECT MASK 1 43.3585 4.75 43.653 4.79 ;
      RECT MASK 1 80.052 4.765 92.2115 5.015 ;
      RECT MASK 1 94.4935 4.765 106.653 5.015 ;
      RECT MASK 1 56.9885 4.777 59.4465 4.817 ;
      RECT MASK 1 62.578 4.78 63.068 4.82 ;
      RECT MASK 1 63.535 4.78 65.033 4.82 ;
      RECT MASK 1 116.256 4.9 128.056 4.94 ;
      RECT MASK 1 3.8695 4.99 7.1295 5.03 ;
      RECT MASK 1 8.4845 4.99 9.1875 5.03 ;
      RECT MASK 1 10.7775 4.99 11.7125 5.03 ;
      RECT MASK 1 35.2245 4.99 36.1595 5.03 ;
      RECT MASK 1 37.7495 4.99 38.4525 5.03 ;
      RECT MASK 1 39.8075 4.99 43.0675 5.03 ;
      RECT MASK 1 60.029 5.02 65.491 5.06 ;
      RECT MASK 1 116.256 5.14 128.056 5.18 ;
      RECT MASK 1 6.2185 5.23 21.2995 5.27 ;
      RECT MASK 1 21.633 5.23 25.304 5.31 ;
      RECT MASK 1 25.6375 5.23 40.7185 5.27 ;
      RECT MASK 1 57.536 5.26 66.237 5.3 ;
      RECT MASK 1 49.3195 5.316 57.138 5.356 ;
      RECT MASK 1 116.256 5.38 128.056 5.42 ;
      RECT MASK 1 49.9515 5.49 52.6775 5.55 ;
      RECT MASK 1 57.536 5.55 66.237 5.73 ;
      RECT MASK 1 66.825 5.6025 90.887 5.6425 ;
      RECT MASK 1 116.256 5.62 128.056 5.66 ;
      RECT MASK 1 116.256 5.86 128.056 5.9 ;
      RECT MASK 1 49.9515 5.97 52.6775 6.03 ;
      RECT MASK 1 46.9405 5.974 47.5485 6.014 ;
      RECT MASK 1 57.536 5.98 60.453 6.02 ;
      RECT MASK 1 63.778 5.98 66.237 6.02 ;
      RECT MASK 1 116.256 6.1 128.056 6.14 ;
      RECT MASK 1 21.633 6.15 25.304 6.23 ;
      RECT MASK 1 6.2185 6.19 21.2995 6.23 ;
      RECT MASK 1 25.6375 6.19 40.7185 6.23 ;
      RECT MASK 1 53.22 6.22 54.5955 6.26 ;
      RECT MASK 1 61.488 6.22 63.793 6.26 ;
      RECT MASK 1 84.541 6.26 88.641 6.4 ;
      RECT MASK 1 89.568 6.26 90.286 6.4 ;
      RECT MASK 1 96.419 6.26 97.137 6.4 ;
      RECT MASK 1 98.064 6.26 102.164 6.4 ;
      RECT MASK 1 90.73 6.31 91.2585 6.35 ;
      RECT MASK 1 116.256 6.34 128.056 6.38 ;
      RECT MASK 1 46.2625 6.358 47.2165 6.398 ;
      RECT MASK 1 52.874 6.412 54.9405 6.452 ;
      RECT MASK 1 55.1495 6.417 56.677 6.457 ;
      RECT MASK 1 3.8695 6.43 7.1295 6.47 ;
      RECT MASK 1 8.4845 6.43 9.1875 6.47 ;
      RECT MASK 1 10.7775 6.43 11.7125 6.47 ;
      RECT MASK 1 35.2245 6.43 36.1595 6.47 ;
      RECT MASK 1 37.7495 6.43 38.4525 6.47 ;
      RECT MASK 1 39.8075 6.43 43.0675 6.47 ;
      RECT MASK 1 49.9515 6.45 52.6775 6.51 ;
      RECT MASK 1 58.74 6.46 59.766 6.5 ;
      RECT MASK 1 61.259 6.46 61.827 6.5 ;
      RECT MASK 1 62.175 6.46 62.743 6.5 ;
      RECT MASK 1 63.708 6.46 63.919 6.5 ;
      RECT MASK 1 64.599 6.46 64.842 6.5 ;
      RECT MASK 1 116.256 6.58 128.056 6.62 ;
      RECT MASK 1 46.1345 6.648 49.0705 6.828 ;
      RECT MASK 1 3.1975 6.67 3.5085 6.71 ;
      RECT MASK 1 3.8695 6.67 9.8545 6.71 ;
      RECT MASK 1 10.0225 6.67 22.5235 6.71 ;
      RECT MASK 1 24.4135 6.67 36.9145 6.71 ;
      RECT MASK 1 37.0825 6.67 43.0675 6.71 ;
      RECT MASK 1 43.3585 6.67 43.653 6.71 ;
      RECT MASK 1 61.03 6.7 63.793 6.74 ;
      RECT MASK 1 84.5045 6.74 90.939 6.88 ;
      RECT MASK 1 95.766 6.74 102.2005 6.88 ;
      RECT MASK 1 53.499 6.768 56.3975 6.948 ;
      RECT MASK 1 116.256 6.82 128.056 6.86 ;
      RECT MASK 1 4.4395 6.91 5.262 6.95 ;
      RECT MASK 1 7.1225 6.91 8.0295 6.95 ;
      RECT MASK 1 38.9075 6.91 39.8145 6.95 ;
      RECT MASK 1 41.9295 6.91 42.4975 6.95 ;
      RECT MASK 1 58.969 6.94 65.033 6.98 ;
      RECT MASK 1 46.1345 7.032 49.0705 7.212 ;
      RECT MASK 1 116.256 7.06 128.056 7.1 ;
      RECT MASK 1 22.0175 7.11 24.8685 7.19 ;
      RECT MASK 1 1.3865 7.15 13.7315 7.19 ;
      RECT MASK 1 14.2605 7.15 21.7575 7.19 ;
      RECT MASK 1 25.1795 7.15 32.6765 7.19 ;
      RECT MASK 1 33.2055 7.15 45.5505 7.19 ;
      RECT MASK 1 116.256 7.3 128.056 7.34 ;
      RECT MASK 1 50.0625 7.41 50.3535 7.47 ;
      RECT MASK 1 50.7265 7.41 51.0175 7.47 ;
      RECT MASK 1 51.3905 7.41 51.6815 7.47 ;
      RECT MASK 1 52.0545 7.41 52.3455 7.47 ;
      RECT MASK 1 58.969 7.42 65.033 7.46 ;
      RECT MASK 1 1.3865 7.44 13.7315 7.62 ;
      RECT MASK 1 14.3195 7.44 21.7575 7.62 ;
      RECT MASK 1 22.0175 7.44 24.8685 7.62 ;
      RECT MASK 1 25.1795 7.44 32.6175 7.62 ;
      RECT MASK 1 33.2055 7.44 45.5505 7.62 ;
      RECT MASK 1 47.4385 7.467 49.7615 7.507 ;
      RECT MASK 1 116.256 7.54 128.056 7.58 ;
      RECT MASK 1 61.03 7.66 63.793 7.7 ;
      RECT MASK 1 47.072 7.6625 49.5955 7.7025 ;
      RECT MASK 1 116.256 7.78 128.056 7.82 ;
      RECT MASK 1 48.055 7.8815 49.2635 7.9215 ;
      RECT MASK 1 50.2835 7.89 50.5795 7.95 ;
      RECT MASK 1 50.9475 7.89 51.2435 7.95 ;
      RECT MASK 1 51.6115 7.89 51.9075 7.95 ;
      RECT MASK 1 52.2755 7.89 52.5715 7.95 ;
      RECT MASK 1 58.74 7.9 59.766 7.94 ;
      RECT MASK 1 61.259 7.9 61.827 7.94 ;
      RECT MASK 1 62.175 7.9 62.743 7.94 ;
      RECT MASK 1 63.708 7.9 63.919 7.94 ;
      RECT MASK 1 64.599 7.9 64.842 7.94 ;
      RECT MASK 1 116.256 8.02 128.056 8.06 ;
      RECT MASK 1 61.488 8.14 63.793 8.18 ;
      RECT MASK 1 35.8005 8.228 42.0895 8.268 ;
      RECT MASK 1 116.256 8.26 128.056 8.3 ;
      RECT MASK 1 1.3865 8.34 13.7315 8.52 ;
      RECT MASK 1 14.3195 8.34 21.7575 8.52 ;
      RECT MASK 1 22.0175 8.34 23.773 8.52 ;
      RECT MASK 1 49.9515 8.37 52.6775 8.43 ;
      RECT MASK 1 57.536 8.38 60.453 8.42 ;
      RECT MASK 1 63.778 8.38 66.237 8.42 ;
      RECT MASK 1 116.256 8.5 128.056 8.54 ;
      RECT MASK 1 57.536 8.67 66.237 8.85 ;
      RECT MASK 1 116.256 8.74 128.056 8.78 ;
      RECT MASK 1 1.3865 8.77 13.7315 8.81 ;
      RECT MASK 1 14.2605 8.77 21.7575 8.81 ;
      RECT MASK 1 22.0175 8.77 23.485 8.85 ;
      RECT MASK 1 52.867 8.7935 55.3905 8.8335 ;
      RECT MASK 1 49.477 8.81 51.1335 8.85 ;
      RECT MASK 1 49.9515 8.97 52.6775 9.03 ;
      RECT MASK 1 116.256 8.98 128.056 9.02 ;
      RECT MASK 1 3.1975 9.01 3.5085 9.05 ;
      RECT MASK 1 4.3095 9.01 5.0075 9.05 ;
      RECT MASK 1 7.1225 9.01 8.0295 9.05 ;
      RECT MASK 1 44.426 9.0255 47.7145 9.0655 ;
      RECT MASK 1 47.9365 9.0255 48.235 9.0655 ;
      RECT MASK 1 57.536 9.1 66.237 9.14 ;
      RECT MASK 1 69.481 9.194 69.79 9.274 ;
      RECT MASK 1 80.151 9.202 81.6775 9.439 ;
      RECT MASK 1 43.311 9.21 43.644 9.25 ;
      RECT MASK 1 116.256 9.22 128.056 9.26 ;
      RECT MASK 1 47.1065 9.238 51.7975 9.278 ;
      RECT MASK 1 26.357 9.246 33.368 9.286 ;
      RECT MASK 1 36.922 9.246 43.0405 9.286 ;
      RECT MASK 1 3.8695 9.25 9.8545 9.29 ;
      RECT MASK 1 10.0225 9.25 22.5235 9.29 ;
      RECT MASK 1 52.984 9.34 54.9915 9.38 ;
      RECT MASK 1 55.1405 9.34 55.3905 9.38 ;
      RECT MASK 1 60.029 9.34 65.491 9.38 ;
      RECT MASK 1 35.4365 9.443 37.261 9.483 ;
      RECT MASK 1 38.067 9.443 42.4975 9.483 ;
      RECT MASK 1 116.256 9.46 128.056 9.5 ;
      RECT MASK 1 3.8695 9.49 7.1295 9.53 ;
      RECT MASK 1 8.4845 9.49 9.1875 9.53 ;
      RECT MASK 1 10.7775 9.49 11.7125 9.53 ;
      RECT MASK 1 66.667 9.502 68.766 9.542 ;
      RECT MASK 1 68.902 9.502 69.8375 9.542 ;
      RECT MASK 1 46.1345 9.528 49.0705 9.708 ;
      RECT MASK 1 54.1575 9.532 54.8985 9.572 ;
      RECT MASK 1 55.0345 9.532 57.024 9.572 ;
      RECT MASK 1 57.241 9.5765 59.4425 9.6165 ;
      RECT MASK 1 63.535 9.58 65.033 9.62 ;
      RECT MASK 1 31.042 9.615 34.513 9.655 ;
      RECT MASK 1 62.535 9.65 63.079 9.69 ;
      RECT MASK 1 116.256 9.7 128.056 9.74 ;
      RECT MASK 1 6.2185 9.73 21.2995 9.77 ;
      RECT MASK 1 21.633 9.73 23.4685 9.81 ;
      RECT MASK 1 31.393 9.817 32.681 9.857 ;
      RECT MASK 1 36.006 9.818 41.241 9.858 ;
      RECT MASK 1 56.914 9.8205 66.2065 9.8605 ;
      RECT MASK 1 116.256 9.94 128.056 9.98 ;
      RECT MASK 1 67.346 10.008 71.009 10.188 ;
      RECT MASK 1 31.3665 10.038 39.3815 10.218 ;
      RECT MASK 1 53.499 10.038 56.4545 10.218 ;
      RECT MASK 1 59.147 10.06 59.308 10.1 ;
      RECT MASK 1 59.656 10.06 60.139 10.1 ;
      RECT MASK 1 63.778 10.06 64.346 10.1 ;
      RECT MASK 1 64.694 10.06 65.262 10.1 ;
      RECT MASK 1 116.256 10.18 128.056 10.22 ;
      RECT MASK 1 43.2725 10.198 52.998 10.238 ;
      RECT MASK 1 5.4865 10.405 31.028 10.445 ;
      RECT MASK 1 116.256 10.42 128.056 10.46 ;
      RECT MASK 1 43.442 10.49 66.829 10.53 ;
      RECT MASK 1 4.72 10.607 31.3495 10.647 ;
      RECT MASK 1 116.256 10.66 128.056 10.7 ;
      RECT MASK 1 31.719 10.79 53.094 10.83 ;
      RECT MASK 1 116.256 10.9 128.056 10.94 ;
      RECT MASK 1 23.348 10.96 31.8905 11 ;
      RECT MASK 1 42.9305 10.982 59.999 11.022 ;
      RECT MASK 1 24.95 11.174 52.977 11.214 ;
      RECT MASK 1 56.0535 11.174 127.253 11.214 ;
      RECT MASK 1 10.587 11.366 102.163 11.406 ;
      RECT MASK 1 24.697 11.558 91.373 11.598 ;
      RECT MASK 1 4.251 11.78 111.8115 11.98 ;
      RECT MASK 1 116.256 11.86 128.056 11.9 ;
      RECT MASK 1 116.256 12.1 128.056 12.14 ;
      RECT MASK 1 4.251 12.202 111.819 12.402 ;
      RECT MASK 1 116.256 12.34 128.056 12.38 ;
      RECT MASK 1 116.256 12.58 128.056 12.62 ;
      RECT MASK 1 27.519 12.582 29.289 12.622 ;
      RECT MASK 1 29.946 12.582 84.567 12.622 ;
      RECT MASK 1 90.765 12.582 91.871 12.622 ;
      RECT MASK 1 9.923 12.772 49.873 12.812 ;
      RECT MASK 1 51.091 12.772 72.947 12.812 ;
      RECT MASK 1 116.256 12.82 128.056 12.86 ;
      RECT MASK 1 101.721 12.868 102.495 12.908 ;
      RECT MASK 1 68.023 12.962 68.299 13.002 ;
      RECT MASK 1 8.263 12.964 46.553 13.004 ;
      RECT MASK 1 47.771 12.964 54.853 13.004 ;
      RECT MASK 1 55.739 12.964 64.716 13.004 ;
      RECT MASK 1 66.861 12.964 67.635 13.004 ;
      RECT MASK 1 68.521 12.964 69.295 13.004 ;
      RECT MASK 1 69.517 12.964 69.793 13.004 ;
      RECT MASK 1 70.181 12.964 72.615 13.004 ;
      RECT MASK 1 77.485 12.964 78.591 13.004 ;
      RECT MASK 1 79.145 12.964 80.251 13.004 ;
      RECT MASK 1 83.461 12.964 84.235 13.004 ;
      RECT MASK 1 89.105 12.964 90.211 13.004 ;
      RECT MASK 1 103.381 12.964 104.155 13.004 ;
      RECT MASK 1 116.256 13.06 128.056 13.1 ;
      RECT MASK 1 52.253 13.15 53.691 13.19 ;
      RECT MASK 1 62.493 13.15 63.153 13.19 ;
      RECT MASK 1 8.761 13.156 9.203 13.196 ;
      RECT MASK 1 10.421 13.156 18.997 13.196 ;
      RECT MASK 1 22.373 13.156 29.787 13.196 ;
      RECT MASK 1 32.333 13.156 33.771 13.196 ;
      RECT MASK 1 34.491 13.156 34.933 13.196 ;
      RECT MASK 1 35.577 13.156 43.067 13.196 ;
      RECT MASK 1 43.953 13.156 45.391 13.196 ;
      RECT MASK 1 46.111 13.156 47.051 13.196 ;
      RECT MASK 1 47.2465 13.156 48.711 13.196 ;
      RECT MASK 1 48.8905 13.156 50.371 13.196 ;
      RECT MASK 1 50.5505 13.156 52.031 13.196 ;
      RECT MASK 1 54.5765 13.156 55.683 13.196 ;
      RECT MASK 1 57.067 13.156 57.509 13.196 ;
      RECT MASK 1 58.063 13.156 59.293 13.196 ;
      RECT MASK 1 60.719 13.156 62.157 13.196 ;
      RECT MASK 1 65.367 13.156 65.809 13.196 ;
      RECT MASK 1 67.027 13.156 67.469 13.196 ;
      RECT MASK 1 68.023 13.156 72.283 13.196 ;
      RECT MASK 1 76.323 13.156 78.757 13.196 ;
      RECT MASK 1 78.979 13.156 84.733 13.196 ;
      RECT MASK 1 88.939 13.156 90.377 13.196 ;
      RECT MASK 1 90.599 13.156 98.013 13.196 ;
      RECT MASK 1 103.547 13.16 110.463 13.2 ;
      RECT MASK 1 101.887 13.1675 102.329 13.2075 ;
      RECT MASK 1 116.256 13.3 128.056 13.34 ;
      RECT MASK 1 116.256 13.54 128.056 13.58 ;
      RECT MASK 1 116.256 13.78 128.056 13.82 ;
      RECT MASK 1 116.256 14.02 128.056 14.06 ;
      RECT MASK 1 116.256 14.26 128.056 14.3 ;
      RECT MASK 1 38.156 14.398 41.626 14.438 ;
      RECT MASK 1 57.072 14.398 70.623 14.438 ;
      RECT MASK 1 45.4475 14.404 51.367 14.444 ;
      RECT MASK 1 116.256 14.5 128.056 14.54 ;
      RECT MASK 1 5.275 14.596 109.633 14.636 ;
      RECT MASK 1 116.256 14.74 128.056 14.78 ;
      RECT MASK 1 8.595 14.788 106.892 14.828 ;
      RECT MASK 1 81.801 14.976 82.575 15.016 ;
      RECT MASK 1 108.361 14.976 109.135 15.016 ;
      RECT MASK 1 10.255 14.978 11.527 15.018 ;
      RECT MASK 1 11.744 14.978 12.689 15.018 ;
      RECT MASK 1 13.077 14.978 14.349 15.018 ;
      RECT MASK 1 15.235 14.978 16.009 15.018 ;
      RECT MASK 1 16.895 14.978 17.669 15.018 ;
      RECT MASK 1 23.535 14.978 24.309 15.018 ;
      RECT MASK 1 25.195 14.978 25.969 15.018 ;
      RECT MASK 1 26.855 14.978 27.629 15.018 ;
      RECT MASK 1 28.515 14.978 29.289 15.018 ;
      RECT MASK 1 30.175 14.978 30.949 15.018 ;
      RECT MASK 1 36.815 14.978 37.589 15.018 ;
      RECT MASK 1 38.475 14.978 39.249 15.018 ;
      RECT MASK 1 40.135 14.978 40.909 15.018 ;
      RECT MASK 1 41.795 14.978 42.569 15.018 ;
      RECT MASK 1 43.455 14.978 44.229 15.018 ;
      RECT MASK 1 50.095 14.978 50.869 15.018 ;
      RECT MASK 1 51.257 14.978 52.529 15.018 ;
      RECT MASK 1 53.415 14.978 54.189 15.018 ;
      RECT MASK 1 55.075 14.978 55.849 15.018 ;
      RECT MASK 1 56.901 14.978 57.675 15.018 ;
      RECT MASK 1 63.541 14.978 64.315 15.018 ;
      RECT MASK 1 65.201 14.978 65.975 15.018 ;
      RECT MASK 1 66.861 14.978 67.635 15.018 ;
      RECT MASK 1 68.521 14.978 69.295 15.018 ;
      RECT MASK 1 70.181 14.978 73.113 15.018 ;
      RECT MASK 1 76.821 14.978 77.595 15.018 ;
      RECT MASK 1 78.481 14.978 79.255 15.018 ;
      RECT MASK 1 79.643 14.978 79.919 15.018 ;
      RECT MASK 1 81.111 14.978 81.3035 15.018 ;
      RECT MASK 1 83.461 14.978 84.235 15.018 ;
      RECT MASK 1 90.101 14.978 90.875 15.018 ;
      RECT MASK 1 91.761 14.978 92.535 15.018 ;
      RECT MASK 1 93.421 14.978 94.195 15.018 ;
      RECT MASK 1 95.081 14.978 95.855 15.018 ;
      RECT MASK 1 96.741 14.978 97.515 15.018 ;
      RECT MASK 1 103.381 14.978 104.155 15.018 ;
      RECT MASK 1 105.041 14.978 105.815 15.018 ;
      RECT MASK 1 106.701 14.978 107.475 15.018 ;
      RECT MASK 1 110.021 14.978 110.795 15.018 ;
      RECT MASK 1 116.256 14.98 128.056 15.02 ;
      RECT MASK 1 4.251 15.198 111.819 15.398 ;
      RECT MASK 1 116.256 15.22 128.056 15.26 ;
      RECT MASK 1 116.256 15.46 128.056 15.5 ;
      RECT MASK 1 116.256 15.7 128.056 15.74 ;
      RECT MASK 1 116.256 15.94 128.056 15.98 ;
      RECT MASK 1 4.251 16.042 111.819 16.242 ;
      RECT MASK 1 116.256 16.18 128.056 16.22 ;
      RECT MASK 1 116.256 16.42 128.056 16.46 ;
      RECT MASK 1 11.417 16.422 105.815 16.462 ;
      RECT MASK 1 107.697 16.606 111.127 16.646 ;
      RECT MASK 1 8.595 16.612 107.143 16.652 ;
      RECT MASK 1 116.256 16.66 128.056 16.7 ;
      RECT MASK 1 4.943 16.804 6.381 16.844 ;
      RECT MASK 1 6.935 16.804 108.803 16.844 ;
      RECT MASK 1 116.256 16.9 128.056 16.94 ;
      RECT MASK 1 5.441 16.996 5.983 17.036 ;
      RECT MASK 1 7.014 16.996 7.543 17.036 ;
      RECT MASK 1 8.176 16.996 9.203 17.036 ;
      RECT MASK 1 10.421 16.996 10.863 17.036 ;
      RECT MASK 1 12.081 16.996 12.58 17.036 ;
      RECT MASK 1 13.632 16.996 14.183 17.036 ;
      RECT MASK 1 14.794 16.996 15.843 17.036 ;
      RECT MASK 1 16.3505 16.996 17.503 17.036 ;
      RECT MASK 1 18.721 16.996 19.198 17.036 ;
      RECT MASK 1 20.25 16.996 20.823 17.036 ;
      RECT MASK 1 22.041 16.996 22.483 17.036 ;
      RECT MASK 1 23.701 16.996 24.143 17.036 ;
      RECT MASK 1 25.361 16.996 25.816 17.036 ;
      RECT MASK 1 26.868 16.996 27.463 17.036 ;
      RECT MASK 1 28.03 16.996 29.123 17.036 ;
      RECT MASK 1 29.677 16.996 30.783 17.036 ;
      RECT MASK 1 32.001 16.996 32.443 17.036 ;
      RECT MASK 1 33.486 16.996 34.103 17.036 ;
      RECT MASK 1 34.648 16.996 35.763 17.036 ;
      RECT MASK 1 36.981 16.996 37.423 17.036 ;
      RECT MASK 1 38.641 16.996 39.083 17.036 ;
      RECT MASK 1 40.104 16.996 40.743 17.036 ;
      RECT MASK 1 41.266 16.996 42.403 17.036 ;
      RECT MASK 1 42.957 16.996 44.063 17.036 ;
      RECT MASK 1 45.281 16.996 45.723 17.036 ;
      RECT MASK 1 46.722 16.996 47.383 17.036 ;
      RECT MASK 1 47.884 16.996 49.043 17.036 ;
      RECT MASK 1 50.261 16.996 50.703 17.036 ;
      RECT MASK 1 51.921 16.996 53.072 17.036 ;
      RECT MASK 1 53.34 16.996 54.023 17.036 ;
      RECT MASK 1 54.502 16.996 55.683 17.036 ;
      RECT MASK 1 56.403 16.996 57.509 17.036 ;
      RECT MASK 1 58.727 16.996 59.169 17.036 ;
      RECT MASK 1 59.958 16.996 60.829 17.036 ;
      RECT MASK 1 61.12 16.996 62.489 17.036 ;
      RECT MASK 1 63.707 16.996 64.149 17.036 ;
      RECT MASK 1 65.367 16.996 65.809 17.036 ;
      RECT MASK 1 66.576 16.996 67.469 17.036 ;
      RECT MASK 1 67.738 16.996 69.129 17.036 ;
      RECT MASK 1 69.6805 16.996 70.789 17.036 ;
      RECT MASK 1 72.007 16.996 72.449 17.036 ;
      RECT MASK 1 73.194 16.996 74.109 17.036 ;
      RECT MASK 1 74.356 16.996 75.769 17.036 ;
      RECT MASK 1 76.987 16.996 77.429 17.036 ;
      RECT MASK 1 78.647 16.996 79.089 17.036 ;
      RECT MASK 1 79.812 16.996 80.749 17.036 ;
      RECT MASK 1 81.297 16.996 82.409 17.036 ;
      RECT MASK 1 82.963 16.996 84.069 17.036 ;
      RECT MASK 1 85.268 16.996 85.729 17.036 ;
      RECT MASK 1 86.43 16.996 87.389 17.036 ;
      RECT MASK 1 87.592 16.996 89.049 17.036 ;
      RECT MASK 1 90.267 16.996 90.709 17.036 ;
      RECT MASK 1 91.886 16.996 92.369 17.036 ;
      RECT MASK 1 93.048 16.996 94.029 17.036 ;
      RECT MASK 1 94.21 16.996 95.689 17.036 ;
      RECT MASK 1 96.243 16.996 97.349 17.036 ;
      RECT MASK 1 98.504 16.996 99.009 17.036 ;
      RECT MASK 1 99.666 16.996 100.669 17.036 ;
      RECT MASK 1 100.828 16.996 102.329 17.036 ;
      RECT MASK 1 103.547 16.996 103.989 17.036 ;
      RECT MASK 1 105.122 16.996 105.649 17.036 ;
      RECT MASK 1 106.284 16.996 107.309 17.036 ;
      RECT MASK 1 107.446 16.996 108.969 17.036 ;
      RECT MASK 1 109.5195 16.996 110.629 17.036 ;
      RECT MASK 1 116.256 17.14 128.056 17.18 ;
      RECT MASK 1 9.338 17.374 10.697 17.414 ;
      RECT MASK 1 11.722 17.374 12.202 17.414 ;
      RECT MASK 1 15.956 17.374 16.507 17.414 ;
      RECT MASK 1 18.246 17.374 18.82 17.414 ;
      RECT MASK 1 21.412 17.374 22.317 17.414 ;
      RECT MASK 1 22.574 17.374 23.9735 17.414 ;
      RECT MASK 1 24.56 17.374 25.438 17.414 ;
      RECT MASK 1 29.192 17.374 29.787 17.414 ;
      RECT MASK 1 31.337 17.374 32.056 17.414 ;
      RECT MASK 1 35.81 17.374 37.257 17.414 ;
      RECT MASK 1 37.566 17.374 38.674 17.414 ;
      RECT MASK 1 42.428 17.374 43.067 17.414 ;
      RECT MASK 1 44.166 17.374 45.292 17.414 ;
      RECT MASK 1 49.046 17.374 50.537 17.414 ;
      RECT MASK 1 51.004 17.374 51.91 17.414 ;
      RECT MASK 1 55.664 17.374 56.513 17.414 ;
      RECT MASK 1 58.063 17.374 58.528 17.414 ;
      RECT MASK 1 62.282 17.374 63.983 17.414 ;
      RECT MASK 1 64.314 17.374 65.146 17.414 ;
      RECT MASK 1 68.9 17.374 69.793 17.414 ;
      RECT MASK 1 71.343 17.374 71.764 17.414 ;
      RECT MASK 1 75.518 17.374 77.263 17.414 ;
      RECT MASK 1 77.983 17.374 78.382 17.414 ;
      RECT MASK 1 80.596 17.374 81.413 17.414 ;
      RECT MASK 1 82.136 17.374 83.073 17.414 ;
      RECT MASK 1 84.052 17.374 85 17.414 ;
      RECT MASK 1 88.754 17.374 90.543 17.414 ;
      RECT MASK 1 90.892 17.374 91.618 17.414 ;
      RECT MASK 1 95.372 17.374 96.353 17.414 ;
      RECT MASK 1 97.588 17.374 98.236 17.414 ;
      RECT MASK 1 101.99 17.374 103.823 17.414 ;
      RECT MASK 1 104.104 17.374 104.854 17.414 ;
      RECT MASK 1 108.608 17.374 109.633 17.414 ;
      RECT MASK 1 116.256 17.38 128.056 17.42 ;
      RECT MASK 1 116.256 17.62 128.056 17.66 ;
      RECT MASK 1 116.256 17.86 128.056 17.9 ;
      RECT MASK 1 116.256 18.1 128.056 18.14 ;
      RECT MASK 1 116.256 18.34 128.056 18.38 ;
      RECT MASK 1 116.256 18.58 128.056 18.62 ;
      RECT MASK 1 116.256 18.82 128.056 18.86 ;
      RECT MASK 1 116.256 19.06 128.056 19.1 ;
      RECT MASK 1 116.256 19.3 128.056 19.34 ;
      RECT MASK 1 116.256 19.54 128.056 19.58 ;
      RECT MASK 1 5.031 19.542 109.945 19.722 ;
      RECT MASK 1 2.327 19.66 3.827 19.7 ;
      RECT MASK 1 116.256 19.78 128.056 19.82 ;
      RECT MASK 1 2.327 19.9 3.827 19.94 ;
      RECT MASK 1 116.256 20.02 128.056 20.06 ;
      RECT MASK 1 2.327 20.14 3.827 20.18 ;
      RECT MASK 1 116.256 20.26 128.056 20.3 ;
      RECT MASK 1 2.327 20.38 3.827 20.42 ;
      RECT MASK 1 56.4625 20.42 58.3775 20.48 ;
      RECT MASK 1 5.6945 20.44 6.023 20.54 ;
      RECT MASK 1 6.8565 20.44 7.185 20.54 ;
      RECT MASK 1 8.0185 20.44 8.347 20.54 ;
      RECT MASK 1 9.1805 20.44 9.509 20.54 ;
      RECT MASK 1 12.3125 20.44 12.641 20.54 ;
      RECT MASK 1 13.4745 20.44 13.803 20.54 ;
      RECT MASK 1 14.6365 20.44 14.965 20.54 ;
      RECT MASK 1 15.7985 20.44 16.127 20.54 ;
      RECT MASK 1 18.9305 20.44 19.259 20.54 ;
      RECT MASK 1 20.0925 20.44 20.421 20.54 ;
      RECT MASK 1 21.2545 20.44 21.583 20.54 ;
      RECT MASK 1 22.4165 20.44 22.745 20.54 ;
      RECT MASK 1 25.5485 20.44 25.877 20.54 ;
      RECT MASK 1 26.7105 20.44 27.039 20.54 ;
      RECT MASK 1 27.8725 20.44 28.201 20.54 ;
      RECT MASK 1 29.0345 20.44 29.363 20.54 ;
      RECT MASK 1 32.1665 20.44 32.495 20.54 ;
      RECT MASK 1 33.3285 20.44 33.657 20.54 ;
      RECT MASK 1 34.4905 20.44 34.819 20.54 ;
      RECT MASK 1 35.6525 20.44 35.981 20.54 ;
      RECT MASK 1 38.7845 20.44 39.113 20.54 ;
      RECT MASK 1 39.9465 20.44 40.275 20.54 ;
      RECT MASK 1 41.1085 20.44 41.437 20.54 ;
      RECT MASK 1 42.2705 20.44 42.599 20.54 ;
      RECT MASK 1 45.4025 20.44 45.731 20.54 ;
      RECT MASK 1 46.5645 20.44 46.893 20.54 ;
      RECT MASK 1 47.7265 20.44 48.055 20.54 ;
      RECT MASK 1 48.8885 20.44 49.217 20.54 ;
      RECT MASK 1 52.0205 20.44 52.349 20.54 ;
      RECT MASK 1 53.1825 20.44 53.511 20.54 ;
      RECT MASK 1 54.3445 20.44 54.673 20.54 ;
      RECT MASK 1 55.5065 20.44 55.835 20.54 ;
      RECT MASK 1 58.6385 20.44 58.967 20.54 ;
      RECT MASK 1 59.8005 20.44 60.129 20.54 ;
      RECT MASK 1 60.9625 20.44 61.291 20.54 ;
      RECT MASK 1 62.1245 20.44 62.453 20.54 ;
      RECT MASK 1 65.2565 20.44 65.585 20.54 ;
      RECT MASK 1 66.4185 20.44 66.747 20.54 ;
      RECT MASK 1 67.5805 20.44 67.909 20.54 ;
      RECT MASK 1 68.7425 20.44 69.071 20.54 ;
      RECT MASK 1 71.8745 20.44 72.203 20.54 ;
      RECT MASK 1 73.0365 20.44 73.365 20.54 ;
      RECT MASK 1 74.1985 20.44 74.527 20.54 ;
      RECT MASK 1 75.3605 20.44 75.689 20.54 ;
      RECT MASK 1 78.4925 20.44 78.821 20.54 ;
      RECT MASK 1 79.6545 20.44 79.983 20.54 ;
      RECT MASK 1 80.8165 20.44 81.145 20.54 ;
      RECT MASK 1 81.9785 20.44 82.307 20.54 ;
      RECT MASK 1 85.1105 20.44 85.439 20.54 ;
      RECT MASK 1 86.2725 20.44 86.601 20.54 ;
      RECT MASK 1 87.4345 20.44 87.763 20.54 ;
      RECT MASK 1 88.5965 20.44 88.925 20.54 ;
      RECT MASK 1 91.7285 20.44 92.057 20.54 ;
      RECT MASK 1 92.8905 20.44 93.219 20.54 ;
      RECT MASK 1 94.0525 20.44 94.381 20.54 ;
      RECT MASK 1 95.2145 20.44 95.543 20.54 ;
      RECT MASK 1 98.3465 20.44 98.675 20.54 ;
      RECT MASK 1 99.5085 20.44 99.837 20.54 ;
      RECT MASK 1 100.6705 20.44 100.999 20.54 ;
      RECT MASK 1 101.8325 20.44 102.161 20.54 ;
      RECT MASK 1 104.9645 20.44 105.293 20.54 ;
      RECT MASK 1 106.1265 20.44 106.455 20.54 ;
      RECT MASK 1 107.2885 20.44 107.617 20.54 ;
      RECT MASK 1 108.4505 20.44 108.779 20.54 ;
      RECT MASK 1 116.256 20.5 128.056 20.54 ;
      RECT MASK 1 2.327 20.62 3.827 20.66 ;
      RECT MASK 1 56.4625 20.66 58.3775 20.72 ;
      RECT MASK 1 116.256 20.74 128.056 20.78 ;
      RECT MASK 1 2.327 20.86 3.827 20.9 ;
      RECT MASK 1 5.031 20.9 109.945 21.1 ;
      RECT MASK 1 116.256 20.98 128.056 21.02 ;
      RECT MASK 1 2.327 21.1 3.827 21.14 ;
      RECT MASK 1 116.256 21.22 128.056 21.26 ;
      RECT MASK 1 2.327 21.34 3.827 21.38 ;
      RECT MASK 1 116.256 21.46 128.056 21.5 ;
      RECT MASK 1 2.327 21.58 3.827 21.62 ;
      RECT MASK 1 56.722 21.625 58.9155 21.685 ;
      RECT MASK 1 6.212 21.657 6.6935 21.717 ;
      RECT MASK 1 7.374 21.657 7.8555 21.717 ;
      RECT MASK 1 8.536 21.657 9.0175 21.717 ;
      RECT MASK 1 9.698 21.657 10.1795 21.717 ;
      RECT MASK 1 12.83 21.657 13.3115 21.717 ;
      RECT MASK 1 13.992 21.657 14.4735 21.717 ;
      RECT MASK 1 15.154 21.657 15.6355 21.717 ;
      RECT MASK 1 16.316 21.657 16.7975 21.717 ;
      RECT MASK 1 19.448 21.657 19.9295 21.717 ;
      RECT MASK 1 20.61 21.657 21.0915 21.717 ;
      RECT MASK 1 21.772 21.657 22.2535 21.717 ;
      RECT MASK 1 22.934 21.657 23.4155 21.717 ;
      RECT MASK 1 26.066 21.657 26.5475 21.717 ;
      RECT MASK 1 27.228 21.657 27.7095 21.717 ;
      RECT MASK 1 28.39 21.657 28.8715 21.717 ;
      RECT MASK 1 29.552 21.657 30.0335 21.717 ;
      RECT MASK 1 32.684 21.657 33.1655 21.717 ;
      RECT MASK 1 33.846 21.657 34.3275 21.717 ;
      RECT MASK 1 35.008 21.657 35.4895 21.717 ;
      RECT MASK 1 36.17 21.657 36.6515 21.717 ;
      RECT MASK 1 39.302 21.657 39.7835 21.717 ;
      RECT MASK 1 40.464 21.657 40.9455 21.717 ;
      RECT MASK 1 41.626 21.657 42.1075 21.717 ;
      RECT MASK 1 42.788 21.657 43.2695 21.717 ;
      RECT MASK 1 45.92 21.657 46.4015 21.717 ;
      RECT MASK 1 47.082 21.657 47.5635 21.717 ;
      RECT MASK 1 48.244 21.657 48.7255 21.717 ;
      RECT MASK 1 49.406 21.657 49.8875 21.717 ;
      RECT MASK 1 52.538 21.657 53.0195 21.717 ;
      RECT MASK 1 53.7 21.657 54.1815 21.717 ;
      RECT MASK 1 54.862 21.657 55.3435 21.717 ;
      RECT MASK 1 56.024 21.657 56.5055 21.717 ;
      RECT MASK 1 59.156 21.657 59.6375 21.717 ;
      RECT MASK 1 60.318 21.657 60.7995 21.717 ;
      RECT MASK 1 61.48 21.657 61.9615 21.717 ;
      RECT MASK 1 62.642 21.657 63.1235 21.717 ;
      RECT MASK 1 65.774 21.657 66.2555 21.717 ;
      RECT MASK 1 66.936 21.657 67.4175 21.717 ;
      RECT MASK 1 68.098 21.657 68.5795 21.717 ;
      RECT MASK 1 69.26 21.657 69.7415 21.717 ;
      RECT MASK 1 72.392 21.657 72.8735 21.717 ;
      RECT MASK 1 73.554 21.657 74.0355 21.717 ;
      RECT MASK 1 74.716 21.657 75.1975 21.717 ;
      RECT MASK 1 75.878 21.657 76.3595 21.717 ;
      RECT MASK 1 79.01 21.657 79.4915 21.717 ;
      RECT MASK 1 80.172 21.657 80.6535 21.717 ;
      RECT MASK 1 81.334 21.657 81.8155 21.717 ;
      RECT MASK 1 82.496 21.657 82.9775 21.717 ;
      RECT MASK 1 85.628 21.657 86.1095 21.717 ;
      RECT MASK 1 86.79 21.657 87.2715 21.717 ;
      RECT MASK 1 87.952 21.657 88.4335 21.717 ;
      RECT MASK 1 89.114 21.657 89.5955 21.717 ;
      RECT MASK 1 92.246 21.657 92.7275 21.717 ;
      RECT MASK 1 93.408 21.657 93.8895 21.717 ;
      RECT MASK 1 94.57 21.657 95.0515 21.717 ;
      RECT MASK 1 95.732 21.657 96.2135 21.717 ;
      RECT MASK 1 98.864 21.657 99.3455 21.717 ;
      RECT MASK 1 100.026 21.657 100.5075 21.717 ;
      RECT MASK 1 101.188 21.657 101.6695 21.717 ;
      RECT MASK 1 102.35 21.657 102.8315 21.717 ;
      RECT MASK 1 105.482 21.657 105.9635 21.717 ;
      RECT MASK 1 106.644 21.657 107.1255 21.717 ;
      RECT MASK 1 107.806 21.657 108.2875 21.717 ;
      RECT MASK 1 108.968 21.657 109.4495 21.717 ;
      RECT MASK 1 116.256 21.7 128.056 21.74 ;
      RECT MASK 1 2.327 21.82 3.827 21.86 ;
      RECT MASK 1 56.722 21.865 58.9155 21.925 ;
      RECT MASK 1 116.256 21.94 128.056 21.98 ;
      RECT MASK 1 2.327 22.06 3.827 22.1 ;
      RECT MASK 1 5.645 22.17 109.165 22.23 ;
      RECT MASK 1 116.256 22.18 128.056 22.22 ;
      RECT MASK 1 2.327 22.3 3.827 22.34 ;
      RECT MASK 1 116.256 22.42 128.056 22.46 ;
      RECT MASK 1 10.177 22.51 12.147 22.61 ;
      RECT MASK 1 16.795 22.51 18.765 22.61 ;
      RECT MASK 1 23.413 22.51 25.383 22.61 ;
      RECT MASK 1 30.031 22.51 32.001 22.61 ;
      RECT MASK 1 36.649 22.51 38.619 22.61 ;
      RECT MASK 1 43.267 22.51 45.237 22.61 ;
      RECT MASK 1 49.885 22.51 51.855 22.61 ;
      RECT MASK 1 56.503 22.51 58.473 22.61 ;
      RECT MASK 1 63.121 22.51 65.091 22.61 ;
      RECT MASK 1 69.739 22.51 71.709 22.61 ;
      RECT MASK 1 76.357 22.51 78.327 22.61 ;
      RECT MASK 1 82.975 22.51 84.945 22.61 ;
      RECT MASK 1 89.593 22.51 91.563 22.61 ;
      RECT MASK 1 96.211 22.51 98.181 22.61 ;
      RECT MASK 1 102.829 22.51 104.799 22.61 ;
      RECT MASK 1 109.447 22.51 112.744 22.61 ;
      RECT MASK 1 2.327 22.54 3.827 22.58 ;
      RECT MASK 1 116.256 22.66 128.056 22.7 ;
      RECT MASK 1 2.327 22.78 3.827 22.82 ;
      RECT MASK 1 5.645 22.89 109.165 22.95 ;
      RECT MASK 1 116.256 22.9 128.056 22.94 ;
      RECT MASK 1 2.327 23.02 3.827 23.06 ;
      RECT MASK 1 116.256 23.14 128.056 23.18 ;
      RECT MASK 1 2.327 23.26 3.827 23.3 ;
      RECT MASK 1 116.256 23.38 128.056 23.42 ;
      RECT MASK 1 2.327 23.5 3.827 23.54 ;
      RECT MASK 1 2.327 23.74 3.827 23.78 ;
      RECT MASK 1 2.327 23.98 3.827 24.02 ;
      RECT MASK 1 2.327 24.22 3.827 24.26 ;
      RECT MASK 1 10.177 24.234 12.147 24.334 ;
      RECT MASK 1 16.795 24.234 18.765 24.334 ;
      RECT MASK 1 23.413 24.234 25.383 24.334 ;
      RECT MASK 1 30.031 24.234 32.001 24.334 ;
      RECT MASK 1 36.649 24.234 38.619 24.334 ;
      RECT MASK 1 43.267 24.234 45.237 24.334 ;
      RECT MASK 1 49.885 24.234 51.855 24.334 ;
      RECT MASK 1 56.503 24.234 58.473 24.334 ;
      RECT MASK 1 63.121 24.234 65.091 24.334 ;
      RECT MASK 1 69.739 24.234 71.709 24.334 ;
      RECT MASK 1 76.357 24.234 78.327 24.334 ;
      RECT MASK 1 82.975 24.234 84.945 24.334 ;
      RECT MASK 1 89.593 24.234 91.563 24.334 ;
      RECT MASK 1 96.211 24.234 98.181 24.334 ;
      RECT MASK 1 102.829 24.234 104.799 24.334 ;
      RECT MASK 1 109.447 24.234 111.839 24.334 ;
      RECT MASK 1 2.327 24.46 3.827 24.5 ;
      RECT MASK 1 5.645 24.569 109.165 24.629 ;
      RECT MASK 1 5.645 25.289 109.165 25.349 ;
      RECT MASK 1 0.567 26.265 114.04 26.385 ;
      RECT MASK 1 115.506 26.505 126.992 26.625 ;
      RECT MASK 1 126.561 26.87 127.29 26.93 ;
      RECT MASK 1 116.318 26.94 126.334 27.14 ;
      RECT MASK 1 116.074 27.536 126.301 27.596 ;
      RECT MASK 1 126.561 27.65 127.29 27.71 ;
      RECT MASK 1 113.368 27.98 126.9585 28.18 ;
      RECT MASK 1 4.681 28.28 10.961 28.38 ;
      RECT MASK 1 11.299 28.28 17.579 28.38 ;
      RECT MASK 1 17.917 28.28 24.197 28.38 ;
      RECT MASK 1 24.535 28.28 30.815 28.38 ;
      RECT MASK 1 31.153 28.28 37.433 28.38 ;
      RECT MASK 1 37.771 28.28 44.051 28.38 ;
      RECT MASK 1 44.389 28.28 50.669 28.38 ;
      RECT MASK 1 51.007 28.28 57.287 28.38 ;
      RECT MASK 1 57.625 28.28 63.905 28.38 ;
      RECT MASK 1 64.243 28.28 70.523 28.38 ;
      RECT MASK 1 70.861 28.28 77.141 28.38 ;
      RECT MASK 1 77.479 28.28 83.759 28.38 ;
      RECT MASK 1 84.097 28.28 90.377 28.38 ;
      RECT MASK 1 90.715 28.28 96.995 28.38 ;
      RECT MASK 1 97.333 28.28 103.613 28.38 ;
      RECT MASK 1 103.951 28.28 110.231 28.38 ;
      RECT MASK 1 126.561 28.43 127.491 28.49 ;
      RECT MASK 1 116.317 28.5 126.333 28.7 ;
      RECT MASK 1 4.672 28.655 10.96 28.755 ;
      RECT MASK 1 11.29 28.655 17.578 28.755 ;
      RECT MASK 1 17.908 28.655 24.196 28.755 ;
      RECT MASK 1 24.526 28.655 30.814 28.755 ;
      RECT MASK 1 31.144 28.655 37.432 28.755 ;
      RECT MASK 1 37.762 28.655 44.05 28.755 ;
      RECT MASK 1 44.38 28.655 50.668 28.755 ;
      RECT MASK 1 50.998 28.655 57.286 28.755 ;
      RECT MASK 1 57.616 28.655 63.904 28.755 ;
      RECT MASK 1 64.234 28.655 70.522 28.755 ;
      RECT MASK 1 70.852 28.655 77.14 28.755 ;
      RECT MASK 1 77.47 28.655 83.758 28.755 ;
      RECT MASK 1 84.088 28.655 90.376 28.755 ;
      RECT MASK 1 90.706 28.655 96.994 28.755 ;
      RECT MASK 1 97.324 28.655 103.612 28.755 ;
      RECT MASK 1 103.942 28.655 110.23 28.755 ;
      RECT MASK 1 4.672 29.025 10.96 29.125 ;
      RECT MASK 1 11.29 29.025 17.578 29.125 ;
      RECT MASK 1 17.908 29.025 24.196 29.125 ;
      RECT MASK 1 24.526 29.025 30.814 29.125 ;
      RECT MASK 1 31.144 29.025 37.432 29.125 ;
      RECT MASK 1 37.762 29.025 44.05 29.125 ;
      RECT MASK 1 44.38 29.025 50.668 29.125 ;
      RECT MASK 1 50.998 29.025 57.286 29.125 ;
      RECT MASK 1 57.616 29.025 63.904 29.125 ;
      RECT MASK 1 64.234 29.025 70.522 29.125 ;
      RECT MASK 1 70.852 29.025 77.14 29.125 ;
      RECT MASK 1 77.47 29.025 83.758 29.125 ;
      RECT MASK 1 84.088 29.025 90.376 29.125 ;
      RECT MASK 1 90.706 29.025 96.994 29.125 ;
      RECT MASK 1 97.324 29.025 103.612 29.125 ;
      RECT MASK 1 103.942 29.025 110.23 29.125 ;
      RECT MASK 1 116.074 29.083 126.312 29.143 ;
      RECT MASK 1 126.561 29.2105 127.491 29.2705 ;
      RECT MASK 1 4.681 29.4 10.961 29.5 ;
      RECT MASK 1 11.299 29.4 17.579 29.5 ;
      RECT MASK 1 17.917 29.4 24.197 29.5 ;
      RECT MASK 1 24.535 29.4 30.815 29.5 ;
      RECT MASK 1 31.153 29.4 37.433 29.5 ;
      RECT MASK 1 37.771 29.4 44.051 29.5 ;
      RECT MASK 1 44.389 29.4 50.669 29.5 ;
      RECT MASK 1 51.007 29.4 57.287 29.5 ;
      RECT MASK 1 57.625 29.4 63.905 29.5 ;
      RECT MASK 1 64.243 29.4 70.523 29.5 ;
      RECT MASK 1 70.861 29.4 77.141 29.5 ;
      RECT MASK 1 77.479 29.4 83.759 29.5 ;
      RECT MASK 1 84.097 29.4 90.377 29.5 ;
      RECT MASK 1 90.715 29.4 96.995 29.5 ;
      RECT MASK 1 97.333 29.4 103.613 29.5 ;
      RECT MASK 1 103.951 29.4 110.231 29.5 ;
      RECT MASK 1 116.2105 29.54 126.3345 29.74 ;
      RECT MASK 1 4.672 29.775 10.96 29.875 ;
      RECT MASK 1 11.29 29.775 17.578 29.875 ;
      RECT MASK 1 17.908 29.775 24.196 29.875 ;
      RECT MASK 1 24.526 29.775 30.814 29.875 ;
      RECT MASK 1 31.144 29.775 37.432 29.875 ;
      RECT MASK 1 37.762 29.775 44.05 29.875 ;
      RECT MASK 1 44.38 29.775 50.668 29.875 ;
      RECT MASK 1 50.998 29.775 57.286 29.875 ;
      RECT MASK 1 57.616 29.775 63.904 29.875 ;
      RECT MASK 1 64.234 29.775 70.522 29.875 ;
      RECT MASK 1 70.852 29.775 77.14 29.875 ;
      RECT MASK 1 77.47 29.775 83.758 29.875 ;
      RECT MASK 1 84.088 29.775 90.376 29.875 ;
      RECT MASK 1 90.706 29.775 96.994 29.875 ;
      RECT MASK 1 97.324 29.775 103.612 29.875 ;
      RECT MASK 1 103.942 29.775 110.23 29.875 ;
      RECT MASK 1 4.672 30.145 10.96 30.245 ;
      RECT MASK 1 11.29 30.145 17.578 30.245 ;
      RECT MASK 1 17.908 30.145 24.196 30.245 ;
      RECT MASK 1 24.526 30.145 30.814 30.245 ;
      RECT MASK 1 31.144 30.145 37.432 30.245 ;
      RECT MASK 1 37.762 30.145 44.05 30.245 ;
      RECT MASK 1 44.38 30.145 50.668 30.245 ;
      RECT MASK 1 50.998 30.145 57.286 30.245 ;
      RECT MASK 1 57.616 30.145 63.904 30.245 ;
      RECT MASK 1 64.234 30.145 70.522 30.245 ;
      RECT MASK 1 70.852 30.145 77.14 30.245 ;
      RECT MASK 1 77.47 30.145 83.758 30.245 ;
      RECT MASK 1 84.088 30.145 90.376 30.245 ;
      RECT MASK 1 90.706 30.145 96.994 30.245 ;
      RECT MASK 1 97.324 30.145 103.612 30.245 ;
      RECT MASK 1 103.942 30.145 110.23 30.245 ;
      RECT MASK 1 115.506 30.315 127.11 30.435 ;
      RECT MASK 1 4.681 30.52 10.961 30.62 ;
      RECT MASK 1 11.299 30.52 17.579 30.62 ;
      RECT MASK 1 17.917 30.52 24.197 30.62 ;
      RECT MASK 1 24.535 30.52 30.815 30.62 ;
      RECT MASK 1 31.153 30.52 37.433 30.62 ;
      RECT MASK 1 37.771 30.52 44.051 30.62 ;
      RECT MASK 1 44.389 30.52 50.669 30.62 ;
      RECT MASK 1 51.007 30.52 57.287 30.62 ;
      RECT MASK 1 57.625 30.52 63.905 30.62 ;
      RECT MASK 1 64.243 30.52 70.523 30.62 ;
      RECT MASK 1 70.861 30.52 77.141 30.62 ;
      RECT MASK 1 77.479 30.52 83.759 30.62 ;
      RECT MASK 1 84.097 30.52 90.377 30.62 ;
      RECT MASK 1 90.715 30.52 96.995 30.62 ;
      RECT MASK 1 97.333 30.52 103.613 30.62 ;
      RECT MASK 1 103.951 30.52 110.231 30.62 ;
      RECT MASK 1 4.672 30.895 10.96 30.995 ;
      RECT MASK 1 11.29 30.895 17.578 30.995 ;
      RECT MASK 1 17.908 30.895 24.196 30.995 ;
      RECT MASK 1 24.526 30.895 30.814 30.995 ;
      RECT MASK 1 31.144 30.895 37.432 30.995 ;
      RECT MASK 1 37.762 30.895 44.05 30.995 ;
      RECT MASK 1 44.38 30.895 50.668 30.995 ;
      RECT MASK 1 50.998 30.895 57.286 30.995 ;
      RECT MASK 1 57.616 30.895 63.904 30.995 ;
      RECT MASK 1 64.234 30.895 70.522 30.995 ;
      RECT MASK 1 70.852 30.895 77.14 30.995 ;
      RECT MASK 1 77.47 30.895 83.758 30.995 ;
      RECT MASK 1 84.088 30.895 90.376 30.995 ;
      RECT MASK 1 90.706 30.895 96.994 30.995 ;
      RECT MASK 1 97.324 30.895 103.612 30.995 ;
      RECT MASK 1 103.942 30.895 110.23 30.995 ;
      RECT MASK 1 4.672 31.265 10.96 31.365 ;
      RECT MASK 1 11.29 31.265 17.578 31.365 ;
      RECT MASK 1 17.908 31.265 24.196 31.365 ;
      RECT MASK 1 24.526 31.265 30.814 31.365 ;
      RECT MASK 1 31.144 31.265 37.432 31.365 ;
      RECT MASK 1 37.762 31.265 44.05 31.365 ;
      RECT MASK 1 44.38 31.265 50.668 31.365 ;
      RECT MASK 1 50.998 31.265 57.286 31.365 ;
      RECT MASK 1 57.616 31.265 63.904 31.365 ;
      RECT MASK 1 64.234 31.265 70.522 31.365 ;
      RECT MASK 1 70.852 31.265 77.14 31.365 ;
      RECT MASK 1 77.47 31.265 83.758 31.365 ;
      RECT MASK 1 84.088 31.265 90.376 31.365 ;
      RECT MASK 1 90.706 31.265 96.994 31.365 ;
      RECT MASK 1 97.324 31.265 103.612 31.365 ;
      RECT MASK 1 103.942 31.265 110.23 31.365 ;
      RECT MASK 1 4.681 31.64 10.961 31.74 ;
      RECT MASK 1 11.299 31.64 17.579 31.74 ;
      RECT MASK 1 17.917 31.64 24.197 31.74 ;
      RECT MASK 1 24.535 31.64 30.815 31.74 ;
      RECT MASK 1 31.153 31.64 37.433 31.74 ;
      RECT MASK 1 37.771 31.64 44.051 31.74 ;
      RECT MASK 1 44.389 31.64 50.669 31.74 ;
      RECT MASK 1 51.007 31.64 57.287 31.74 ;
      RECT MASK 1 57.625 31.64 63.905 31.74 ;
      RECT MASK 1 64.243 31.64 70.523 31.74 ;
      RECT MASK 1 70.861 31.64 77.141 31.74 ;
      RECT MASK 1 77.479 31.64 83.759 31.74 ;
      RECT MASK 1 84.097 31.64 90.377 31.74 ;
      RECT MASK 1 90.715 31.64 96.995 31.74 ;
      RECT MASK 1 97.333 31.64 103.613 31.74 ;
      RECT MASK 1 103.951 31.64 110.231 31.74 ;
      RECT MASK 1 4.672 32.015 10.96 32.115 ;
      RECT MASK 1 11.29 32.015 17.578 32.115 ;
      RECT MASK 1 17.908 32.015 24.196 32.115 ;
      RECT MASK 1 24.526 32.015 30.814 32.115 ;
      RECT MASK 1 31.144 32.015 37.432 32.115 ;
      RECT MASK 1 37.762 32.015 44.05 32.115 ;
      RECT MASK 1 44.38 32.015 50.668 32.115 ;
      RECT MASK 1 50.998 32.015 57.286 32.115 ;
      RECT MASK 1 57.616 32.015 63.904 32.115 ;
      RECT MASK 1 64.234 32.015 70.522 32.115 ;
      RECT MASK 1 70.852 32.015 77.14 32.115 ;
      RECT MASK 1 77.47 32.015 83.758 32.115 ;
      RECT MASK 1 84.088 32.015 90.376 32.115 ;
      RECT MASK 1 90.706 32.015 96.994 32.115 ;
      RECT MASK 1 97.324 32.015 103.612 32.115 ;
      RECT MASK 1 103.942 32.015 110.23 32.115 ;
      RECT MASK 1 4.672 32.385 10.96 32.485 ;
      RECT MASK 1 11.29 32.385 17.578 32.485 ;
      RECT MASK 1 17.908 32.385 24.196 32.485 ;
      RECT MASK 1 24.526 32.385 30.814 32.485 ;
      RECT MASK 1 31.144 32.385 37.432 32.485 ;
      RECT MASK 1 37.762 32.385 44.05 32.485 ;
      RECT MASK 1 44.38 32.385 50.668 32.485 ;
      RECT MASK 1 50.998 32.385 57.286 32.485 ;
      RECT MASK 1 57.616 32.385 63.904 32.485 ;
      RECT MASK 1 64.234 32.385 70.522 32.485 ;
      RECT MASK 1 70.852 32.385 77.14 32.485 ;
      RECT MASK 1 77.47 32.385 83.758 32.485 ;
      RECT MASK 1 84.088 32.385 90.376 32.485 ;
      RECT MASK 1 90.706 32.385 96.994 32.485 ;
      RECT MASK 1 97.324 32.385 103.612 32.485 ;
      RECT MASK 1 103.942 32.385 110.23 32.485 ;
      RECT MASK 1 111.044 32.615 129.1315 32.675 ;
      RECT MASK 1 4.681 32.76 10.961 32.86 ;
      RECT MASK 1 11.299 32.76 17.579 32.86 ;
      RECT MASK 1 17.917 32.76 24.197 32.86 ;
      RECT MASK 1 24.535 32.76 30.815 32.86 ;
      RECT MASK 1 31.153 32.76 37.433 32.86 ;
      RECT MASK 1 37.771 32.76 44.051 32.86 ;
      RECT MASK 1 44.389 32.76 50.669 32.86 ;
      RECT MASK 1 51.007 32.76 57.287 32.86 ;
      RECT MASK 1 57.625 32.76 63.905 32.86 ;
      RECT MASK 1 64.243 32.76 70.523 32.86 ;
      RECT MASK 1 70.861 32.76 77.141 32.86 ;
      RECT MASK 1 77.479 32.76 83.759 32.86 ;
      RECT MASK 1 84.097 32.76 90.377 32.86 ;
      RECT MASK 1 90.715 32.76 96.995 32.86 ;
      RECT MASK 1 97.333 32.76 103.613 32.86 ;
      RECT MASK 1 103.951 32.76 110.231 32.86 ;
      RECT MASK 1 117.268 33.375 129.1315 33.435 ;
      RECT MASK 1 111.044 33.9725 127.58 34.0725 ;
      RECT MASK 1 111.044 34.2925 129.1315 34.5425 ;
      RECT MASK 1 4.681 34.37 10.961 34.47 ;
      RECT MASK 1 11.299 34.37 17.579 34.47 ;
      RECT MASK 1 17.917 34.37 24.197 34.47 ;
      RECT MASK 1 24.535 34.37 30.815 34.47 ;
      RECT MASK 1 31.153 34.37 37.433 34.47 ;
      RECT MASK 1 37.771 34.37 44.051 34.47 ;
      RECT MASK 1 44.389 34.37 50.669 34.47 ;
      RECT MASK 1 51.007 34.37 57.287 34.47 ;
      RECT MASK 1 57.625 34.37 63.905 34.47 ;
      RECT MASK 1 64.243 34.37 70.523 34.47 ;
      RECT MASK 1 70.861 34.37 77.141 34.47 ;
      RECT MASK 1 77.479 34.37 83.759 34.47 ;
      RECT MASK 1 84.097 34.37 90.377 34.47 ;
      RECT MASK 1 90.715 34.37 96.995 34.47 ;
      RECT MASK 1 97.333 34.37 103.613 34.47 ;
      RECT MASK 1 103.951 34.37 110.231 34.47 ;
      RECT MASK 1 4.672 34.745 10.96 34.845 ;
      RECT MASK 1 11.29 34.745 17.578 34.845 ;
      RECT MASK 1 17.908 34.745 24.196 34.845 ;
      RECT MASK 1 24.526 34.745 30.814 34.845 ;
      RECT MASK 1 31.144 34.745 37.432 34.845 ;
      RECT MASK 1 37.762 34.745 44.05 34.845 ;
      RECT MASK 1 44.38 34.745 50.668 34.845 ;
      RECT MASK 1 50.998 34.745 57.286 34.845 ;
      RECT MASK 1 57.616 34.745 63.904 34.845 ;
      RECT MASK 1 64.234 34.745 70.522 34.845 ;
      RECT MASK 1 70.852 34.745 77.14 34.845 ;
      RECT MASK 1 77.47 34.745 83.758 34.845 ;
      RECT MASK 1 84.088 34.745 90.376 34.845 ;
      RECT MASK 1 90.706 34.745 96.994 34.845 ;
      RECT MASK 1 97.324 34.745 103.612 34.845 ;
      RECT MASK 1 103.942 34.745 110.23 34.845 ;
      RECT MASK 1 111.044 34.8075 129.1315 34.9075 ;
      RECT MASK 1 4.672 35.115 10.96 35.215 ;
      RECT MASK 1 11.29 35.115 17.578 35.215 ;
      RECT MASK 1 17.908 35.115 24.196 35.215 ;
      RECT MASK 1 24.526 35.115 30.814 35.215 ;
      RECT MASK 1 31.144 35.115 37.432 35.215 ;
      RECT MASK 1 37.762 35.115 44.05 35.215 ;
      RECT MASK 1 44.38 35.115 50.668 35.215 ;
      RECT MASK 1 50.998 35.115 57.286 35.215 ;
      RECT MASK 1 57.616 35.115 63.904 35.215 ;
      RECT MASK 1 64.234 35.115 70.522 35.215 ;
      RECT MASK 1 70.852 35.115 77.14 35.215 ;
      RECT MASK 1 77.47 35.115 83.758 35.215 ;
      RECT MASK 1 84.088 35.115 90.376 35.215 ;
      RECT MASK 1 90.706 35.115 96.994 35.215 ;
      RECT MASK 1 97.324 35.115 103.612 35.215 ;
      RECT MASK 1 103.942 35.115 110.23 35.215 ;
      RECT MASK 1 111.044 35.3225 127.58 35.4225 ;
      RECT MASK 1 4.681 35.49 10.961 35.59 ;
      RECT MASK 1 11.299 35.49 17.579 35.59 ;
      RECT MASK 1 17.917 35.49 24.197 35.59 ;
      RECT MASK 1 24.535 35.49 30.815 35.59 ;
      RECT MASK 1 31.153 35.49 37.433 35.59 ;
      RECT MASK 1 37.771 35.49 44.051 35.59 ;
      RECT MASK 1 44.389 35.49 50.669 35.59 ;
      RECT MASK 1 51.007 35.49 57.287 35.59 ;
      RECT MASK 1 57.625 35.49 63.905 35.59 ;
      RECT MASK 1 64.243 35.49 70.523 35.59 ;
      RECT MASK 1 70.861 35.49 77.141 35.59 ;
      RECT MASK 1 77.479 35.49 83.759 35.59 ;
      RECT MASK 1 84.097 35.49 90.377 35.59 ;
      RECT MASK 1 90.715 35.49 96.995 35.59 ;
      RECT MASK 1 97.333 35.49 103.613 35.59 ;
      RECT MASK 1 103.951 35.49 110.231 35.59 ;
      RECT MASK 1 111.044 35.6425 129.1315 35.8925 ;
      RECT MASK 1 4.672 35.865 10.96 35.965 ;
      RECT MASK 1 11.29 35.865 17.578 35.965 ;
      RECT MASK 1 17.908 35.865 24.196 35.965 ;
      RECT MASK 1 24.526 35.865 30.814 35.965 ;
      RECT MASK 1 31.144 35.865 37.432 35.965 ;
      RECT MASK 1 37.762 35.865 44.05 35.965 ;
      RECT MASK 1 44.38 35.865 50.668 35.965 ;
      RECT MASK 1 50.998 35.865 57.286 35.965 ;
      RECT MASK 1 57.616 35.865 63.904 35.965 ;
      RECT MASK 1 64.234 35.865 70.522 35.965 ;
      RECT MASK 1 70.852 35.865 77.14 35.965 ;
      RECT MASK 1 77.47 35.865 83.758 35.965 ;
      RECT MASK 1 84.088 35.865 90.376 35.965 ;
      RECT MASK 1 90.706 35.865 96.994 35.965 ;
      RECT MASK 1 97.324 35.865 103.612 35.965 ;
      RECT MASK 1 103.942 35.865 110.23 35.965 ;
      RECT MASK 1 111.044 36.1575 129.1315 36.2575 ;
      RECT MASK 1 4.672 36.235 10.96 36.335 ;
      RECT MASK 1 11.29 36.235 17.578 36.335 ;
      RECT MASK 1 17.908 36.235 24.196 36.335 ;
      RECT MASK 1 24.526 36.235 30.814 36.335 ;
      RECT MASK 1 31.144 36.235 37.432 36.335 ;
      RECT MASK 1 37.762 36.235 44.05 36.335 ;
      RECT MASK 1 44.38 36.235 50.668 36.335 ;
      RECT MASK 1 50.998 36.235 57.286 36.335 ;
      RECT MASK 1 57.616 36.235 63.904 36.335 ;
      RECT MASK 1 64.234 36.235 70.522 36.335 ;
      RECT MASK 1 70.852 36.235 77.14 36.335 ;
      RECT MASK 1 77.47 36.235 83.758 36.335 ;
      RECT MASK 1 84.088 36.235 90.376 36.335 ;
      RECT MASK 1 90.706 36.235 96.994 36.335 ;
      RECT MASK 1 97.324 36.235 103.612 36.335 ;
      RECT MASK 1 103.942 36.235 110.23 36.335 ;
      RECT MASK 1 4.681 36.61 10.961 36.71 ;
      RECT MASK 1 11.299 36.61 17.579 36.71 ;
      RECT MASK 1 17.917 36.61 24.197 36.71 ;
      RECT MASK 1 24.535 36.61 30.815 36.71 ;
      RECT MASK 1 31.153 36.61 37.433 36.71 ;
      RECT MASK 1 37.771 36.61 44.051 36.71 ;
      RECT MASK 1 44.389 36.61 50.669 36.71 ;
      RECT MASK 1 51.007 36.61 57.287 36.71 ;
      RECT MASK 1 57.625 36.61 63.905 36.71 ;
      RECT MASK 1 64.243 36.61 70.523 36.71 ;
      RECT MASK 1 70.861 36.61 77.141 36.71 ;
      RECT MASK 1 77.479 36.61 83.759 36.71 ;
      RECT MASK 1 84.097 36.61 90.377 36.71 ;
      RECT MASK 1 90.715 36.61 96.995 36.71 ;
      RECT MASK 1 97.333 36.61 103.613 36.71 ;
      RECT MASK 1 103.951 36.61 110.231 36.71 ;
      RECT MASK 1 111.044 36.7075 127.58 36.8075 ;
      RECT MASK 1 4.672 36.985 10.96 37.085 ;
      RECT MASK 1 11.29 36.985 17.578 37.085 ;
      RECT MASK 1 17.908 36.985 24.196 37.085 ;
      RECT MASK 1 24.526 36.985 30.814 37.085 ;
      RECT MASK 1 31.144 36.985 37.432 37.085 ;
      RECT MASK 1 37.762 36.985 44.05 37.085 ;
      RECT MASK 1 44.38 36.985 50.668 37.085 ;
      RECT MASK 1 50.998 36.985 57.286 37.085 ;
      RECT MASK 1 57.616 36.985 63.904 37.085 ;
      RECT MASK 1 64.234 36.985 70.522 37.085 ;
      RECT MASK 1 70.852 36.985 77.14 37.085 ;
      RECT MASK 1 77.47 36.985 83.758 37.085 ;
      RECT MASK 1 84.088 36.985 90.376 37.085 ;
      RECT MASK 1 90.706 36.985 96.994 37.085 ;
      RECT MASK 1 97.324 36.985 103.612 37.085 ;
      RECT MASK 1 103.942 36.985 110.23 37.085 ;
      RECT MASK 1 111.044 37.0275 129.1315 37.2775 ;
      RECT MASK 1 4.672 37.355 10.96 37.455 ;
      RECT MASK 1 11.29 37.355 17.578 37.455 ;
      RECT MASK 1 17.908 37.355 24.196 37.455 ;
      RECT MASK 1 24.526 37.355 30.814 37.455 ;
      RECT MASK 1 31.144 37.355 37.432 37.455 ;
      RECT MASK 1 37.762 37.355 44.05 37.455 ;
      RECT MASK 1 44.38 37.355 50.668 37.455 ;
      RECT MASK 1 50.998 37.355 57.286 37.455 ;
      RECT MASK 1 57.616 37.355 63.904 37.455 ;
      RECT MASK 1 64.234 37.355 70.522 37.455 ;
      RECT MASK 1 70.852 37.355 77.14 37.455 ;
      RECT MASK 1 77.47 37.355 83.758 37.455 ;
      RECT MASK 1 84.088 37.355 90.376 37.455 ;
      RECT MASK 1 90.706 37.355 96.994 37.455 ;
      RECT MASK 1 97.324 37.355 103.612 37.455 ;
      RECT MASK 1 103.942 37.355 110.23 37.455 ;
      RECT MASK 1 111.044 37.5075 129.1315 37.6075 ;
      RECT MASK 1 4.681 37.73 10.961 37.83 ;
      RECT MASK 1 11.299 37.73 17.579 37.83 ;
      RECT MASK 1 17.917 37.73 24.197 37.83 ;
      RECT MASK 1 24.535 37.73 30.815 37.83 ;
      RECT MASK 1 31.153 37.73 37.433 37.83 ;
      RECT MASK 1 37.771 37.73 44.051 37.83 ;
      RECT MASK 1 44.389 37.73 50.669 37.83 ;
      RECT MASK 1 51.007 37.73 57.287 37.83 ;
      RECT MASK 1 57.625 37.73 63.905 37.83 ;
      RECT MASK 1 64.243 37.73 70.523 37.83 ;
      RECT MASK 1 70.861 37.73 77.141 37.83 ;
      RECT MASK 1 77.479 37.73 83.759 37.83 ;
      RECT MASK 1 84.097 37.73 90.377 37.83 ;
      RECT MASK 1 90.715 37.73 96.995 37.83 ;
      RECT MASK 1 97.333 37.73 103.613 37.83 ;
      RECT MASK 1 103.951 37.73 110.231 37.83 ;
      RECT MASK 1 111.044 38.0225 127.58 38.1225 ;
      RECT MASK 1 4.672 38.105 10.96 38.205 ;
      RECT MASK 1 11.29 38.105 17.578 38.205 ;
      RECT MASK 1 17.908 38.105 24.196 38.205 ;
      RECT MASK 1 24.526 38.105 30.814 38.205 ;
      RECT MASK 1 31.144 38.105 37.432 38.205 ;
      RECT MASK 1 37.762 38.105 44.05 38.205 ;
      RECT MASK 1 44.38 38.105 50.668 38.205 ;
      RECT MASK 1 50.998 38.105 57.286 38.205 ;
      RECT MASK 1 57.616 38.105 63.904 38.205 ;
      RECT MASK 1 64.234 38.105 70.522 38.205 ;
      RECT MASK 1 70.852 38.105 77.14 38.205 ;
      RECT MASK 1 77.47 38.105 83.758 38.205 ;
      RECT MASK 1 84.088 38.105 90.376 38.205 ;
      RECT MASK 1 90.706 38.105 96.994 38.205 ;
      RECT MASK 1 97.324 38.105 103.612 38.205 ;
      RECT MASK 1 103.942 38.105 110.23 38.205 ;
      RECT MASK 1 111.044 38.3425 129.1315 38.5925 ;
      RECT MASK 1 4.672 38.475 10.96 38.575 ;
      RECT MASK 1 11.29 38.475 17.578 38.575 ;
      RECT MASK 1 17.908 38.475 24.196 38.575 ;
      RECT MASK 1 24.526 38.475 30.814 38.575 ;
      RECT MASK 1 31.144 38.475 37.432 38.575 ;
      RECT MASK 1 37.762 38.475 44.05 38.575 ;
      RECT MASK 1 44.38 38.475 50.668 38.575 ;
      RECT MASK 1 50.998 38.475 57.286 38.575 ;
      RECT MASK 1 57.616 38.475 63.904 38.575 ;
      RECT MASK 1 64.234 38.475 70.522 38.575 ;
      RECT MASK 1 70.852 38.475 77.14 38.575 ;
      RECT MASK 1 77.47 38.475 83.758 38.575 ;
      RECT MASK 1 84.088 38.475 90.376 38.575 ;
      RECT MASK 1 90.706 38.475 96.994 38.575 ;
      RECT MASK 1 97.324 38.475 103.612 38.575 ;
      RECT MASK 1 103.942 38.475 110.23 38.575 ;
      RECT MASK 1 4.681 38.85 10.961 38.95 ;
      RECT MASK 1 11.299 38.85 17.579 38.95 ;
      RECT MASK 1 17.917 38.85 24.197 38.95 ;
      RECT MASK 1 24.535 38.85 30.815 38.95 ;
      RECT MASK 1 31.153 38.85 37.433 38.95 ;
      RECT MASK 1 37.771 38.85 44.051 38.95 ;
      RECT MASK 1 44.389 38.85 50.669 38.95 ;
      RECT MASK 1 51.007 38.85 57.287 38.95 ;
      RECT MASK 1 57.625 38.85 63.905 38.95 ;
      RECT MASK 1 64.243 38.85 70.523 38.95 ;
      RECT MASK 1 70.861 38.85 77.141 38.95 ;
      RECT MASK 1 77.479 38.85 83.759 38.95 ;
      RECT MASK 1 84.097 38.85 90.377 38.95 ;
      RECT MASK 1 90.715 38.85 96.995 38.95 ;
      RECT MASK 1 97.333 38.85 103.613 38.95 ;
      RECT MASK 1 103.951 38.85 110.231 38.95 ;
      RECT MASK 1 111.044 38.8575 129.1315 38.9575 ;
      RECT MASK 1 117.268 39.3725 127.58 39.4725 ;
      RECT MASK 1 117.268 39.6925 129.1315 39.9425 ;
      RECT MASK 1 111.044 40.2675 129.1315 40.3675 ;
      RECT MASK 1 4.681 40.49 10.961 40.59 ;
      RECT MASK 1 11.299 40.49 17.579 40.59 ;
      RECT MASK 1 17.917 40.49 24.197 40.59 ;
      RECT MASK 1 24.535 40.49 30.815 40.59 ;
      RECT MASK 1 31.153 40.49 37.433 40.59 ;
      RECT MASK 1 37.771 40.49 44.051 40.59 ;
      RECT MASK 1 44.389 40.49 50.669 40.59 ;
      RECT MASK 1 51.007 40.49 57.287 40.59 ;
      RECT MASK 1 57.625 40.49 63.905 40.59 ;
      RECT MASK 1 64.243 40.49 70.523 40.59 ;
      RECT MASK 1 70.861 40.49 77.141 40.59 ;
      RECT MASK 1 77.479 40.49 83.759 40.59 ;
      RECT MASK 1 84.097 40.49 90.377 40.59 ;
      RECT MASK 1 90.715 40.49 96.995 40.59 ;
      RECT MASK 1 97.333 40.49 103.613 40.59 ;
      RECT MASK 1 103.951 40.49 110.231 40.59 ;
      RECT MASK 1 111.044 40.7825 129.1315 40.8825 ;
      RECT MASK 1 4.672 40.865 10.96 40.965 ;
      RECT MASK 1 11.29 40.865 17.578 40.965 ;
      RECT MASK 1 17.908 40.865 24.196 40.965 ;
      RECT MASK 1 24.526 40.865 30.814 40.965 ;
      RECT MASK 1 31.144 40.865 37.432 40.965 ;
      RECT MASK 1 37.762 40.865 44.05 40.965 ;
      RECT MASK 1 44.38 40.865 50.668 40.965 ;
      RECT MASK 1 50.998 40.865 57.286 40.965 ;
      RECT MASK 1 57.616 40.865 63.904 40.965 ;
      RECT MASK 1 64.234 40.865 70.522 40.965 ;
      RECT MASK 1 70.852 40.865 77.14 40.965 ;
      RECT MASK 1 77.47 40.865 83.758 40.965 ;
      RECT MASK 1 84.088 40.865 90.376 40.965 ;
      RECT MASK 1 90.706 40.865 96.994 40.965 ;
      RECT MASK 1 97.324 40.865 103.612 40.965 ;
      RECT MASK 1 103.942 40.865 110.23 40.965 ;
      RECT MASK 1 111.044 41.1025 129.1315 41.3525 ;
      RECT MASK 1 4.672 41.235 10.96 41.335 ;
      RECT MASK 1 11.29 41.235 17.578 41.335 ;
      RECT MASK 1 17.908 41.235 24.196 41.335 ;
      RECT MASK 1 24.526 41.235 30.814 41.335 ;
      RECT MASK 1 31.144 41.235 37.432 41.335 ;
      RECT MASK 1 37.762 41.235 44.05 41.335 ;
      RECT MASK 1 44.38 41.235 50.668 41.335 ;
      RECT MASK 1 50.998 41.235 57.286 41.335 ;
      RECT MASK 1 57.616 41.235 63.904 41.335 ;
      RECT MASK 1 64.234 41.235 70.522 41.335 ;
      RECT MASK 1 70.852 41.235 77.14 41.335 ;
      RECT MASK 1 77.47 41.235 83.758 41.335 ;
      RECT MASK 1 84.088 41.235 90.376 41.335 ;
      RECT MASK 1 90.706 41.235 96.994 41.335 ;
      RECT MASK 1 97.324 41.235 103.612 41.335 ;
      RECT MASK 1 103.942 41.235 110.23 41.335 ;
      RECT MASK 1 4.681 41.61 10.961 41.71 ;
      RECT MASK 1 11.299 41.61 17.579 41.71 ;
      RECT MASK 1 17.917 41.61 24.197 41.71 ;
      RECT MASK 1 24.535 41.61 30.815 41.71 ;
      RECT MASK 1 31.153 41.61 37.433 41.71 ;
      RECT MASK 1 37.771 41.61 44.051 41.71 ;
      RECT MASK 1 44.389 41.61 50.669 41.71 ;
      RECT MASK 1 51.007 41.61 57.287 41.71 ;
      RECT MASK 1 57.625 41.61 63.905 41.71 ;
      RECT MASK 1 64.243 41.61 70.523 41.71 ;
      RECT MASK 1 70.861 41.61 77.141 41.71 ;
      RECT MASK 1 77.479 41.61 83.759 41.71 ;
      RECT MASK 1 84.097 41.61 90.377 41.71 ;
      RECT MASK 1 90.715 41.61 96.995 41.71 ;
      RECT MASK 1 97.333 41.61 103.613 41.71 ;
      RECT MASK 1 103.951 41.61 110.231 41.71 ;
      RECT MASK 1 111.044 41.6175 127.58 41.7175 ;
      RECT MASK 1 4.672 41.985 10.96 42.085 ;
      RECT MASK 1 11.29 41.985 17.578 42.085 ;
      RECT MASK 1 17.908 41.985 24.196 42.085 ;
      RECT MASK 1 24.526 41.985 30.814 42.085 ;
      RECT MASK 1 31.144 41.985 37.432 42.085 ;
      RECT MASK 1 37.762 41.985 44.05 42.085 ;
      RECT MASK 1 44.38 41.985 50.668 42.085 ;
      RECT MASK 1 50.998 41.985 57.286 42.085 ;
      RECT MASK 1 57.616 41.985 63.904 42.085 ;
      RECT MASK 1 64.234 41.985 70.522 42.085 ;
      RECT MASK 1 70.852 41.985 77.14 42.085 ;
      RECT MASK 1 77.47 41.985 83.758 42.085 ;
      RECT MASK 1 84.088 41.985 90.376 42.085 ;
      RECT MASK 1 90.706 41.985 96.994 42.085 ;
      RECT MASK 1 97.324 41.985 103.612 42.085 ;
      RECT MASK 1 103.942 41.985 110.23 42.085 ;
      RECT MASK 1 111.044 42.1325 129.1315 42.2325 ;
      RECT MASK 1 4.672 42.355 10.96 42.455 ;
      RECT MASK 1 11.29 42.355 17.578 42.455 ;
      RECT MASK 1 17.908 42.355 24.196 42.455 ;
      RECT MASK 1 24.526 42.355 30.814 42.455 ;
      RECT MASK 1 31.144 42.355 37.432 42.455 ;
      RECT MASK 1 37.762 42.355 44.05 42.455 ;
      RECT MASK 1 44.38 42.355 50.668 42.455 ;
      RECT MASK 1 50.998 42.355 57.286 42.455 ;
      RECT MASK 1 57.616 42.355 63.904 42.455 ;
      RECT MASK 1 64.234 42.355 70.522 42.455 ;
      RECT MASK 1 70.852 42.355 77.14 42.455 ;
      RECT MASK 1 77.47 42.355 83.758 42.455 ;
      RECT MASK 1 84.088 42.355 90.376 42.455 ;
      RECT MASK 1 90.706 42.355 96.994 42.455 ;
      RECT MASK 1 97.324 42.355 103.612 42.455 ;
      RECT MASK 1 103.942 42.355 110.23 42.455 ;
      RECT MASK 1 111.044 42.4525 129.1315 42.7025 ;
      RECT MASK 1 4.681 42.73 10.961 42.83 ;
      RECT MASK 1 11.299 42.73 17.579 42.83 ;
      RECT MASK 1 17.917 42.73 24.197 42.83 ;
      RECT MASK 1 24.535 42.73 30.815 42.83 ;
      RECT MASK 1 31.153 42.73 37.433 42.83 ;
      RECT MASK 1 37.771 42.73 44.051 42.83 ;
      RECT MASK 1 44.389 42.73 50.669 42.83 ;
      RECT MASK 1 51.007 42.73 57.287 42.83 ;
      RECT MASK 1 57.625 42.73 63.905 42.83 ;
      RECT MASK 1 64.243 42.73 70.523 42.83 ;
      RECT MASK 1 70.861 42.73 77.141 42.83 ;
      RECT MASK 1 77.479 42.73 83.759 42.83 ;
      RECT MASK 1 84.097 42.73 90.377 42.83 ;
      RECT MASK 1 90.715 42.73 96.995 42.83 ;
      RECT MASK 1 97.333 42.73 103.613 42.83 ;
      RECT MASK 1 103.951 42.73 110.231 42.83 ;
      RECT MASK 1 111.044 42.9675 129.1315 43.0675 ;
      RECT MASK 1 4.672 43.105 10.96 43.205 ;
      RECT MASK 1 11.29 43.105 17.578 43.205 ;
      RECT MASK 1 17.908 43.105 24.196 43.205 ;
      RECT MASK 1 24.526 43.105 30.814 43.205 ;
      RECT MASK 1 31.144 43.105 37.432 43.205 ;
      RECT MASK 1 37.762 43.105 44.05 43.205 ;
      RECT MASK 1 44.38 43.105 50.668 43.205 ;
      RECT MASK 1 50.998 43.105 57.286 43.205 ;
      RECT MASK 1 57.616 43.105 63.904 43.205 ;
      RECT MASK 1 64.234 43.105 70.522 43.205 ;
      RECT MASK 1 70.852 43.105 77.14 43.205 ;
      RECT MASK 1 77.47 43.105 83.758 43.205 ;
      RECT MASK 1 84.088 43.105 90.376 43.205 ;
      RECT MASK 1 90.706 43.105 96.994 43.205 ;
      RECT MASK 1 97.324 43.105 103.612 43.205 ;
      RECT MASK 1 103.942 43.105 110.23 43.205 ;
      RECT MASK 1 4.672 43.475 10.96 43.575 ;
      RECT MASK 1 11.29 43.475 17.578 43.575 ;
      RECT MASK 1 17.908 43.475 24.196 43.575 ;
      RECT MASK 1 24.526 43.475 30.814 43.575 ;
      RECT MASK 1 31.144 43.475 37.432 43.575 ;
      RECT MASK 1 37.762 43.475 44.05 43.575 ;
      RECT MASK 1 44.38 43.475 50.668 43.575 ;
      RECT MASK 1 50.998 43.475 57.286 43.575 ;
      RECT MASK 1 57.616 43.475 63.904 43.575 ;
      RECT MASK 1 64.234 43.475 70.522 43.575 ;
      RECT MASK 1 70.852 43.475 77.14 43.575 ;
      RECT MASK 1 77.47 43.475 83.758 43.575 ;
      RECT MASK 1 84.088 43.475 90.376 43.575 ;
      RECT MASK 1 90.706 43.475 96.994 43.575 ;
      RECT MASK 1 97.324 43.475 103.612 43.575 ;
      RECT MASK 1 103.942 43.475 110.23 43.575 ;
      RECT MASK 1 111.044 43.4825 129.1315 43.5825 ;
      RECT MASK 1 111.044 43.8025 129.1315 44.0525 ;
      RECT MASK 1 4.681 43.85 10.961 43.95 ;
      RECT MASK 1 11.299 43.85 17.579 43.95 ;
      RECT MASK 1 17.917 43.85 24.197 43.95 ;
      RECT MASK 1 24.535 43.85 30.815 43.95 ;
      RECT MASK 1 31.153 43.85 37.433 43.95 ;
      RECT MASK 1 37.771 43.85 44.051 43.95 ;
      RECT MASK 1 44.389 43.85 50.669 43.95 ;
      RECT MASK 1 51.007 43.85 57.287 43.95 ;
      RECT MASK 1 57.625 43.85 63.905 43.95 ;
      RECT MASK 1 64.243 43.85 70.523 43.95 ;
      RECT MASK 1 70.861 43.85 77.141 43.95 ;
      RECT MASK 1 77.479 43.85 83.759 43.95 ;
      RECT MASK 1 84.097 43.85 90.377 43.95 ;
      RECT MASK 1 90.715 43.85 96.995 43.95 ;
      RECT MASK 1 97.333 43.85 103.613 43.95 ;
      RECT MASK 1 103.951 43.85 110.231 43.95 ;
      RECT MASK 1 4.672 44.225 10.96 44.325 ;
      RECT MASK 1 11.29 44.225 17.578 44.325 ;
      RECT MASK 1 17.908 44.225 24.196 44.325 ;
      RECT MASK 1 24.526 44.225 30.814 44.325 ;
      RECT MASK 1 31.144 44.225 37.432 44.325 ;
      RECT MASK 1 37.762 44.225 44.05 44.325 ;
      RECT MASK 1 44.38 44.225 50.668 44.325 ;
      RECT MASK 1 50.998 44.225 57.286 44.325 ;
      RECT MASK 1 57.616 44.225 63.904 44.325 ;
      RECT MASK 1 64.234 44.225 70.522 44.325 ;
      RECT MASK 1 70.852 44.225 77.14 44.325 ;
      RECT MASK 1 77.47 44.225 83.758 44.325 ;
      RECT MASK 1 84.088 44.225 90.376 44.325 ;
      RECT MASK 1 90.706 44.225 96.994 44.325 ;
      RECT MASK 1 97.324 44.225 103.612 44.325 ;
      RECT MASK 1 103.942 44.225 110.23 44.325 ;
      RECT MASK 1 111.044 44.3175 129.1315 44.4175 ;
      RECT MASK 1 4.672 44.595 10.96 44.695 ;
      RECT MASK 1 11.29 44.595 17.578 44.695 ;
      RECT MASK 1 17.908 44.595 24.196 44.695 ;
      RECT MASK 1 24.526 44.595 30.814 44.695 ;
      RECT MASK 1 31.144 44.595 37.432 44.695 ;
      RECT MASK 1 37.762 44.595 44.05 44.695 ;
      RECT MASK 1 44.38 44.595 50.668 44.695 ;
      RECT MASK 1 50.998 44.595 57.286 44.695 ;
      RECT MASK 1 57.616 44.595 63.904 44.695 ;
      RECT MASK 1 64.234 44.595 70.522 44.695 ;
      RECT MASK 1 70.852 44.595 77.14 44.695 ;
      RECT MASK 1 77.47 44.595 83.758 44.695 ;
      RECT MASK 1 84.088 44.595 90.376 44.695 ;
      RECT MASK 1 90.706 44.595 96.994 44.695 ;
      RECT MASK 1 97.324 44.595 103.612 44.695 ;
      RECT MASK 1 103.942 44.595 110.23 44.695 ;
      RECT MASK 1 111.044 44.7875 129.1315 44.8875 ;
      RECT MASK 1 4.681 44.97 10.961 45.07 ;
      RECT MASK 1 11.299 44.97 17.579 45.07 ;
      RECT MASK 1 17.917 44.97 24.197 45.07 ;
      RECT MASK 1 24.535 44.97 30.815 45.07 ;
      RECT MASK 1 31.153 44.97 37.433 45.07 ;
      RECT MASK 1 37.771 44.97 44.051 45.07 ;
      RECT MASK 1 44.389 44.97 50.669 45.07 ;
      RECT MASK 1 51.007 44.97 57.287 45.07 ;
      RECT MASK 1 57.625 44.97 63.905 45.07 ;
      RECT MASK 1 64.243 44.97 70.523 45.07 ;
      RECT MASK 1 70.861 44.97 77.141 45.07 ;
      RECT MASK 1 77.479 44.97 83.759 45.07 ;
      RECT MASK 1 84.097 44.97 90.377 45.07 ;
      RECT MASK 1 90.715 44.97 96.995 45.07 ;
      RECT MASK 1 97.333 44.97 103.613 45.07 ;
      RECT MASK 1 103.951 44.97 110.231 45.07 ;
      RECT MASK 1 117.268 45.1525 129.1315 45.4025 ;
      RECT MASK 1 117.181 45.779 129.1315 45.819 ;
      RECT MASK 1 117.181 45.939 129.1315 45.979 ;
      RECT MASK 1 117.181 46.099 129.1315 46.139 ;
      RECT MASK 1 117.181 46.259 129.1315 46.299 ;
      RECT MASK 1 111.044 46.59 129.1315 46.65 ;
      RECT MASK 1 4.681 46.61 10.961 46.71 ;
      RECT MASK 1 11.299 46.61 17.579 46.71 ;
      RECT MASK 1 17.917 46.61 24.197 46.71 ;
      RECT MASK 1 24.535 46.61 30.815 46.71 ;
      RECT MASK 1 31.153 46.61 37.433 46.71 ;
      RECT MASK 1 37.771 46.61 44.051 46.71 ;
      RECT MASK 1 44.389 46.61 50.669 46.71 ;
      RECT MASK 1 51.007 46.61 57.287 46.71 ;
      RECT MASK 1 57.625 46.61 63.905 46.71 ;
      RECT MASK 1 64.243 46.61 70.523 46.71 ;
      RECT MASK 1 70.861 46.61 77.141 46.71 ;
      RECT MASK 1 77.479 46.61 83.759 46.71 ;
      RECT MASK 1 84.097 46.61 90.377 46.71 ;
      RECT MASK 1 90.715 46.61 96.995 46.71 ;
      RECT MASK 1 97.333 46.61 103.613 46.71 ;
      RECT MASK 1 103.951 46.61 110.231 46.71 ;
      RECT MASK 1 4.672 46.985 10.96 47.085 ;
      RECT MASK 1 11.29 46.985 17.578 47.085 ;
      RECT MASK 1 17.908 46.985 24.196 47.085 ;
      RECT MASK 1 24.526 46.985 30.814 47.085 ;
      RECT MASK 1 31.144 46.985 37.432 47.085 ;
      RECT MASK 1 37.762 46.985 44.05 47.085 ;
      RECT MASK 1 44.38 46.985 50.668 47.085 ;
      RECT MASK 1 50.998 46.985 57.286 47.085 ;
      RECT MASK 1 57.616 46.985 63.904 47.085 ;
      RECT MASK 1 64.234 46.985 70.522 47.085 ;
      RECT MASK 1 70.852 46.985 77.14 47.085 ;
      RECT MASK 1 77.47 46.985 83.758 47.085 ;
      RECT MASK 1 84.088 46.985 90.376 47.085 ;
      RECT MASK 1 90.706 46.985 96.994 47.085 ;
      RECT MASK 1 97.324 46.985 103.612 47.085 ;
      RECT MASK 1 103.942 46.985 110.23 47.085 ;
      RECT MASK 1 111.044 46.985 129.1315 47.085 ;
      RECT MASK 1 4.672 47.355 10.96 47.455 ;
      RECT MASK 1 11.29 47.355 17.578 47.455 ;
      RECT MASK 1 17.908 47.355 24.196 47.455 ;
      RECT MASK 1 24.526 47.355 30.814 47.455 ;
      RECT MASK 1 31.144 47.355 37.432 47.455 ;
      RECT MASK 1 37.762 47.355 44.05 47.455 ;
      RECT MASK 1 44.38 47.355 50.668 47.455 ;
      RECT MASK 1 50.998 47.355 57.286 47.455 ;
      RECT MASK 1 57.616 47.355 63.904 47.455 ;
      RECT MASK 1 64.234 47.355 70.522 47.455 ;
      RECT MASK 1 70.852 47.355 77.14 47.455 ;
      RECT MASK 1 77.47 47.355 83.758 47.455 ;
      RECT MASK 1 84.088 47.355 90.376 47.455 ;
      RECT MASK 1 90.706 47.355 96.994 47.455 ;
      RECT MASK 1 97.324 47.355 103.612 47.455 ;
      RECT MASK 1 103.942 47.355 110.23 47.455 ;
      RECT MASK 1 111.044 47.355 129.1315 47.455 ;
      RECT MASK 1 4.681 47.73 10.961 47.83 ;
      RECT MASK 1 11.299 47.73 17.579 47.83 ;
      RECT MASK 1 17.917 47.73 24.197 47.83 ;
      RECT MASK 1 24.535 47.73 30.815 47.83 ;
      RECT MASK 1 31.153 47.73 37.433 47.83 ;
      RECT MASK 1 37.771 47.73 44.051 47.83 ;
      RECT MASK 1 44.389 47.73 50.669 47.83 ;
      RECT MASK 1 51.007 47.73 57.287 47.83 ;
      RECT MASK 1 57.625 47.73 63.905 47.83 ;
      RECT MASK 1 64.243 47.73 70.523 47.83 ;
      RECT MASK 1 70.861 47.73 77.141 47.83 ;
      RECT MASK 1 77.479 47.73 83.759 47.83 ;
      RECT MASK 1 84.097 47.73 90.377 47.83 ;
      RECT MASK 1 90.715 47.73 96.995 47.83 ;
      RECT MASK 1 97.333 47.73 103.613 47.83 ;
      RECT MASK 1 103.951 47.73 110.231 47.83 ;
      RECT MASK 1 111.044 47.73 129.1315 47.83 ;
      RECT MASK 1 4.672 48.105 10.96 48.205 ;
      RECT MASK 1 11.29 48.105 17.578 48.205 ;
      RECT MASK 1 17.908 48.105 24.196 48.205 ;
      RECT MASK 1 24.526 48.105 30.814 48.205 ;
      RECT MASK 1 31.144 48.105 37.432 48.205 ;
      RECT MASK 1 37.762 48.105 44.05 48.205 ;
      RECT MASK 1 44.38 48.105 50.668 48.205 ;
      RECT MASK 1 50.998 48.105 57.286 48.205 ;
      RECT MASK 1 57.616 48.105 63.904 48.205 ;
      RECT MASK 1 64.234 48.105 70.522 48.205 ;
      RECT MASK 1 70.852 48.105 77.14 48.205 ;
      RECT MASK 1 77.47 48.105 83.758 48.205 ;
      RECT MASK 1 84.088 48.105 90.376 48.205 ;
      RECT MASK 1 90.706 48.105 96.994 48.205 ;
      RECT MASK 1 97.324 48.105 103.612 48.205 ;
      RECT MASK 1 103.942 48.105 110.23 48.205 ;
      RECT MASK 1 111.044 48.105 129.1315 48.205 ;
      RECT MASK 1 4.672 48.475 10.96 48.575 ;
      RECT MASK 1 11.29 48.475 17.578 48.575 ;
      RECT MASK 1 17.908 48.475 24.196 48.575 ;
      RECT MASK 1 24.526 48.475 30.814 48.575 ;
      RECT MASK 1 31.144 48.475 37.432 48.575 ;
      RECT MASK 1 37.762 48.475 44.05 48.575 ;
      RECT MASK 1 44.38 48.475 50.668 48.575 ;
      RECT MASK 1 50.998 48.475 57.286 48.575 ;
      RECT MASK 1 57.616 48.475 63.904 48.575 ;
      RECT MASK 1 64.234 48.475 70.522 48.575 ;
      RECT MASK 1 70.852 48.475 77.14 48.575 ;
      RECT MASK 1 77.47 48.475 83.758 48.575 ;
      RECT MASK 1 84.088 48.475 90.376 48.575 ;
      RECT MASK 1 90.706 48.475 96.994 48.575 ;
      RECT MASK 1 97.324 48.475 103.612 48.575 ;
      RECT MASK 1 103.942 48.475 110.23 48.575 ;
      RECT MASK 1 111.044 48.475 129.1315 48.575 ;
      RECT MASK 1 4.681 48.85 10.961 48.95 ;
      RECT MASK 1 11.299 48.85 17.579 48.95 ;
      RECT MASK 1 17.917 48.85 24.197 48.95 ;
      RECT MASK 1 24.535 48.85 30.815 48.95 ;
      RECT MASK 1 31.153 48.85 37.433 48.95 ;
      RECT MASK 1 37.771 48.85 44.051 48.95 ;
      RECT MASK 1 44.389 48.85 50.669 48.95 ;
      RECT MASK 1 51.007 48.85 57.287 48.95 ;
      RECT MASK 1 57.625 48.85 63.905 48.95 ;
      RECT MASK 1 64.243 48.85 70.523 48.95 ;
      RECT MASK 1 70.861 48.85 77.141 48.95 ;
      RECT MASK 1 77.479 48.85 83.759 48.95 ;
      RECT MASK 1 84.097 48.85 90.377 48.95 ;
      RECT MASK 1 90.715 48.85 96.995 48.95 ;
      RECT MASK 1 97.333 48.85 103.613 48.95 ;
      RECT MASK 1 103.951 48.85 110.231 48.95 ;
      RECT MASK 1 111.044 48.85 129.1315 48.95 ;
      RECT MASK 1 4.672 49.225 10.96 49.325 ;
      RECT MASK 1 11.29 49.225 17.578 49.325 ;
      RECT MASK 1 17.908 49.225 24.196 49.325 ;
      RECT MASK 1 24.526 49.225 30.814 49.325 ;
      RECT MASK 1 31.144 49.225 37.432 49.325 ;
      RECT MASK 1 37.762 49.225 44.05 49.325 ;
      RECT MASK 1 44.38 49.225 50.668 49.325 ;
      RECT MASK 1 50.998 49.225 57.286 49.325 ;
      RECT MASK 1 57.616 49.225 63.904 49.325 ;
      RECT MASK 1 64.234 49.225 70.522 49.325 ;
      RECT MASK 1 70.852 49.225 77.14 49.325 ;
      RECT MASK 1 77.47 49.225 83.758 49.325 ;
      RECT MASK 1 84.088 49.225 90.376 49.325 ;
      RECT MASK 1 90.706 49.225 96.994 49.325 ;
      RECT MASK 1 97.324 49.225 103.612 49.325 ;
      RECT MASK 1 103.942 49.225 110.23 49.325 ;
      RECT MASK 1 111.044 49.225 129.1315 49.325 ;
      RECT MASK 1 4.672 49.595 10.96 49.695 ;
      RECT MASK 1 11.29 49.595 17.578 49.695 ;
      RECT MASK 1 17.908 49.595 24.196 49.695 ;
      RECT MASK 1 24.526 49.595 30.814 49.695 ;
      RECT MASK 1 31.144 49.595 37.432 49.695 ;
      RECT MASK 1 37.762 49.595 44.05 49.695 ;
      RECT MASK 1 44.38 49.595 50.668 49.695 ;
      RECT MASK 1 50.998 49.595 57.286 49.695 ;
      RECT MASK 1 57.616 49.595 63.904 49.695 ;
      RECT MASK 1 64.234 49.595 70.522 49.695 ;
      RECT MASK 1 70.852 49.595 77.14 49.695 ;
      RECT MASK 1 77.47 49.595 83.758 49.695 ;
      RECT MASK 1 84.088 49.595 90.376 49.695 ;
      RECT MASK 1 90.706 49.595 96.994 49.695 ;
      RECT MASK 1 97.324 49.595 103.612 49.695 ;
      RECT MASK 1 103.942 49.595 110.23 49.695 ;
      RECT MASK 1 117.4265 49.595 127.58 49.695 ;
      RECT MASK 1 4.681 49.97 10.961 50.07 ;
      RECT MASK 1 11.299 49.97 17.579 50.07 ;
      RECT MASK 1 17.917 49.97 24.197 50.07 ;
      RECT MASK 1 24.535 49.97 30.815 50.07 ;
      RECT MASK 1 31.153 49.97 37.433 50.07 ;
      RECT MASK 1 37.771 49.97 44.051 50.07 ;
      RECT MASK 1 44.389 49.97 50.669 50.07 ;
      RECT MASK 1 51.007 49.97 57.287 50.07 ;
      RECT MASK 1 57.625 49.97 63.905 50.07 ;
      RECT MASK 1 64.243 49.97 70.523 50.07 ;
      RECT MASK 1 70.861 49.97 77.141 50.07 ;
      RECT MASK 1 77.479 49.97 83.759 50.07 ;
      RECT MASK 1 84.097 49.97 90.377 50.07 ;
      RECT MASK 1 90.715 49.97 96.995 50.07 ;
      RECT MASK 1 97.333 49.97 103.613 50.07 ;
      RECT MASK 1 103.951 49.97 110.231 50.07 ;
      RECT MASK 1 117.4265 49.97 127.58 50.07 ;
      RECT MASK 1 4.672 50.345 10.96 50.445 ;
      RECT MASK 1 11.29 50.345 17.578 50.445 ;
      RECT MASK 1 17.908 50.345 24.196 50.445 ;
      RECT MASK 1 24.526 50.345 30.814 50.445 ;
      RECT MASK 1 31.144 50.345 37.432 50.445 ;
      RECT MASK 1 37.762 50.345 44.05 50.445 ;
      RECT MASK 1 44.38 50.345 50.668 50.445 ;
      RECT MASK 1 50.998 50.345 57.286 50.445 ;
      RECT MASK 1 57.616 50.345 63.904 50.445 ;
      RECT MASK 1 64.234 50.345 70.522 50.445 ;
      RECT MASK 1 70.852 50.345 77.14 50.445 ;
      RECT MASK 1 77.47 50.345 83.758 50.445 ;
      RECT MASK 1 84.088 50.345 90.376 50.445 ;
      RECT MASK 1 90.706 50.345 96.994 50.445 ;
      RECT MASK 1 97.324 50.345 103.612 50.445 ;
      RECT MASK 1 103.942 50.345 110.23 50.445 ;
      RECT MASK 1 117.4265 50.345 127.58 50.445 ;
      RECT MASK 1 4.672 50.715 10.96 50.815 ;
      RECT MASK 1 11.29 50.715 17.578 50.815 ;
      RECT MASK 1 17.908 50.715 24.196 50.815 ;
      RECT MASK 1 24.526 50.715 30.814 50.815 ;
      RECT MASK 1 31.144 50.715 37.432 50.815 ;
      RECT MASK 1 37.762 50.715 44.05 50.815 ;
      RECT MASK 1 44.38 50.715 50.668 50.815 ;
      RECT MASK 1 50.998 50.715 57.286 50.815 ;
      RECT MASK 1 57.616 50.715 63.904 50.815 ;
      RECT MASK 1 64.234 50.715 70.522 50.815 ;
      RECT MASK 1 70.852 50.715 77.14 50.815 ;
      RECT MASK 1 77.47 50.715 83.758 50.815 ;
      RECT MASK 1 84.088 50.715 90.376 50.815 ;
      RECT MASK 1 90.706 50.715 96.994 50.815 ;
      RECT MASK 1 97.324 50.715 103.612 50.815 ;
      RECT MASK 1 103.942 50.715 110.23 50.815 ;
      RECT MASK 1 111.044 50.715 129.1315 50.815 ;
      RECT MASK 1 4.681 51.09 10.961 51.19 ;
      RECT MASK 1 11.299 51.09 17.579 51.19 ;
      RECT MASK 1 17.917 51.09 24.197 51.19 ;
      RECT MASK 1 24.535 51.09 30.815 51.19 ;
      RECT MASK 1 31.153 51.09 37.433 51.19 ;
      RECT MASK 1 37.771 51.09 44.051 51.19 ;
      RECT MASK 1 44.389 51.09 50.669 51.19 ;
      RECT MASK 1 51.007 51.09 57.287 51.19 ;
      RECT MASK 1 57.625 51.09 63.905 51.19 ;
      RECT MASK 1 64.243 51.09 70.523 51.19 ;
      RECT MASK 1 70.861 51.09 77.141 51.19 ;
      RECT MASK 1 77.479 51.09 83.759 51.19 ;
      RECT MASK 1 84.097 51.09 90.377 51.19 ;
      RECT MASK 1 90.715 51.09 96.995 51.19 ;
      RECT MASK 1 97.333 51.09 103.613 51.19 ;
      RECT MASK 1 103.951 51.09 110.231 51.19 ;
      RECT MASK 1 111.044 51.09 129.1315 51.19 ;
      RECT MASK 1 117.181 51.34 129.1315 51.38 ;
      RECT MASK 1 117.181 51.5 129.1315 51.54 ;
      RECT MASK 1 117.181 51.66 129.1315 51.7 ;
      RECT MASK 1 117.181 51.82 129.1315 51.86 ;
      RECT MASK 1 117.181 51.98 129.1315 52.02 ;
      RECT MASK 1 117.181 52.14 129.1315 52.18 ;
      RECT MASK 1 117.181 52.3 129.1315 52.34 ;
      RECT MASK 1 111.044 52.725 129.1315 52.825 ;
      RECT MASK 1 4.681 52.73 10.961 52.83 ;
      RECT MASK 1 11.299 52.73 17.579 52.83 ;
      RECT MASK 1 17.917 52.73 24.197 52.83 ;
      RECT MASK 1 24.535 52.73 30.815 52.83 ;
      RECT MASK 1 31.153 52.73 37.433 52.83 ;
      RECT MASK 1 37.771 52.73 44.051 52.83 ;
      RECT MASK 1 44.389 52.73 50.669 52.83 ;
      RECT MASK 1 51.007 52.73 57.287 52.83 ;
      RECT MASK 1 57.625 52.73 63.905 52.83 ;
      RECT MASK 1 64.243 52.73 70.523 52.83 ;
      RECT MASK 1 70.861 52.73 77.141 52.83 ;
      RECT MASK 1 77.479 52.73 83.759 52.83 ;
      RECT MASK 1 84.097 52.73 90.377 52.83 ;
      RECT MASK 1 90.715 52.73 96.995 52.83 ;
      RECT MASK 1 97.333 52.73 103.613 52.83 ;
      RECT MASK 1 103.951 52.73 110.231 52.83 ;
      RECT MASK 1 4.672 53.105 10.96 53.205 ;
      RECT MASK 1 11.29 53.105 17.578 53.205 ;
      RECT MASK 1 17.908 53.105 24.196 53.205 ;
      RECT MASK 1 24.526 53.105 30.814 53.205 ;
      RECT MASK 1 31.144 53.105 37.432 53.205 ;
      RECT MASK 1 37.762 53.105 44.05 53.205 ;
      RECT MASK 1 44.38 53.105 50.668 53.205 ;
      RECT MASK 1 50.998 53.105 57.286 53.205 ;
      RECT MASK 1 57.616 53.105 63.904 53.205 ;
      RECT MASK 1 64.234 53.105 70.522 53.205 ;
      RECT MASK 1 70.852 53.105 77.14 53.205 ;
      RECT MASK 1 77.47 53.105 83.758 53.205 ;
      RECT MASK 1 84.088 53.105 90.376 53.205 ;
      RECT MASK 1 90.706 53.105 96.994 53.205 ;
      RECT MASK 1 97.324 53.105 103.612 53.205 ;
      RECT MASK 1 103.942 53.105 110.23 53.205 ;
      RECT MASK 1 111.044 53.105 129.1315 53.205 ;
      RECT MASK 1 4.672 53.475 10.96 53.575 ;
      RECT MASK 1 11.29 53.475 17.578 53.575 ;
      RECT MASK 1 17.908 53.475 24.196 53.575 ;
      RECT MASK 1 24.526 53.475 30.814 53.575 ;
      RECT MASK 1 31.144 53.475 37.432 53.575 ;
      RECT MASK 1 37.762 53.475 44.05 53.575 ;
      RECT MASK 1 44.38 53.475 50.668 53.575 ;
      RECT MASK 1 50.998 53.475 57.286 53.575 ;
      RECT MASK 1 57.616 53.475 63.904 53.575 ;
      RECT MASK 1 64.234 53.475 70.522 53.575 ;
      RECT MASK 1 70.852 53.475 77.14 53.575 ;
      RECT MASK 1 77.47 53.475 83.758 53.575 ;
      RECT MASK 1 84.088 53.475 90.376 53.575 ;
      RECT MASK 1 90.706 53.475 96.994 53.575 ;
      RECT MASK 1 97.324 53.475 103.612 53.575 ;
      RECT MASK 1 103.942 53.475 110.23 53.575 ;
      RECT MASK 1 111.044 53.475 129.1315 53.575 ;
      RECT MASK 1 4.681 53.85 10.961 53.95 ;
      RECT MASK 1 11.299 53.85 17.579 53.95 ;
      RECT MASK 1 17.917 53.85 24.197 53.95 ;
      RECT MASK 1 24.535 53.85 30.815 53.95 ;
      RECT MASK 1 31.153 53.85 37.433 53.95 ;
      RECT MASK 1 37.771 53.85 44.051 53.95 ;
      RECT MASK 1 44.389 53.85 50.669 53.95 ;
      RECT MASK 1 51.007 53.85 57.287 53.95 ;
      RECT MASK 1 57.625 53.85 63.905 53.95 ;
      RECT MASK 1 64.243 53.85 70.523 53.95 ;
      RECT MASK 1 70.861 53.85 77.141 53.95 ;
      RECT MASK 1 77.479 53.85 83.759 53.95 ;
      RECT MASK 1 84.097 53.85 90.377 53.95 ;
      RECT MASK 1 90.715 53.85 96.995 53.95 ;
      RECT MASK 1 97.333 53.85 103.613 53.95 ;
      RECT MASK 1 103.951 53.85 110.231 53.95 ;
      RECT MASK 1 111.044 53.85 129.1315 53.95 ;
      RECT MASK 1 4.672 54.225 10.96 54.325 ;
      RECT MASK 1 11.29 54.225 17.578 54.325 ;
      RECT MASK 1 17.908 54.225 24.196 54.325 ;
      RECT MASK 1 24.526 54.225 30.814 54.325 ;
      RECT MASK 1 31.144 54.225 37.432 54.325 ;
      RECT MASK 1 37.762 54.225 44.05 54.325 ;
      RECT MASK 1 44.38 54.225 50.668 54.325 ;
      RECT MASK 1 50.998 54.225 57.286 54.325 ;
      RECT MASK 1 57.616 54.225 63.904 54.325 ;
      RECT MASK 1 64.234 54.225 70.522 54.325 ;
      RECT MASK 1 70.852 54.225 77.14 54.325 ;
      RECT MASK 1 77.47 54.225 83.758 54.325 ;
      RECT MASK 1 84.088 54.225 90.376 54.325 ;
      RECT MASK 1 90.706 54.225 96.994 54.325 ;
      RECT MASK 1 97.324 54.225 103.612 54.325 ;
      RECT MASK 1 103.942 54.225 110.23 54.325 ;
      RECT MASK 1 111.044 54.225 129.1315 54.325 ;
      RECT MASK 1 4.672 54.595 10.96 54.695 ;
      RECT MASK 1 11.29 54.595 17.578 54.695 ;
      RECT MASK 1 17.908 54.595 24.196 54.695 ;
      RECT MASK 1 24.526 54.595 30.814 54.695 ;
      RECT MASK 1 31.144 54.595 37.432 54.695 ;
      RECT MASK 1 37.762 54.595 44.05 54.695 ;
      RECT MASK 1 44.38 54.595 50.668 54.695 ;
      RECT MASK 1 50.998 54.595 57.286 54.695 ;
      RECT MASK 1 57.616 54.595 63.904 54.695 ;
      RECT MASK 1 64.234 54.595 70.522 54.695 ;
      RECT MASK 1 70.852 54.595 77.14 54.695 ;
      RECT MASK 1 77.47 54.595 83.758 54.695 ;
      RECT MASK 1 84.088 54.595 90.376 54.695 ;
      RECT MASK 1 90.706 54.595 96.994 54.695 ;
      RECT MASK 1 97.324 54.595 103.612 54.695 ;
      RECT MASK 1 103.942 54.595 110.23 54.695 ;
      RECT MASK 1 111.044 54.595 129.1315 54.695 ;
      RECT MASK 1 4.681 54.97 10.961 55.07 ;
      RECT MASK 1 11.299 54.97 17.579 55.07 ;
      RECT MASK 1 17.917 54.97 24.197 55.07 ;
      RECT MASK 1 24.535 54.97 30.815 55.07 ;
      RECT MASK 1 31.153 54.97 37.433 55.07 ;
      RECT MASK 1 37.771 54.97 44.051 55.07 ;
      RECT MASK 1 44.389 54.97 50.669 55.07 ;
      RECT MASK 1 51.007 54.97 57.287 55.07 ;
      RECT MASK 1 57.625 54.97 63.905 55.07 ;
      RECT MASK 1 64.243 54.97 70.523 55.07 ;
      RECT MASK 1 70.861 54.97 77.141 55.07 ;
      RECT MASK 1 77.479 54.97 83.759 55.07 ;
      RECT MASK 1 84.097 54.97 90.377 55.07 ;
      RECT MASK 1 90.715 54.97 96.995 55.07 ;
      RECT MASK 1 97.333 54.97 103.613 55.07 ;
      RECT MASK 1 103.951 54.97 110.231 55.07 ;
      RECT MASK 1 111.044 54.97 129.1315 55.07 ;
      RECT MASK 1 4.672 55.345 10.96 55.445 ;
      RECT MASK 1 11.29 55.345 17.578 55.445 ;
      RECT MASK 1 17.908 55.345 24.196 55.445 ;
      RECT MASK 1 24.526 55.345 30.814 55.445 ;
      RECT MASK 1 31.144 55.345 37.432 55.445 ;
      RECT MASK 1 37.762 55.345 44.05 55.445 ;
      RECT MASK 1 44.38 55.345 50.668 55.445 ;
      RECT MASK 1 50.998 55.345 57.286 55.445 ;
      RECT MASK 1 57.616 55.345 63.904 55.445 ;
      RECT MASK 1 64.234 55.345 70.522 55.445 ;
      RECT MASK 1 70.852 55.345 77.14 55.445 ;
      RECT MASK 1 77.47 55.345 83.758 55.445 ;
      RECT MASK 1 84.088 55.345 90.376 55.445 ;
      RECT MASK 1 90.706 55.345 96.994 55.445 ;
      RECT MASK 1 97.324 55.345 103.612 55.445 ;
      RECT MASK 1 103.942 55.345 110.23 55.445 ;
      RECT MASK 1 111.044 55.345 129.1315 55.445 ;
      RECT MASK 1 4.672 55.715 10.96 55.815 ;
      RECT MASK 1 11.29 55.715 17.578 55.815 ;
      RECT MASK 1 17.908 55.715 24.196 55.815 ;
      RECT MASK 1 24.526 55.715 30.814 55.815 ;
      RECT MASK 1 31.144 55.715 37.432 55.815 ;
      RECT MASK 1 37.762 55.715 44.05 55.815 ;
      RECT MASK 1 44.38 55.715 50.668 55.815 ;
      RECT MASK 1 50.998 55.715 57.286 55.815 ;
      RECT MASK 1 57.616 55.715 63.904 55.815 ;
      RECT MASK 1 64.234 55.715 70.522 55.815 ;
      RECT MASK 1 70.852 55.715 77.14 55.815 ;
      RECT MASK 1 77.47 55.715 83.758 55.815 ;
      RECT MASK 1 84.088 55.715 90.376 55.815 ;
      RECT MASK 1 90.706 55.715 96.994 55.815 ;
      RECT MASK 1 97.324 55.715 103.612 55.815 ;
      RECT MASK 1 103.942 55.715 110.23 55.815 ;
      RECT MASK 1 111.044 55.715 129.1315 55.815 ;
      RECT MASK 1 4.681 56.09 10.961 56.19 ;
      RECT MASK 1 11.299 56.09 17.579 56.19 ;
      RECT MASK 1 17.917 56.09 24.197 56.19 ;
      RECT MASK 1 24.535 56.09 30.815 56.19 ;
      RECT MASK 1 31.153 56.09 37.433 56.19 ;
      RECT MASK 1 37.771 56.09 44.051 56.19 ;
      RECT MASK 1 44.389 56.09 50.669 56.19 ;
      RECT MASK 1 51.007 56.09 57.287 56.19 ;
      RECT MASK 1 57.625 56.09 63.905 56.19 ;
      RECT MASK 1 64.243 56.09 70.523 56.19 ;
      RECT MASK 1 70.861 56.09 77.141 56.19 ;
      RECT MASK 1 77.479 56.09 83.759 56.19 ;
      RECT MASK 1 84.097 56.09 90.377 56.19 ;
      RECT MASK 1 90.715 56.09 96.995 56.19 ;
      RECT MASK 1 97.333 56.09 103.613 56.19 ;
      RECT MASK 1 103.951 56.09 110.231 56.19 ;
      RECT MASK 1 111.044 56.09 129.1315 56.19 ;
      RECT MASK 1 4.672 56.465 10.96 56.565 ;
      RECT MASK 1 11.29 56.465 17.578 56.565 ;
      RECT MASK 1 17.908 56.465 24.196 56.565 ;
      RECT MASK 1 24.526 56.465 30.814 56.565 ;
      RECT MASK 1 31.144 56.465 37.432 56.565 ;
      RECT MASK 1 37.762 56.465 44.05 56.565 ;
      RECT MASK 1 44.38 56.465 50.668 56.565 ;
      RECT MASK 1 50.998 56.465 57.286 56.565 ;
      RECT MASK 1 57.616 56.465 63.904 56.565 ;
      RECT MASK 1 64.234 56.465 70.522 56.565 ;
      RECT MASK 1 70.852 56.465 77.14 56.565 ;
      RECT MASK 1 77.47 56.465 83.758 56.565 ;
      RECT MASK 1 84.088 56.465 90.376 56.565 ;
      RECT MASK 1 90.706 56.465 96.994 56.565 ;
      RECT MASK 1 97.324 56.465 103.612 56.565 ;
      RECT MASK 1 103.942 56.465 110.23 56.565 ;
      RECT MASK 1 111.044 56.465 129.1315 56.565 ;
      RECT MASK 1 4.672 56.835 10.96 56.935 ;
      RECT MASK 1 11.29 56.835 17.578 56.935 ;
      RECT MASK 1 17.908 56.835 24.196 56.935 ;
      RECT MASK 1 24.526 56.835 30.814 56.935 ;
      RECT MASK 1 31.144 56.835 37.432 56.935 ;
      RECT MASK 1 37.762 56.835 44.05 56.935 ;
      RECT MASK 1 44.38 56.835 50.668 56.935 ;
      RECT MASK 1 50.998 56.835 57.286 56.935 ;
      RECT MASK 1 57.616 56.835 63.904 56.935 ;
      RECT MASK 1 64.234 56.835 70.522 56.935 ;
      RECT MASK 1 70.852 56.835 77.14 56.935 ;
      RECT MASK 1 77.47 56.835 83.758 56.935 ;
      RECT MASK 1 84.088 56.835 90.376 56.935 ;
      RECT MASK 1 90.706 56.835 96.994 56.935 ;
      RECT MASK 1 97.324 56.835 103.612 56.935 ;
      RECT MASK 1 103.942 56.835 110.23 56.935 ;
      RECT MASK 1 111.044 56.835 129.1315 56.935 ;
      RECT MASK 1 4.681 57.21 10.961 57.31 ;
      RECT MASK 1 11.299 57.21 17.579 57.31 ;
      RECT MASK 1 17.917 57.21 24.197 57.31 ;
      RECT MASK 1 24.535 57.21 30.815 57.31 ;
      RECT MASK 1 31.153 57.21 37.433 57.31 ;
      RECT MASK 1 37.771 57.21 44.051 57.31 ;
      RECT MASK 1 44.389 57.21 50.669 57.31 ;
      RECT MASK 1 51.007 57.21 57.287 57.31 ;
      RECT MASK 1 57.625 57.21 63.905 57.31 ;
      RECT MASK 1 64.243 57.21 70.523 57.31 ;
      RECT MASK 1 70.861 57.21 77.141 57.31 ;
      RECT MASK 1 77.479 57.21 83.759 57.31 ;
      RECT MASK 1 84.097 57.21 90.377 57.31 ;
      RECT MASK 1 90.715 57.21 96.995 57.31 ;
      RECT MASK 1 97.333 57.21 103.613 57.31 ;
      RECT MASK 1 103.951 57.21 110.231 57.31 ;
      RECT MASK 1 111.044 57.21 129.1315 57.31 ;
      RECT MASK 1 117.181 57.55 129.1315 57.59 ;
      RECT MASK 1 117.181 57.71 129.1315 57.75 ;
      RECT MASK 1 117.181 57.87 129.1315 57.91 ;
      RECT MASK 1 117.181 58.03 129.1315 58.07 ;
      RECT MASK 1 117.268 58.385 129.1315 58.485 ;
      RECT MASK 1 111.044 58.62 129.1315 58.68 ;
      RECT MASK 1 4.681 58.85 10.961 58.95 ;
      RECT MASK 1 11.299 58.85 17.579 58.95 ;
      RECT MASK 1 17.917 58.85 24.197 58.95 ;
      RECT MASK 1 24.535 58.85 30.815 58.95 ;
      RECT MASK 1 31.153 58.85 37.433 58.95 ;
      RECT MASK 1 37.771 58.85 44.051 58.95 ;
      RECT MASK 1 44.389 58.85 50.669 58.95 ;
      RECT MASK 1 51.007 58.85 57.287 58.95 ;
      RECT MASK 1 57.625 58.85 63.905 58.95 ;
      RECT MASK 1 64.243 58.85 70.523 58.95 ;
      RECT MASK 1 70.861 58.85 77.141 58.95 ;
      RECT MASK 1 77.479 58.85 83.759 58.95 ;
      RECT MASK 1 84.097 58.85 90.377 58.95 ;
      RECT MASK 1 90.715 58.85 96.995 58.95 ;
      RECT MASK 1 97.333 58.85 103.613 58.95 ;
      RECT MASK 1 103.951 58.85 110.231 58.95 ;
      RECT MASK 1 4.672 59.225 10.96 59.325 ;
      RECT MASK 1 11.29 59.225 17.578 59.325 ;
      RECT MASK 1 17.908 59.225 24.196 59.325 ;
      RECT MASK 1 24.526 59.225 30.814 59.325 ;
      RECT MASK 1 31.144 59.225 37.432 59.325 ;
      RECT MASK 1 37.762 59.225 44.05 59.325 ;
      RECT MASK 1 44.38 59.225 50.668 59.325 ;
      RECT MASK 1 50.998 59.225 57.286 59.325 ;
      RECT MASK 1 57.616 59.225 63.904 59.325 ;
      RECT MASK 1 64.234 59.225 70.522 59.325 ;
      RECT MASK 1 70.852 59.225 77.14 59.325 ;
      RECT MASK 1 77.47 59.225 83.758 59.325 ;
      RECT MASK 1 84.088 59.225 90.376 59.325 ;
      RECT MASK 1 90.706 59.225 96.994 59.325 ;
      RECT MASK 1 97.324 59.225 103.612 59.325 ;
      RECT MASK 1 103.942 59.225 110.23 59.325 ;
      RECT MASK 1 111.044 59.2625 127.58 59.3625 ;
      RECT MASK 1 117.268 59.5825 129.1315 59.8325 ;
      RECT MASK 1 4.672 59.595 10.96 59.695 ;
      RECT MASK 1 11.29 59.595 17.578 59.695 ;
      RECT MASK 1 17.908 59.595 24.196 59.695 ;
      RECT MASK 1 24.526 59.595 30.814 59.695 ;
      RECT MASK 1 31.144 59.595 37.432 59.695 ;
      RECT MASK 1 37.762 59.595 44.05 59.695 ;
      RECT MASK 1 44.38 59.595 50.668 59.695 ;
      RECT MASK 1 50.998 59.595 57.286 59.695 ;
      RECT MASK 1 57.616 59.595 63.904 59.695 ;
      RECT MASK 1 64.234 59.595 70.522 59.695 ;
      RECT MASK 1 70.852 59.595 77.14 59.695 ;
      RECT MASK 1 77.47 59.595 83.758 59.695 ;
      RECT MASK 1 84.088 59.595 90.376 59.695 ;
      RECT MASK 1 90.706 59.595 96.994 59.695 ;
      RECT MASK 1 97.324 59.595 103.612 59.695 ;
      RECT MASK 1 103.942 59.595 110.23 59.695 ;
      RECT MASK 1 4.681 59.97 10.961 60.07 ;
      RECT MASK 1 11.299 59.97 17.579 60.07 ;
      RECT MASK 1 17.917 59.97 24.197 60.07 ;
      RECT MASK 1 24.535 59.97 30.815 60.07 ;
      RECT MASK 1 31.153 59.97 37.433 60.07 ;
      RECT MASK 1 37.771 59.97 44.051 60.07 ;
      RECT MASK 1 44.389 59.97 50.669 60.07 ;
      RECT MASK 1 51.007 59.97 57.287 60.07 ;
      RECT MASK 1 57.625 59.97 63.905 60.07 ;
      RECT MASK 1 64.243 59.97 70.523 60.07 ;
      RECT MASK 1 70.861 59.97 77.141 60.07 ;
      RECT MASK 1 77.479 59.97 83.759 60.07 ;
      RECT MASK 1 84.097 59.97 90.377 60.07 ;
      RECT MASK 1 90.715 59.97 96.995 60.07 ;
      RECT MASK 1 97.333 59.97 103.613 60.07 ;
      RECT MASK 1 103.951 59.97 110.231 60.07 ;
      RECT MASK 1 111.044 60.0975 129.1315 60.1975 ;
      RECT MASK 1 4.672 60.345 10.96 60.445 ;
      RECT MASK 1 11.29 60.345 17.578 60.445 ;
      RECT MASK 1 17.908 60.345 24.196 60.445 ;
      RECT MASK 1 24.526 60.345 30.814 60.445 ;
      RECT MASK 1 31.144 60.345 37.432 60.445 ;
      RECT MASK 1 37.762 60.345 44.05 60.445 ;
      RECT MASK 1 44.38 60.345 50.668 60.445 ;
      RECT MASK 1 50.998 60.345 57.286 60.445 ;
      RECT MASK 1 57.616 60.345 63.904 60.445 ;
      RECT MASK 1 64.234 60.345 70.522 60.445 ;
      RECT MASK 1 70.852 60.345 77.14 60.445 ;
      RECT MASK 1 77.47 60.345 83.758 60.445 ;
      RECT MASK 1 84.088 60.345 90.376 60.445 ;
      RECT MASK 1 90.706 60.345 96.994 60.445 ;
      RECT MASK 1 97.324 60.345 103.612 60.445 ;
      RECT MASK 1 103.942 60.345 110.23 60.445 ;
      RECT MASK 1 111.044 60.6125 127.58 60.7125 ;
      RECT MASK 1 4.672 60.715 10.96 60.815 ;
      RECT MASK 1 11.29 60.715 17.578 60.815 ;
      RECT MASK 1 17.908 60.715 24.196 60.815 ;
      RECT MASK 1 24.526 60.715 30.814 60.815 ;
      RECT MASK 1 31.144 60.715 37.432 60.815 ;
      RECT MASK 1 37.762 60.715 44.05 60.815 ;
      RECT MASK 1 44.38 60.715 50.668 60.815 ;
      RECT MASK 1 50.998 60.715 57.286 60.815 ;
      RECT MASK 1 57.616 60.715 63.904 60.815 ;
      RECT MASK 1 64.234 60.715 70.522 60.815 ;
      RECT MASK 1 70.852 60.715 77.14 60.815 ;
      RECT MASK 1 77.47 60.715 83.758 60.815 ;
      RECT MASK 1 84.088 60.715 90.376 60.815 ;
      RECT MASK 1 90.706 60.715 96.994 60.815 ;
      RECT MASK 1 97.324 60.715 103.612 60.815 ;
      RECT MASK 1 103.942 60.715 110.23 60.815 ;
      RECT MASK 1 111.044 60.9325 129.1315 61.1825 ;
      RECT MASK 1 4.681 61.09 10.961 61.19 ;
      RECT MASK 1 11.299 61.09 17.579 61.19 ;
      RECT MASK 1 17.917 61.09 24.197 61.19 ;
      RECT MASK 1 24.535 61.09 30.815 61.19 ;
      RECT MASK 1 31.153 61.09 37.433 61.19 ;
      RECT MASK 1 37.771 61.09 44.051 61.19 ;
      RECT MASK 1 44.389 61.09 50.669 61.19 ;
      RECT MASK 1 51.007 61.09 57.287 61.19 ;
      RECT MASK 1 57.625 61.09 63.905 61.19 ;
      RECT MASK 1 64.243 61.09 70.523 61.19 ;
      RECT MASK 1 70.861 61.09 77.141 61.19 ;
      RECT MASK 1 77.479 61.09 83.759 61.19 ;
      RECT MASK 1 84.097 61.09 90.377 61.19 ;
      RECT MASK 1 90.715 61.09 96.995 61.19 ;
      RECT MASK 1 97.333 61.09 103.613 61.19 ;
      RECT MASK 1 103.951 61.09 110.231 61.19 ;
      RECT MASK 1 111.044 61.4475 129.1315 61.5475 ;
      RECT MASK 1 4.672 61.465 10.96 61.565 ;
      RECT MASK 1 11.29 61.465 17.578 61.565 ;
      RECT MASK 1 17.908 61.465 24.196 61.565 ;
      RECT MASK 1 24.526 61.465 30.814 61.565 ;
      RECT MASK 1 31.144 61.465 37.432 61.565 ;
      RECT MASK 1 37.762 61.465 44.05 61.565 ;
      RECT MASK 1 44.38 61.465 50.668 61.565 ;
      RECT MASK 1 50.998 61.465 57.286 61.565 ;
      RECT MASK 1 57.616 61.465 63.904 61.565 ;
      RECT MASK 1 64.234 61.465 70.522 61.565 ;
      RECT MASK 1 70.852 61.465 77.14 61.565 ;
      RECT MASK 1 77.47 61.465 83.758 61.565 ;
      RECT MASK 1 84.088 61.465 90.376 61.565 ;
      RECT MASK 1 90.706 61.465 96.994 61.565 ;
      RECT MASK 1 97.324 61.465 103.612 61.565 ;
      RECT MASK 1 103.942 61.465 110.23 61.565 ;
      RECT MASK 1 4.672 61.835 10.96 61.935 ;
      RECT MASK 1 11.29 61.835 17.578 61.935 ;
      RECT MASK 1 17.908 61.835 24.196 61.935 ;
      RECT MASK 1 24.526 61.835 30.814 61.935 ;
      RECT MASK 1 31.144 61.835 37.432 61.935 ;
      RECT MASK 1 37.762 61.835 44.05 61.935 ;
      RECT MASK 1 44.38 61.835 50.668 61.935 ;
      RECT MASK 1 50.998 61.835 57.286 61.935 ;
      RECT MASK 1 57.616 61.835 63.904 61.935 ;
      RECT MASK 1 64.234 61.835 70.522 61.935 ;
      RECT MASK 1 70.852 61.835 77.14 61.935 ;
      RECT MASK 1 77.47 61.835 83.758 61.935 ;
      RECT MASK 1 84.088 61.835 90.376 61.935 ;
      RECT MASK 1 90.706 61.835 96.994 61.935 ;
      RECT MASK 1 97.324 61.835 103.612 61.935 ;
      RECT MASK 1 103.942 61.835 110.23 61.935 ;
      RECT MASK 1 111.044 61.9625 127.58 62.0625 ;
      RECT MASK 1 4.681 62.21 10.961 62.31 ;
      RECT MASK 1 11.299 62.21 17.579 62.31 ;
      RECT MASK 1 17.917 62.21 24.197 62.31 ;
      RECT MASK 1 24.535 62.21 30.815 62.31 ;
      RECT MASK 1 31.153 62.21 37.433 62.31 ;
      RECT MASK 1 37.771 62.21 44.051 62.31 ;
      RECT MASK 1 44.389 62.21 50.669 62.31 ;
      RECT MASK 1 51.007 62.21 57.287 62.31 ;
      RECT MASK 1 57.625 62.21 63.905 62.31 ;
      RECT MASK 1 64.243 62.21 70.523 62.31 ;
      RECT MASK 1 70.861 62.21 77.141 62.31 ;
      RECT MASK 1 77.479 62.21 83.759 62.31 ;
      RECT MASK 1 84.097 62.21 90.377 62.31 ;
      RECT MASK 1 90.715 62.21 96.995 62.31 ;
      RECT MASK 1 97.333 62.21 103.613 62.31 ;
      RECT MASK 1 103.951 62.21 110.231 62.31 ;
      RECT MASK 1 111.044 62.2825 129.1315 62.5325 ;
      RECT MASK 1 4.672 62.585 10.96 62.685 ;
      RECT MASK 1 11.29 62.585 17.578 62.685 ;
      RECT MASK 1 17.908 62.585 24.196 62.685 ;
      RECT MASK 1 24.526 62.585 30.814 62.685 ;
      RECT MASK 1 31.144 62.585 37.432 62.685 ;
      RECT MASK 1 37.762 62.585 44.05 62.685 ;
      RECT MASK 1 44.38 62.585 50.668 62.685 ;
      RECT MASK 1 50.998 62.585 57.286 62.685 ;
      RECT MASK 1 57.616 62.585 63.904 62.685 ;
      RECT MASK 1 64.234 62.585 70.522 62.685 ;
      RECT MASK 1 70.852 62.585 77.14 62.685 ;
      RECT MASK 1 77.47 62.585 83.758 62.685 ;
      RECT MASK 1 84.088 62.585 90.376 62.685 ;
      RECT MASK 1 90.706 62.585 96.994 62.685 ;
      RECT MASK 1 97.324 62.585 103.612 62.685 ;
      RECT MASK 1 103.942 62.585 110.23 62.685 ;
      RECT MASK 1 111.044 62.7975 129.1315 62.8975 ;
      RECT MASK 1 4.672 62.955 10.96 63.055 ;
      RECT MASK 1 11.29 62.955 17.578 63.055 ;
      RECT MASK 1 17.908 62.955 24.196 63.055 ;
      RECT MASK 1 24.526 62.955 30.814 63.055 ;
      RECT MASK 1 31.144 62.955 37.432 63.055 ;
      RECT MASK 1 37.762 62.955 44.05 63.055 ;
      RECT MASK 1 44.38 62.955 50.668 63.055 ;
      RECT MASK 1 50.998 62.955 57.286 63.055 ;
      RECT MASK 1 57.616 62.955 63.904 63.055 ;
      RECT MASK 1 64.234 62.955 70.522 63.055 ;
      RECT MASK 1 70.852 62.955 77.14 63.055 ;
      RECT MASK 1 77.47 62.955 83.758 63.055 ;
      RECT MASK 1 84.088 62.955 90.376 63.055 ;
      RECT MASK 1 90.706 62.955 96.994 63.055 ;
      RECT MASK 1 97.324 62.955 103.612 63.055 ;
      RECT MASK 1 103.942 62.955 110.23 63.055 ;
      RECT MASK 1 111.044 63.3125 127.58 63.4125 ;
      RECT MASK 1 4.681 63.33 10.961 63.43 ;
      RECT MASK 1 11.299 63.33 17.579 63.43 ;
      RECT MASK 1 17.917 63.33 24.197 63.43 ;
      RECT MASK 1 24.535 63.33 30.815 63.43 ;
      RECT MASK 1 31.153 63.33 37.433 63.43 ;
      RECT MASK 1 37.771 63.33 44.051 63.43 ;
      RECT MASK 1 44.389 63.33 50.669 63.43 ;
      RECT MASK 1 51.007 63.33 57.287 63.43 ;
      RECT MASK 1 57.625 63.33 63.905 63.43 ;
      RECT MASK 1 64.243 63.33 70.523 63.43 ;
      RECT MASK 1 70.861 63.33 77.141 63.43 ;
      RECT MASK 1 77.479 63.33 83.759 63.43 ;
      RECT MASK 1 84.097 63.33 90.377 63.43 ;
      RECT MASK 1 90.715 63.33 96.995 63.43 ;
      RECT MASK 1 97.333 63.33 103.613 63.43 ;
      RECT MASK 1 103.951 63.33 110.231 63.43 ;
      RECT MASK 1 117.268 63.6325 129.1315 63.8825 ;
      RECT MASK 1 117.268 64.1775 129.1315 64.2775 ;
      RECT MASK 1 111.044 64.6925 127.58 64.7925 ;
      RECT MASK 1 4.681 64.97 10.961 65.07 ;
      RECT MASK 1 11.299 64.97 17.579 65.07 ;
      RECT MASK 1 17.917 64.97 24.197 65.07 ;
      RECT MASK 1 24.535 64.97 30.815 65.07 ;
      RECT MASK 1 31.153 64.97 37.433 65.07 ;
      RECT MASK 1 37.771 64.97 44.051 65.07 ;
      RECT MASK 1 44.389 64.97 50.669 65.07 ;
      RECT MASK 1 51.007 64.97 57.287 65.07 ;
      RECT MASK 1 57.625 64.97 63.905 65.07 ;
      RECT MASK 1 64.243 64.97 70.523 65.07 ;
      RECT MASK 1 70.861 64.97 77.141 65.07 ;
      RECT MASK 1 77.479 64.97 83.759 65.07 ;
      RECT MASK 1 84.097 64.97 90.377 65.07 ;
      RECT MASK 1 90.715 64.97 96.995 65.07 ;
      RECT MASK 1 97.333 64.97 103.613 65.07 ;
      RECT MASK 1 103.951 64.97 110.231 65.07 ;
      RECT MASK 1 111.044 65.0125 129.1315 65.2625 ;
      RECT MASK 1 4.672 65.345 10.96 65.445 ;
      RECT MASK 1 11.29 65.345 17.578 65.445 ;
      RECT MASK 1 17.908 65.345 24.196 65.445 ;
      RECT MASK 1 24.526 65.345 30.814 65.445 ;
      RECT MASK 1 31.144 65.345 37.432 65.445 ;
      RECT MASK 1 37.762 65.345 44.05 65.445 ;
      RECT MASK 1 44.38 65.345 50.668 65.445 ;
      RECT MASK 1 50.998 65.345 57.286 65.445 ;
      RECT MASK 1 57.616 65.345 63.904 65.445 ;
      RECT MASK 1 64.234 65.345 70.522 65.445 ;
      RECT MASK 1 70.852 65.345 77.14 65.445 ;
      RECT MASK 1 77.47 65.345 83.758 65.445 ;
      RECT MASK 1 84.088 65.345 90.376 65.445 ;
      RECT MASK 1 90.706 65.345 96.994 65.445 ;
      RECT MASK 1 97.324 65.345 103.612 65.445 ;
      RECT MASK 1 103.942 65.345 110.23 65.445 ;
      RECT MASK 1 111.044 65.5275 129.1315 65.6275 ;
      RECT MASK 1 4.672 65.715 10.96 65.815 ;
      RECT MASK 1 11.29 65.715 17.578 65.815 ;
      RECT MASK 1 17.908 65.715 24.196 65.815 ;
      RECT MASK 1 24.526 65.715 30.814 65.815 ;
      RECT MASK 1 31.144 65.715 37.432 65.815 ;
      RECT MASK 1 37.762 65.715 44.05 65.815 ;
      RECT MASK 1 44.38 65.715 50.668 65.815 ;
      RECT MASK 1 50.998 65.715 57.286 65.815 ;
      RECT MASK 1 57.616 65.715 63.904 65.815 ;
      RECT MASK 1 64.234 65.715 70.522 65.815 ;
      RECT MASK 1 70.852 65.715 77.14 65.815 ;
      RECT MASK 1 77.47 65.715 83.758 65.815 ;
      RECT MASK 1 84.088 65.715 90.376 65.815 ;
      RECT MASK 1 90.706 65.715 96.994 65.815 ;
      RECT MASK 1 97.324 65.715 103.612 65.815 ;
      RECT MASK 1 103.942 65.715 110.23 65.815 ;
      RECT MASK 1 111.044 66.0425 127.58 66.1425 ;
      RECT MASK 1 4.681 66.09 10.961 66.19 ;
      RECT MASK 1 11.299 66.09 17.579 66.19 ;
      RECT MASK 1 17.917 66.09 24.197 66.19 ;
      RECT MASK 1 24.535 66.09 30.815 66.19 ;
      RECT MASK 1 31.153 66.09 37.433 66.19 ;
      RECT MASK 1 37.771 66.09 44.051 66.19 ;
      RECT MASK 1 44.389 66.09 50.669 66.19 ;
      RECT MASK 1 51.007 66.09 57.287 66.19 ;
      RECT MASK 1 57.625 66.09 63.905 66.19 ;
      RECT MASK 1 64.243 66.09 70.523 66.19 ;
      RECT MASK 1 70.861 66.09 77.141 66.19 ;
      RECT MASK 1 77.479 66.09 83.759 66.19 ;
      RECT MASK 1 84.097 66.09 90.377 66.19 ;
      RECT MASK 1 90.715 66.09 96.995 66.19 ;
      RECT MASK 1 97.333 66.09 103.613 66.19 ;
      RECT MASK 1 103.951 66.09 110.231 66.19 ;
      RECT MASK 1 111.044 66.3625 129.1315 66.6125 ;
      RECT MASK 1 4.672 66.465 10.96 66.565 ;
      RECT MASK 1 11.29 66.465 17.578 66.565 ;
      RECT MASK 1 17.908 66.465 24.196 66.565 ;
      RECT MASK 1 24.526 66.465 30.814 66.565 ;
      RECT MASK 1 31.144 66.465 37.432 66.565 ;
      RECT MASK 1 37.762 66.465 44.05 66.565 ;
      RECT MASK 1 44.38 66.465 50.668 66.565 ;
      RECT MASK 1 50.998 66.465 57.286 66.565 ;
      RECT MASK 1 57.616 66.465 63.904 66.565 ;
      RECT MASK 1 64.234 66.465 70.522 66.565 ;
      RECT MASK 1 70.852 66.465 77.14 66.565 ;
      RECT MASK 1 77.47 66.465 83.758 66.565 ;
      RECT MASK 1 84.088 66.465 90.376 66.565 ;
      RECT MASK 1 90.706 66.465 96.994 66.565 ;
      RECT MASK 1 97.324 66.465 103.612 66.565 ;
      RECT MASK 1 103.942 66.465 110.23 66.565 ;
      RECT MASK 1 4.672 66.835 10.96 66.935 ;
      RECT MASK 1 11.29 66.835 17.578 66.935 ;
      RECT MASK 1 17.908 66.835 24.196 66.935 ;
      RECT MASK 1 24.526 66.835 30.814 66.935 ;
      RECT MASK 1 31.144 66.835 37.432 66.935 ;
      RECT MASK 1 37.762 66.835 44.05 66.935 ;
      RECT MASK 1 44.38 66.835 50.668 66.935 ;
      RECT MASK 1 50.998 66.835 57.286 66.935 ;
      RECT MASK 1 57.616 66.835 63.904 66.935 ;
      RECT MASK 1 64.234 66.835 70.522 66.935 ;
      RECT MASK 1 70.852 66.835 77.14 66.935 ;
      RECT MASK 1 77.47 66.835 83.758 66.935 ;
      RECT MASK 1 84.088 66.835 90.376 66.935 ;
      RECT MASK 1 90.706 66.835 96.994 66.935 ;
      RECT MASK 1 97.324 66.835 103.612 66.935 ;
      RECT MASK 1 103.942 66.835 110.23 66.935 ;
      RECT MASK 1 111.044 66.8775 129.1315 66.9775 ;
      RECT MASK 1 4.681 67.21 10.961 67.31 ;
      RECT MASK 1 11.299 67.21 17.579 67.31 ;
      RECT MASK 1 17.917 67.21 24.197 67.31 ;
      RECT MASK 1 24.535 67.21 30.815 67.31 ;
      RECT MASK 1 31.153 67.21 37.433 67.31 ;
      RECT MASK 1 37.771 67.21 44.051 67.31 ;
      RECT MASK 1 44.389 67.21 50.669 67.31 ;
      RECT MASK 1 51.007 67.21 57.287 67.31 ;
      RECT MASK 1 57.625 67.21 63.905 67.31 ;
      RECT MASK 1 64.243 67.21 70.523 67.31 ;
      RECT MASK 1 70.861 67.21 77.141 67.31 ;
      RECT MASK 1 77.479 67.21 83.759 67.31 ;
      RECT MASK 1 84.097 67.21 90.377 67.31 ;
      RECT MASK 1 90.715 67.21 96.995 67.31 ;
      RECT MASK 1 97.333 67.21 103.613 67.31 ;
      RECT MASK 1 103.951 67.21 110.231 67.31 ;
      RECT MASK 1 111.044 67.3925 127.58 67.4925 ;
      RECT MASK 1 4.672 67.585 10.96 67.685 ;
      RECT MASK 1 11.29 67.585 17.578 67.685 ;
      RECT MASK 1 17.908 67.585 24.196 67.685 ;
      RECT MASK 1 24.526 67.585 30.814 67.685 ;
      RECT MASK 1 31.144 67.585 37.432 67.685 ;
      RECT MASK 1 37.762 67.585 44.05 67.685 ;
      RECT MASK 1 44.38 67.585 50.668 67.685 ;
      RECT MASK 1 50.998 67.585 57.286 67.685 ;
      RECT MASK 1 57.616 67.585 63.904 67.685 ;
      RECT MASK 1 64.234 67.585 70.522 67.685 ;
      RECT MASK 1 70.852 67.585 77.14 67.685 ;
      RECT MASK 1 77.47 67.585 83.758 67.685 ;
      RECT MASK 1 84.088 67.585 90.376 67.685 ;
      RECT MASK 1 90.706 67.585 96.994 67.685 ;
      RECT MASK 1 97.324 67.585 103.612 67.685 ;
      RECT MASK 1 103.942 67.585 110.23 67.685 ;
      RECT MASK 1 111.044 67.7125 129.1315 67.9625 ;
      RECT MASK 1 4.672 67.955 10.96 68.055 ;
      RECT MASK 1 11.29 67.955 17.578 68.055 ;
      RECT MASK 1 17.908 67.955 24.196 68.055 ;
      RECT MASK 1 24.526 67.955 30.814 68.055 ;
      RECT MASK 1 31.144 67.955 37.432 68.055 ;
      RECT MASK 1 37.762 67.955 44.05 68.055 ;
      RECT MASK 1 44.38 67.955 50.668 68.055 ;
      RECT MASK 1 50.998 67.955 57.286 68.055 ;
      RECT MASK 1 57.616 67.955 63.904 68.055 ;
      RECT MASK 1 64.234 67.955 70.522 68.055 ;
      RECT MASK 1 70.852 67.955 77.14 68.055 ;
      RECT MASK 1 77.47 67.955 83.758 68.055 ;
      RECT MASK 1 84.088 67.955 90.376 68.055 ;
      RECT MASK 1 90.706 67.955 96.994 68.055 ;
      RECT MASK 1 97.324 67.955 103.612 68.055 ;
      RECT MASK 1 103.942 67.955 110.23 68.055 ;
      RECT MASK 1 111.044 68.2275 129.1315 68.3275 ;
      RECT MASK 1 4.681 68.33 10.961 68.43 ;
      RECT MASK 1 11.299 68.33 17.579 68.43 ;
      RECT MASK 1 17.917 68.33 24.197 68.43 ;
      RECT MASK 1 24.535 68.33 30.815 68.43 ;
      RECT MASK 1 31.153 68.33 37.433 68.43 ;
      RECT MASK 1 37.771 68.33 44.051 68.43 ;
      RECT MASK 1 44.389 68.33 50.669 68.43 ;
      RECT MASK 1 51.007 68.33 57.287 68.43 ;
      RECT MASK 1 57.625 68.33 63.905 68.43 ;
      RECT MASK 1 64.243 68.33 70.523 68.43 ;
      RECT MASK 1 70.861 68.33 77.141 68.43 ;
      RECT MASK 1 77.479 68.33 83.759 68.43 ;
      RECT MASK 1 84.097 68.33 90.377 68.43 ;
      RECT MASK 1 90.715 68.33 96.995 68.43 ;
      RECT MASK 1 97.333 68.33 103.613 68.43 ;
      RECT MASK 1 103.951 68.33 110.231 68.43 ;
      RECT MASK 1 4.672 68.705 10.96 68.805 ;
      RECT MASK 1 11.29 68.705 17.578 68.805 ;
      RECT MASK 1 17.908 68.705 24.196 68.805 ;
      RECT MASK 1 24.526 68.705 30.814 68.805 ;
      RECT MASK 1 31.144 68.705 37.432 68.805 ;
      RECT MASK 1 37.762 68.705 44.05 68.805 ;
      RECT MASK 1 44.38 68.705 50.668 68.805 ;
      RECT MASK 1 50.998 68.705 57.286 68.805 ;
      RECT MASK 1 57.616 68.705 63.904 68.805 ;
      RECT MASK 1 64.234 68.705 70.522 68.805 ;
      RECT MASK 1 70.852 68.705 77.14 68.805 ;
      RECT MASK 1 77.47 68.705 83.758 68.805 ;
      RECT MASK 1 84.088 68.705 90.376 68.805 ;
      RECT MASK 1 90.706 68.705 96.994 68.805 ;
      RECT MASK 1 97.324 68.705 103.612 68.805 ;
      RECT MASK 1 103.942 68.705 110.23 68.805 ;
      RECT MASK 1 111.044 68.7425 127.58 68.8425 ;
      RECT MASK 1 111.044 69.0625 129.1315 69.3125 ;
      RECT MASK 1 4.672 69.075 10.96 69.175 ;
      RECT MASK 1 11.29 69.075 17.578 69.175 ;
      RECT MASK 1 17.908 69.075 24.196 69.175 ;
      RECT MASK 1 24.526 69.075 30.814 69.175 ;
      RECT MASK 1 31.144 69.075 37.432 69.175 ;
      RECT MASK 1 37.762 69.075 44.05 69.175 ;
      RECT MASK 1 44.38 69.075 50.668 69.175 ;
      RECT MASK 1 50.998 69.075 57.286 69.175 ;
      RECT MASK 1 57.616 69.075 63.904 69.175 ;
      RECT MASK 1 64.234 69.075 70.522 69.175 ;
      RECT MASK 1 70.852 69.075 77.14 69.175 ;
      RECT MASK 1 77.47 69.075 83.758 69.175 ;
      RECT MASK 1 84.088 69.075 90.376 69.175 ;
      RECT MASK 1 90.706 69.075 96.994 69.175 ;
      RECT MASK 1 97.324 69.075 103.612 69.175 ;
      RECT MASK 1 103.942 69.075 110.23 69.175 ;
      RECT MASK 1 4.681 69.45 10.961 69.55 ;
      RECT MASK 1 11.299 69.45 17.579 69.55 ;
      RECT MASK 1 17.917 69.45 24.197 69.55 ;
      RECT MASK 1 24.535 69.45 30.815 69.55 ;
      RECT MASK 1 31.153 69.45 37.433 69.55 ;
      RECT MASK 1 37.771 69.45 44.051 69.55 ;
      RECT MASK 1 44.389 69.45 50.669 69.55 ;
      RECT MASK 1 51.007 69.45 57.287 69.55 ;
      RECT MASK 1 57.625 69.45 63.905 69.55 ;
      RECT MASK 1 64.243 69.45 70.523 69.55 ;
      RECT MASK 1 70.861 69.45 77.141 69.55 ;
      RECT MASK 1 77.479 69.45 83.759 69.55 ;
      RECT MASK 1 84.097 69.45 90.377 69.55 ;
      RECT MASK 1 90.715 69.45 96.995 69.55 ;
      RECT MASK 1 97.333 69.45 103.613 69.55 ;
      RECT MASK 1 103.951 69.45 110.231 69.55 ;
      RECT MASK 1 111.044 69.5775 129.1315 69.6775 ;
      RECT MASK 1 113.0865 70.8925 127.58 71.1425 ;
      RECT MASK 1 4.681 71.09 10.961 71.19 ;
      RECT MASK 1 11.299 71.09 17.579 71.19 ;
      RECT MASK 1 17.917 71.09 24.197 71.19 ;
      RECT MASK 1 24.535 71.09 30.815 71.19 ;
      RECT MASK 1 31.153 71.09 37.433 71.19 ;
      RECT MASK 1 37.771 71.09 44.051 71.19 ;
      RECT MASK 1 44.389 71.09 50.669 71.19 ;
      RECT MASK 1 51.007 71.09 57.287 71.19 ;
      RECT MASK 1 57.625 71.09 63.905 71.19 ;
      RECT MASK 1 64.243 71.09 70.523 71.19 ;
      RECT MASK 1 70.861 71.09 77.141 71.19 ;
      RECT MASK 1 77.479 71.09 83.759 71.19 ;
      RECT MASK 1 84.097 71.09 90.377 71.19 ;
      RECT MASK 1 90.715 71.09 96.995 71.19 ;
      RECT MASK 1 97.333 71.09 103.613 71.19 ;
      RECT MASK 1 103.951 71.09 110.231 71.19 ;
      RECT MASK 1 111.044 71.325 129.1315 71.385 ;
      RECT MASK 1 4.672 71.465 10.96 71.565 ;
      RECT MASK 1 11.29 71.465 17.578 71.565 ;
      RECT MASK 1 17.908 71.465 24.196 71.565 ;
      RECT MASK 1 24.526 71.465 30.814 71.565 ;
      RECT MASK 1 31.144 71.465 37.432 71.565 ;
      RECT MASK 1 37.762 71.465 44.05 71.565 ;
      RECT MASK 1 44.38 71.465 50.668 71.565 ;
      RECT MASK 1 50.998 71.465 57.286 71.565 ;
      RECT MASK 1 57.616 71.465 63.904 71.565 ;
      RECT MASK 1 64.234 71.465 70.522 71.565 ;
      RECT MASK 1 70.852 71.465 77.14 71.565 ;
      RECT MASK 1 77.47 71.465 83.758 71.565 ;
      RECT MASK 1 84.088 71.465 90.376 71.565 ;
      RECT MASK 1 90.706 71.465 96.994 71.565 ;
      RECT MASK 1 97.324 71.465 103.612 71.565 ;
      RECT MASK 1 103.942 71.465 110.23 71.565 ;
      RECT MASK 1 111.044 71.5675 129.1315 71.8175 ;
      RECT MASK 1 4.672 71.835 10.96 71.935 ;
      RECT MASK 1 11.29 71.835 17.578 71.935 ;
      RECT MASK 1 17.908 71.835 24.196 71.935 ;
      RECT MASK 1 24.526 71.835 30.814 71.935 ;
      RECT MASK 1 31.144 71.835 37.432 71.935 ;
      RECT MASK 1 37.762 71.835 44.05 71.935 ;
      RECT MASK 1 44.38 71.835 50.668 71.935 ;
      RECT MASK 1 50.998 71.835 57.286 71.935 ;
      RECT MASK 1 57.616 71.835 63.904 71.935 ;
      RECT MASK 1 64.234 71.835 70.522 71.935 ;
      RECT MASK 1 70.852 71.835 77.14 71.935 ;
      RECT MASK 1 77.47 71.835 83.758 71.935 ;
      RECT MASK 1 84.088 71.835 90.376 71.935 ;
      RECT MASK 1 90.706 71.835 96.994 71.935 ;
      RECT MASK 1 97.324 71.835 103.612 71.935 ;
      RECT MASK 1 103.942 71.835 110.23 71.935 ;
      RECT MASK 1 4.681 72.21 10.961 72.31 ;
      RECT MASK 1 11.299 72.21 17.579 72.31 ;
      RECT MASK 1 17.917 72.21 24.197 72.31 ;
      RECT MASK 1 24.535 72.21 30.815 72.31 ;
      RECT MASK 1 31.153 72.21 37.433 72.31 ;
      RECT MASK 1 37.771 72.21 44.051 72.31 ;
      RECT MASK 1 44.389 72.21 50.669 72.31 ;
      RECT MASK 1 51.007 72.21 57.287 72.31 ;
      RECT MASK 1 57.625 72.21 63.905 72.31 ;
      RECT MASK 1 64.243 72.21 70.523 72.31 ;
      RECT MASK 1 70.861 72.21 77.141 72.31 ;
      RECT MASK 1 77.479 72.21 83.759 72.31 ;
      RECT MASK 1 84.097 72.21 90.377 72.31 ;
      RECT MASK 1 90.715 72.21 96.995 72.31 ;
      RECT MASK 1 97.333 72.21 103.613 72.31 ;
      RECT MASK 1 103.951 72.21 110.231 72.31 ;
      RECT MASK 1 111.0245 72.345 129.1315 72.465 ;
      RECT MASK 1 4.672 72.585 10.96 72.685 ;
      RECT MASK 1 11.29 72.585 17.578 72.685 ;
      RECT MASK 1 17.908 72.585 24.196 72.685 ;
      RECT MASK 1 24.526 72.585 30.814 72.685 ;
      RECT MASK 1 31.144 72.585 37.432 72.685 ;
      RECT MASK 1 37.762 72.585 44.05 72.685 ;
      RECT MASK 1 44.38 72.585 50.668 72.685 ;
      RECT MASK 1 50.998 72.585 57.286 72.685 ;
      RECT MASK 1 57.616 72.585 63.904 72.685 ;
      RECT MASK 1 64.234 72.585 70.522 72.685 ;
      RECT MASK 1 70.852 72.585 77.14 72.685 ;
      RECT MASK 1 77.47 72.585 83.758 72.685 ;
      RECT MASK 1 84.088 72.585 90.376 72.685 ;
      RECT MASK 1 90.706 72.585 96.994 72.685 ;
      RECT MASK 1 97.324 72.585 103.612 72.685 ;
      RECT MASK 1 103.942 72.585 110.23 72.685 ;
      RECT MASK 1 113.84 72.845 114.583 72.965 ;
      RECT MASK 1 4.672 72.955 10.96 73.055 ;
      RECT MASK 1 11.29 72.955 17.578 73.055 ;
      RECT MASK 1 17.908 72.955 24.196 73.055 ;
      RECT MASK 1 24.526 72.955 30.814 73.055 ;
      RECT MASK 1 31.144 72.955 37.432 73.055 ;
      RECT MASK 1 37.762 72.955 44.05 73.055 ;
      RECT MASK 1 44.38 72.955 50.668 73.055 ;
      RECT MASK 1 50.998 72.955 57.286 73.055 ;
      RECT MASK 1 57.616 72.955 63.904 73.055 ;
      RECT MASK 1 64.234 72.955 70.522 73.055 ;
      RECT MASK 1 70.852 72.955 77.14 73.055 ;
      RECT MASK 1 77.47 72.955 83.758 73.055 ;
      RECT MASK 1 84.088 72.955 90.376 73.055 ;
      RECT MASK 1 90.706 72.955 96.994 73.055 ;
      RECT MASK 1 97.324 72.955 103.612 73.055 ;
      RECT MASK 1 103.942 72.955 110.23 73.055 ;
      RECT MASK 1 115.506 73.305 126.992 73.425 ;
      RECT MASK 1 4.681 73.33 10.961 73.43 ;
      RECT MASK 1 11.299 73.33 17.579 73.43 ;
      RECT MASK 1 17.917 73.33 24.197 73.43 ;
      RECT MASK 1 24.535 73.33 30.815 73.43 ;
      RECT MASK 1 31.153 73.33 37.433 73.43 ;
      RECT MASK 1 37.771 73.33 44.051 73.43 ;
      RECT MASK 1 44.389 73.33 50.669 73.43 ;
      RECT MASK 1 51.007 73.33 57.287 73.43 ;
      RECT MASK 1 57.625 73.33 63.905 73.43 ;
      RECT MASK 1 64.243 73.33 70.523 73.43 ;
      RECT MASK 1 70.861 73.33 77.141 73.43 ;
      RECT MASK 1 77.479 73.33 83.759 73.43 ;
      RECT MASK 1 84.097 73.33 90.377 73.43 ;
      RECT MASK 1 90.715 73.33 96.995 73.43 ;
      RECT MASK 1 97.333 73.33 103.613 73.43 ;
      RECT MASK 1 103.951 73.33 110.231 73.43 ;
      RECT MASK 1 4.672 73.705 10.96 73.805 ;
      RECT MASK 1 11.29 73.705 17.578 73.805 ;
      RECT MASK 1 17.908 73.705 24.196 73.805 ;
      RECT MASK 1 24.526 73.705 30.814 73.805 ;
      RECT MASK 1 31.144 73.705 37.432 73.805 ;
      RECT MASK 1 37.762 73.705 44.05 73.805 ;
      RECT MASK 1 44.38 73.705 50.668 73.805 ;
      RECT MASK 1 50.998 73.705 57.286 73.805 ;
      RECT MASK 1 57.616 73.705 63.904 73.805 ;
      RECT MASK 1 64.234 73.705 70.522 73.805 ;
      RECT MASK 1 70.852 73.705 77.14 73.805 ;
      RECT MASK 1 77.47 73.705 83.758 73.805 ;
      RECT MASK 1 84.088 73.705 90.376 73.805 ;
      RECT MASK 1 90.706 73.705 96.994 73.805 ;
      RECT MASK 1 97.324 73.705 103.612 73.805 ;
      RECT MASK 1 103.942 73.705 110.23 73.805 ;
      RECT MASK 1 116.163 74 126.333 74.2 ;
      RECT MASK 1 4.672 74.075 10.96 74.175 ;
      RECT MASK 1 11.29 74.075 17.578 74.175 ;
      RECT MASK 1 17.908 74.075 24.196 74.175 ;
      RECT MASK 1 24.526 74.075 30.814 74.175 ;
      RECT MASK 1 31.144 74.075 37.432 74.175 ;
      RECT MASK 1 37.762 74.075 44.05 74.175 ;
      RECT MASK 1 44.38 74.075 50.668 74.175 ;
      RECT MASK 1 50.998 74.075 57.286 74.175 ;
      RECT MASK 1 57.616 74.075 63.904 74.175 ;
      RECT MASK 1 64.234 74.075 70.522 74.175 ;
      RECT MASK 1 70.852 74.075 77.14 74.175 ;
      RECT MASK 1 77.47 74.075 83.758 74.175 ;
      RECT MASK 1 84.088 74.075 90.376 74.175 ;
      RECT MASK 1 90.706 74.075 96.994 74.175 ;
      RECT MASK 1 97.324 74.075 103.612 74.175 ;
      RECT MASK 1 103.942 74.075 110.23 74.175 ;
      RECT MASK 1 4.681 74.45 10.961 74.55 ;
      RECT MASK 1 11.299 74.45 17.579 74.55 ;
      RECT MASK 1 17.917 74.45 24.197 74.55 ;
      RECT MASK 1 24.535 74.45 30.815 74.55 ;
      RECT MASK 1 31.153 74.45 37.433 74.55 ;
      RECT MASK 1 37.771 74.45 44.051 74.55 ;
      RECT MASK 1 44.389 74.45 50.669 74.55 ;
      RECT MASK 1 51.007 74.45 57.287 74.55 ;
      RECT MASK 1 57.625 74.45 63.905 74.55 ;
      RECT MASK 1 64.243 74.45 70.523 74.55 ;
      RECT MASK 1 70.861 74.45 77.141 74.55 ;
      RECT MASK 1 77.479 74.45 83.759 74.55 ;
      RECT MASK 1 84.097 74.45 90.377 74.55 ;
      RECT MASK 1 90.715 74.45 96.995 74.55 ;
      RECT MASK 1 97.333 74.45 103.613 74.55 ;
      RECT MASK 1 103.951 74.45 110.231 74.55 ;
      RECT MASK 1 126.538 74.47 127.51 74.53 ;
      RECT MASK 1 116.163 74.52 126.333 74.72 ;
      RECT MASK 1 4.672 74.825 10.96 74.925 ;
      RECT MASK 1 11.29 74.825 17.578 74.925 ;
      RECT MASK 1 17.908 74.825 24.196 74.925 ;
      RECT MASK 1 24.526 74.825 30.814 74.925 ;
      RECT MASK 1 31.144 74.825 37.432 74.925 ;
      RECT MASK 1 37.762 74.825 44.05 74.925 ;
      RECT MASK 1 44.38 74.825 50.668 74.925 ;
      RECT MASK 1 50.998 74.825 57.286 74.925 ;
      RECT MASK 1 57.616 74.825 63.904 74.925 ;
      RECT MASK 1 64.234 74.825 70.522 74.925 ;
      RECT MASK 1 70.852 74.825 77.14 74.925 ;
      RECT MASK 1 77.47 74.825 83.758 74.925 ;
      RECT MASK 1 84.088 74.825 90.376 74.925 ;
      RECT MASK 1 90.706 74.825 96.994 74.925 ;
      RECT MASK 1 97.324 74.825 103.612 74.925 ;
      RECT MASK 1 103.942 74.825 110.23 74.925 ;
      RECT MASK 1 116.218 75.11 126.339 75.17 ;
      RECT MASK 1 4.672 75.195 10.96 75.295 ;
      RECT MASK 1 11.29 75.195 17.578 75.295 ;
      RECT MASK 1 17.908 75.195 24.196 75.295 ;
      RECT MASK 1 24.526 75.195 30.814 75.295 ;
      RECT MASK 1 31.144 75.195 37.432 75.295 ;
      RECT MASK 1 37.762 75.195 44.05 75.295 ;
      RECT MASK 1 44.38 75.195 50.668 75.295 ;
      RECT MASK 1 50.998 75.195 57.286 75.295 ;
      RECT MASK 1 57.616 75.195 63.904 75.295 ;
      RECT MASK 1 64.234 75.195 70.522 75.295 ;
      RECT MASK 1 70.852 75.195 77.14 75.295 ;
      RECT MASK 1 77.47 75.195 83.758 75.295 ;
      RECT MASK 1 84.088 75.195 90.376 75.295 ;
      RECT MASK 1 90.706 75.195 96.994 75.295 ;
      RECT MASK 1 97.324 75.195 103.612 75.295 ;
      RECT MASK 1 103.942 75.195 110.23 75.295 ;
      RECT MASK 1 126.538 75.25 127.51 75.31 ;
      RECT MASK 1 116.162 75.56 126.332 75.76 ;
      RECT MASK 1 4.681 75.57 10.961 75.67 ;
      RECT MASK 1 11.299 75.57 17.579 75.67 ;
      RECT MASK 1 17.917 75.57 24.197 75.67 ;
      RECT MASK 1 24.535 75.57 30.815 75.67 ;
      RECT MASK 1 31.153 75.57 37.433 75.67 ;
      RECT MASK 1 37.771 75.57 44.051 75.67 ;
      RECT MASK 1 44.389 75.57 50.669 75.67 ;
      RECT MASK 1 51.007 75.57 57.287 75.67 ;
      RECT MASK 1 57.625 75.57 63.905 75.67 ;
      RECT MASK 1 64.243 75.57 70.523 75.67 ;
      RECT MASK 1 70.861 75.57 77.141 75.67 ;
      RECT MASK 1 77.479 75.57 83.759 75.67 ;
      RECT MASK 1 84.097 75.57 90.377 75.67 ;
      RECT MASK 1 90.715 75.57 96.995 75.67 ;
      RECT MASK 1 97.333 75.57 103.613 75.67 ;
      RECT MASK 1 103.951 75.57 110.231 75.67 ;
      RECT MASK 1 126.538 76.03 127.51 76.09 ;
      RECT MASK 1 116.163 76.08 126.333 76.28 ;
      RECT MASK 1 116.218 76.655 126.339 76.715 ;
      RECT MASK 1 126.538 76.81 127.51 76.87 ;
      RECT MASK 1 115.515 77.12 126.969 77.32 ;
      RECT MASK 1 126.538 77.59 127.73 77.65 ;
      RECT MASK 1 0.567 77.595 114.583 77.715 ;
      RECT MASK 1 116.163 77.64 126.333 77.84 ;
      RECT MASK 1 116.218 78.24 126.339 78.3 ;
      RECT MASK 1 126.538 78.37 127.73 78.43 ;
      RECT MASK 1 6.807 78.631 109.165 78.691 ;
      RECT MASK 1 115.515 78.68 126.969 78.88 ;
      RECT MASK 1 111.1115 78.87 113.3685 78.99 ;
      RECT MASK 1 2.169 79.15 4.491 79.19 ;
      RECT MASK 1 126.538 79.15 127.73 79.21 ;
      RECT MASK 1 116.163 79.2 126.333 79.4 ;
      RECT MASK 1 6.807 79.351 109.165 79.411 ;
      RECT MASK 1 2.169 79.39 4.491 79.43 ;
      RECT MASK 1 2.169 79.63 4.491 79.67 ;
      RECT MASK 1 10.177 79.646 12.147 79.746 ;
      RECT MASK 1 16.795 79.646 18.765 79.746 ;
      RECT MASK 1 23.413 79.646 25.383 79.746 ;
      RECT MASK 1 30.031 79.646 32.001 79.746 ;
      RECT MASK 1 36.649 79.646 38.619 79.746 ;
      RECT MASK 1 43.267 79.646 45.237 79.746 ;
      RECT MASK 1 49.885 79.646 51.855 79.746 ;
      RECT MASK 1 56.503 79.646 58.473 79.746 ;
      RECT MASK 1 63.121 79.646 65.091 79.746 ;
      RECT MASK 1 69.739 79.646 71.709 79.746 ;
      RECT MASK 1 76.357 79.646 78.327 79.746 ;
      RECT MASK 1 82.975 79.646 84.945 79.746 ;
      RECT MASK 1 89.593 79.646 91.563 79.746 ;
      RECT MASK 1 96.211 79.646 98.181 79.746 ;
      RECT MASK 1 102.829 79.646 104.799 79.746 ;
      RECT MASK 1 109.447 79.646 111.9315 79.746 ;
      RECT MASK 1 2.169 79.87 4.491 79.91 ;
      RECT MASK 1 126.538 79.93 127.73 79.99 ;
      RECT MASK 1 2.169 80.11 4.491 80.15 ;
      RECT MASK 1 115.506 80.235 126.992 80.355 ;
      RECT MASK 1 2.169 80.35 4.491 80.39 ;
      RECT MASK 1 111.186 80.382 113.339 80.562 ;
      RECT MASK 1 2.169 80.59 4.491 80.63 ;
      RECT MASK 1 57.178 80.79 59.7205 80.85 ;
      RECT MASK 1 63.0635 80.79 64.425 80.85 ;
      RECT MASK 1 2.169 80.83 4.491 80.87 ;
      RECT MASK 1 6.807 81.03 109.165 81.09 ;
      RECT MASK 1 2.169 81.07 4.491 81.11 ;
      RECT MASK 1 2.169 81.31 4.491 81.35 ;
      RECT MASK 1 10.177 81.37 12.147 81.47 ;
      RECT MASK 1 16.795 81.37 18.765 81.47 ;
      RECT MASK 1 23.413 81.37 25.383 81.47 ;
      RECT MASK 1 30.031 81.37 32.001 81.47 ;
      RECT MASK 1 36.649 81.37 38.619 81.47 ;
      RECT MASK 1 43.267 81.37 45.237 81.47 ;
      RECT MASK 1 49.885 81.37 51.855 81.47 ;
      RECT MASK 1 56.503 81.37 60.88 81.47 ;
      RECT MASK 1 63.121 81.37 65.091 81.47 ;
      RECT MASK 1 69.739 81.37 71.709 81.47 ;
      RECT MASK 1 76.357 81.37 78.327 81.47 ;
      RECT MASK 1 82.975 81.37 84.945 81.47 ;
      RECT MASK 1 89.593 81.37 91.563 81.47 ;
      RECT MASK 1 96.211 81.37 98.181 81.47 ;
      RECT MASK 1 102.829 81.37 104.799 81.47 ;
      RECT MASK 1 109.447 81.37 112.735 81.47 ;
      RECT MASK 1 2.169 81.55 4.491 81.59 ;
      RECT MASK 1 6.807 81.75 109.165 81.81 ;
      RECT MASK 1 111.1115 81.75 113.3685 81.93 ;
      RECT MASK 1 2.169 81.79 4.491 81.83 ;
      RECT MASK 1 116.564 81.94 127.654 81.98 ;
      RECT MASK 1 57.178 82.023 64.425 82.083 ;
      RECT MASK 1 2.169 82.03 4.491 82.07 ;
      RECT MASK 1 116.564 82.18 127.654 82.22 ;
      RECT MASK 1 111.1115 82.2 113.3685 82.32 ;
      RECT MASK 1 7.374 82.263 7.8555 82.323 ;
      RECT MASK 1 8.536 82.263 9.0175 82.323 ;
      RECT MASK 1 9.698 82.263 10.1795 82.323 ;
      RECT MASK 1 12.83 82.263 13.3115 82.323 ;
      RECT MASK 1 13.992 82.263 14.4735 82.323 ;
      RECT MASK 1 15.154 82.263 15.6355 82.323 ;
      RECT MASK 1 16.316 82.263 16.7975 82.323 ;
      RECT MASK 1 19.448 82.263 19.9295 82.323 ;
      RECT MASK 1 20.61 82.263 21.0915 82.323 ;
      RECT MASK 1 21.772 82.263 22.2535 82.323 ;
      RECT MASK 1 22.934 82.263 23.4155 82.323 ;
      RECT MASK 1 26.066 82.263 26.5475 82.323 ;
      RECT MASK 1 27.228 82.263 27.7095 82.323 ;
      RECT MASK 1 28.39 82.263 28.8715 82.323 ;
      RECT MASK 1 29.552 82.263 30.0335 82.323 ;
      RECT MASK 1 32.684 82.263 33.1655 82.323 ;
      RECT MASK 1 33.846 82.263 34.3275 82.323 ;
      RECT MASK 1 35.008 82.263 35.4895 82.323 ;
      RECT MASK 1 36.17 82.263 36.6515 82.323 ;
      RECT MASK 1 39.302 82.263 39.7835 82.323 ;
      RECT MASK 1 40.464 82.263 40.9455 82.323 ;
      RECT MASK 1 41.626 82.263 42.1075 82.323 ;
      RECT MASK 1 42.788 82.263 43.2695 82.323 ;
      RECT MASK 1 45.92 82.263 46.4015 82.323 ;
      RECT MASK 1 47.082 82.263 47.5635 82.323 ;
      RECT MASK 1 48.244 82.263 48.7255 82.323 ;
      RECT MASK 1 49.406 82.263 49.8875 82.323 ;
      RECT MASK 1 52.538 82.263 53.0195 82.323 ;
      RECT MASK 1 53.7 82.263 54.1815 82.323 ;
      RECT MASK 1 54.862 82.263 55.3435 82.323 ;
      RECT MASK 1 56.024 82.263 56.5055 82.323 ;
      RECT MASK 1 57.178 82.263 58.9205 82.323 ;
      RECT MASK 1 59.156 82.263 59.6375 82.323 ;
      RECT MASK 1 59.8375 82.263 60.118 82.323 ;
      RECT MASK 1 60.318 82.263 60.7995 82.323 ;
      RECT MASK 1 60.9995 82.263 61.28 82.323 ;
      RECT MASK 1 61.48 82.263 61.9615 82.323 ;
      RECT MASK 1 62.1615 82.263 62.442 82.323 ;
      RECT MASK 1 62.642 82.263 63.1235 82.323 ;
      RECT MASK 1 63.3875 82.263 64.425 82.323 ;
      RECT MASK 1 65.774 82.263 66.2555 82.323 ;
      RECT MASK 1 66.936 82.263 67.4175 82.323 ;
      RECT MASK 1 68.098 82.263 68.5795 82.323 ;
      RECT MASK 1 69.26 82.263 69.7415 82.323 ;
      RECT MASK 1 72.392 82.263 72.8735 82.323 ;
      RECT MASK 1 73.554 82.263 74.0355 82.323 ;
      RECT MASK 1 74.716 82.263 75.1975 82.323 ;
      RECT MASK 1 75.878 82.263 76.3595 82.323 ;
      RECT MASK 1 79.01 82.263 79.4915 82.323 ;
      RECT MASK 1 80.172 82.263 80.6535 82.323 ;
      RECT MASK 1 81.334 82.263 81.8155 82.323 ;
      RECT MASK 1 82.496 82.263 82.9775 82.323 ;
      RECT MASK 1 85.628 82.263 86.1095 82.323 ;
      RECT MASK 1 86.79 82.263 87.2715 82.323 ;
      RECT MASK 1 87.952 82.263 88.4335 82.323 ;
      RECT MASK 1 89.114 82.263 89.5955 82.323 ;
      RECT MASK 1 92.246 82.263 92.7275 82.323 ;
      RECT MASK 1 93.408 82.263 93.8895 82.323 ;
      RECT MASK 1 94.57 82.263 95.0515 82.323 ;
      RECT MASK 1 95.732 82.263 96.2135 82.323 ;
      RECT MASK 1 98.864 82.263 99.3455 82.323 ;
      RECT MASK 1 100.026 82.263 100.5075 82.323 ;
      RECT MASK 1 101.188 82.263 101.6695 82.323 ;
      RECT MASK 1 102.35 82.263 102.8315 82.323 ;
      RECT MASK 1 105.482 82.263 105.9635 82.323 ;
      RECT MASK 1 106.644 82.263 107.1255 82.323 ;
      RECT MASK 1 107.806 82.263 108.2875 82.323 ;
      RECT MASK 1 108.968 82.263 109.4495 82.323 ;
      RECT MASK 1 2.169 82.27 4.491 82.31 ;
      RECT MASK 1 116.564 82.42 127.654 82.46 ;
      RECT MASK 1 2.169 82.51 4.491 82.55 ;
      RECT MASK 1 57.178 82.605 64.425 82.665 ;
      RECT MASK 1 116.564 82.66 127.654 82.7 ;
      RECT MASK 1 2.169 82.75 4.491 82.79 ;
      RECT MASK 1 6.181 82.88 56.9 83.08 ;
      RECT MASK 1 57.174 82.88 64.42 83.08 ;
      RECT MASK 1 64.694 82.88 113.072 83.08 ;
      RECT MASK 1 116.564 82.9 127.654 82.94 ;
      RECT MASK 1 2.169 82.99 4.491 83.03 ;
      RECT MASK 1 116.564 83.14 127.654 83.18 ;
      RECT MASK 1 2.169 83.23 4.491 83.27 ;
      RECT MASK 1 57.178 83.26 64.425 83.32 ;
      RECT MASK 1 116.564 83.38 127.654 83.42 ;
      RECT MASK 1 2.169 83.47 4.491 83.51 ;
      RECT MASK 1 6.616 83.584 7 83.684 ;
      RECT MASK 1 7.778 83.584 8.162 83.684 ;
      RECT MASK 1 8.94 83.584 9.324 83.684 ;
      RECT MASK 1 12.072 83.584 12.456 83.684 ;
      RECT MASK 1 13.234 83.584 13.618 83.684 ;
      RECT MASK 1 14.396 83.584 14.78 83.684 ;
      RECT MASK 1 15.558 83.584 15.942 83.684 ;
      RECT MASK 1 18.69 83.584 19.074 83.684 ;
      RECT MASK 1 19.852 83.584 20.236 83.684 ;
      RECT MASK 1 21.014 83.584 21.398 83.684 ;
      RECT MASK 1 22.176 83.584 22.56 83.684 ;
      RECT MASK 1 25.308 83.584 25.692 83.684 ;
      RECT MASK 1 26.47 83.584 26.854 83.684 ;
      RECT MASK 1 27.632 83.584 28.016 83.684 ;
      RECT MASK 1 28.794 83.584 29.178 83.684 ;
      RECT MASK 1 31.926 83.584 32.31 83.684 ;
      RECT MASK 1 33.088 83.584 33.472 83.684 ;
      RECT MASK 1 34.25 83.584 34.634 83.684 ;
      RECT MASK 1 35.412 83.584 35.796 83.684 ;
      RECT MASK 1 38.544 83.584 38.928 83.684 ;
      RECT MASK 1 39.706 83.584 40.09 83.684 ;
      RECT MASK 1 40.868 83.584 41.252 83.684 ;
      RECT MASK 1 42.03 83.584 42.414 83.684 ;
      RECT MASK 1 45.162 83.584 45.546 83.684 ;
      RECT MASK 1 46.324 83.584 46.708 83.684 ;
      RECT MASK 1 47.486 83.584 47.87 83.684 ;
      RECT MASK 1 48.648 83.584 49.032 83.684 ;
      RECT MASK 1 51.78 83.584 52.164 83.684 ;
      RECT MASK 1 52.942 83.584 53.326 83.684 ;
      RECT MASK 1 54.104 83.584 54.488 83.684 ;
      RECT MASK 1 55.266 83.584 55.65 83.684 ;
      RECT MASK 1 57.178 83.584 58.042 83.684 ;
      RECT MASK 1 58.398 83.584 58.782 83.684 ;
      RECT MASK 1 59.56 83.584 59.944 83.684 ;
      RECT MASK 1 60.722 83.584 61.106 83.684 ;
      RECT MASK 1 61.884 83.584 62.268 83.684 ;
      RECT MASK 1 63.004 83.584 64.425 83.684 ;
      RECT MASK 1 65.016 83.584 65.4 83.684 ;
      RECT MASK 1 66.178 83.584 66.562 83.684 ;
      RECT MASK 1 67.34 83.584 67.724 83.684 ;
      RECT MASK 1 68.502 83.584 68.886 83.684 ;
      RECT MASK 1 71.634 83.584 72.018 83.684 ;
      RECT MASK 1 72.796 83.584 73.18 83.684 ;
      RECT MASK 1 73.958 83.584 74.342 83.684 ;
      RECT MASK 1 75.12 83.584 75.504 83.684 ;
      RECT MASK 1 78.252 83.584 78.636 83.684 ;
      RECT MASK 1 79.414 83.584 79.798 83.684 ;
      RECT MASK 1 80.576 83.584 80.96 83.684 ;
      RECT MASK 1 81.738 83.584 82.122 83.684 ;
      RECT MASK 1 84.87 83.584 85.254 83.684 ;
      RECT MASK 1 86.032 83.584 86.416 83.684 ;
      RECT MASK 1 87.194 83.584 87.578 83.684 ;
      RECT MASK 1 88.356 83.584 88.74 83.684 ;
      RECT MASK 1 91.488 83.584 91.872 83.684 ;
      RECT MASK 1 92.65 83.584 93.034 83.684 ;
      RECT MASK 1 93.812 83.584 94.196 83.684 ;
      RECT MASK 1 94.974 83.584 95.358 83.684 ;
      RECT MASK 1 98.106 83.584 98.49 83.684 ;
      RECT MASK 1 99.268 83.584 99.652 83.684 ;
      RECT MASK 1 100.43 83.584 100.814 83.684 ;
      RECT MASK 1 101.592 83.584 101.976 83.684 ;
      RECT MASK 1 104.724 83.584 105.108 83.684 ;
      RECT MASK 1 105.886 83.584 106.27 83.684 ;
      RECT MASK 1 107.048 83.584 107.432 83.684 ;
      RECT MASK 1 108.21 83.584 108.594 83.684 ;
      RECT MASK 1 116.564 83.62 127.654 83.66 ;
      RECT MASK 1 2.169 83.71 4.491 83.75 ;
      RECT MASK 1 116.564 83.86 127.654 83.9 ;
      RECT MASK 1 2.169 83.95 4.491 83.99 ;
      RECT MASK 1 116.564 84.1 127.654 84.14 ;
      RECT MASK 1 2.169 84.19 4.491 84.23 ;
      RECT MASK 1 6.193 84.258 56.89 84.438 ;
      RECT MASK 1 57.174 84.258 64.42 84.438 ;
      RECT MASK 1 64.694 84.258 113.373 84.438 ;
      RECT MASK 1 116.564 84.34 127.654 84.38 ;
      RECT MASK 1 2.169 84.43 4.491 84.47 ;
      RECT MASK 1 116.564 84.58 127.654 84.62 ;
      RECT MASK 1 2.169 84.67 4.491 84.71 ;
      RECT MASK 1 116.564 84.82 127.654 84.86 ;
      RECT MASK 1 2.169 84.91 4.491 84.95 ;
      RECT MASK 1 116.564 85.06 127.654 85.1 ;
      RECT MASK 1 2.169 85.15 4.491 85.19 ;
      RECT MASK 1 116.564 85.3 127.654 85.34 ;
      RECT MASK 1 2.169 85.39 4.491 85.43 ;
      RECT MASK 1 116.564 85.54 127.654 85.58 ;
      RECT MASK 1 2.169 85.63 4.491 85.67 ;
      RECT MASK 1 24.397 85.686 25.055 85.786 ;
      RECT MASK 1 116.564 85.78 127.654 85.82 ;
      RECT MASK 1 2.169 85.87 4.491 85.91 ;
      RECT MASK 1 116.564 86.02 127.654 86.06 ;
      RECT MASK 1 2.169 86.11 4.491 86.15 ;
      RECT MASK 1 72.062 86.242 72.202 95.438 ;
      RECT MASK 1 103.38 86.242 103.52 95.438 ;
      RECT MASK 1 116.564 86.26 127.654 86.3 ;
      RECT MASK 1 69.863 86.285 71.692 86.485 ;
      RECT MASK 1 103.89 86.285 105.719 86.485 ;
      RECT MASK 1 2.169 86.35 4.491 86.39 ;
      RECT MASK 1 35.672 86.35 35.812 95.33 ;
      RECT MASK 1 66.99 86.35 67.13 95.33 ;
      RECT MASK 1 33.473 86.375 35.302 86.575 ;
      RECT MASK 1 67.491 86.375 69.163 86.575 ;
      RECT MASK 1 26.225 86.43 26.285 92.31 ;
      RECT MASK 1 26.495 86.43 26.555 92.31 ;
      RECT MASK 1 26.765 86.43 26.825 92.31 ;
      RECT MASK 1 27.035 86.43 27.095 92.31 ;
      RECT MASK 1 27.305 86.43 27.365 92.31 ;
      RECT MASK 1 27.575 86.43 27.635 92.31 ;
      RECT MASK 1 27.845 86.43 27.905 92.31 ;
      RECT MASK 1 28.115 86.43 28.175 92.31 ;
      RECT MASK 1 28.385 86.43 28.445 92.31 ;
      RECT MASK 1 28.655 86.43 28.715 92.31 ;
      RECT MASK 1 28.925 86.43 28.985 92.31 ;
      RECT MASK 1 29.195 86.43 29.255 92.31 ;
      RECT MASK 1 29.465 86.43 29.525 92.31 ;
      RECT MASK 1 29.735 86.43 29.795 92.31 ;
      RECT MASK 1 30.005 86.43 30.065 92.31 ;
      RECT MASK 1 36.1535 86.469 66.6485 86.569 ;
      RECT MASK 1 72.5435 86.469 103.0385 86.569 ;
      RECT MASK 1 116.564 86.5 127.654 86.54 ;
      RECT MASK 1 2.169 86.59 4.491 86.63 ;
      RECT MASK 1 70.359 86.735 71.692 86.935 ;
      RECT MASK 1 103.89 86.735 105.223 86.935 ;
      RECT MASK 1 69.797 86.745 69.897 94.935 ;
      RECT MASK 1 105.685 86.745 105.785 94.935 ;
      RECT MASK 1 33.969 86.825 35.302 87.025 ;
      RECT MASK 1 67.494 86.825 68.8145 87.025 ;
      RECT MASK 1 2.169 86.83 4.491 86.87 ;
      RECT MASK 1 33.407 86.835 33.507 94.845 ;
      RECT MASK 1 69.129 86.835 69.229 94.845 ;
      RECT MASK 1 2.169 87.07 4.491 87.11 ;
      RECT MASK 1 14.7225 87.07 23.518 87.17 ;
      RECT MASK 1 25.864 87.096 25.924 88.922 ;
      RECT MASK 1 30.366 87.096 30.426 88.922 ;
      RECT MASK 1 70.129 87.1235 70.229 94.5565 ;
      RECT MASK 1 105.353 87.1235 105.453 94.5565 ;
      RECT MASK 1 36.326 87.147 66.476 87.207 ;
      RECT MASK 1 72.716 87.147 102.866 87.207 ;
      RECT MASK 1 33.739 87.285 33.839 94.395 ;
      RECT MASK 1 34.365 87.285 34.465 94.395 ;
      RECT MASK 1 34.697 87.285 34.797 94.395 ;
      RECT MASK 1 35.029 87.285 35.129 94.395 ;
      RECT MASK 1 67.839 87.285 67.939 94.395 ;
      RECT MASK 1 68.171 87.285 68.271 94.395 ;
      RECT MASK 1 68.797 87.285 68.897 94.395 ;
      RECT MASK 1 70.755 87.3 70.855 94.38 ;
      RECT MASK 1 71.087 87.3 71.187 94.38 ;
      RECT MASK 1 71.419 87.3 71.519 94.38 ;
      RECT MASK 1 104.063 87.3 104.163 94.38 ;
      RECT MASK 1 104.395 87.3 104.495 94.38 ;
      RECT MASK 1 104.727 87.3 104.827 94.38 ;
      RECT MASK 1 2.169 87.31 4.491 87.35 ;
      RECT MASK 1 36.326 87.399 66.476 87.459 ;
      RECT MASK 1 72.716 87.399 102.866 87.459 ;
      RECT MASK 1 9.68 87.52 23.924 87.62 ;
      RECT MASK 1 2.169 87.55 4.491 87.59 ;
      RECT MASK 1 2.169 87.79 4.491 87.83 ;
      RECT MASK 1 2.169 88.03 4.491 88.07 ;
      RECT MASK 1 36.326 88.047 36.778 88.107 ;
      RECT MASK 1 37.048 88.047 65.754 88.107 ;
      RECT MASK 1 66.024 88.047 66.476 88.107 ;
      RECT MASK 1 72.716 88.047 73.168 88.107 ;
      RECT MASK 1 73.438 88.047 102.144 88.107 ;
      RECT MASK 1 102.414 88.047 102.866 88.107 ;
      RECT MASK 1 108.344 88.09 127.654 88.13 ;
      RECT MASK 1 13.784 88.155 16.627 88.335 ;
      RECT MASK 1 2.169 88.27 4.491 88.31 ;
      RECT MASK 1 36.326 88.299 36.778 88.359 ;
      RECT MASK 1 37.048 88.299 65.754 88.359 ;
      RECT MASK 1 66.024 88.299 66.476 88.359 ;
      RECT MASK 1 72.716 88.299 73.168 88.359 ;
      RECT MASK 1 73.438 88.299 102.144 88.359 ;
      RECT MASK 1 102.414 88.299 102.866 88.359 ;
      RECT MASK 1 108.344 88.33 127.654 88.37 ;
      RECT MASK 1 2.169 88.51 4.491 88.55 ;
      RECT MASK 1 108.344 88.57 127.654 88.61 ;
      RECT MASK 1 14.6495 88.74 21.734 88.8 ;
      RECT MASK 1 2.169 88.75 4.491 88.79 ;
      RECT MASK 1 108.344 88.81 127.654 88.85 ;
      RECT MASK 1 5.984 88.812 7.422 88.992 ;
      RECT MASK 1 36.326 88.947 66.476 89.007 ;
      RECT MASK 1 72.716 88.947 102.866 89.007 ;
      RECT MASK 1 2.169 88.99 4.491 89.03 ;
      RECT MASK 1 108.344 89.05 127.654 89.09 ;
      RECT MASK 1 9.6585 89.15 11.3185 89.23 ;
      RECT MASK 1 14.7065 89.15 15.7025 89.23 ;
      RECT MASK 1 19.0905 89.15 20.7505 89.23 ;
      RECT MASK 1 36.326 89.199 66.476 89.259 ;
      RECT MASK 1 72.716 89.199 102.866 89.259 ;
      RECT MASK 1 2.169 89.23 4.491 89.27 ;
      RECT MASK 1 108.344 89.29 127.654 89.33 ;
      RECT MASK 1 25.864 89.436 25.924 91.262 ;
      RECT MASK 1 30.366 89.436 30.426 91.262 ;
      RECT MASK 1 2.169 89.47 4.491 89.51 ;
      RECT MASK 1 14.6495 89.49 21.734 89.55 ;
      RECT MASK 1 108.344 89.53 127.654 89.57 ;
      RECT MASK 1 2.169 89.71 4.491 89.75 ;
      RECT MASK 1 9.503 89.73 20.9155 89.79 ;
      RECT MASK 1 108.344 89.77 127.654 89.81 ;
      RECT MASK 1 36.326 89.847 36.778 89.907 ;
      RECT MASK 1 37.048 89.847 65.754 89.907 ;
      RECT MASK 1 66.024 89.847 66.476 89.907 ;
      RECT MASK 1 72.716 89.847 73.168 89.907 ;
      RECT MASK 1 73.438 89.847 102.144 89.907 ;
      RECT MASK 1 102.414 89.847 102.866 89.907 ;
      RECT MASK 1 2.169 89.95 4.491 89.99 ;
      RECT MASK 1 108.344 90.01 127.654 90.05 ;
      RECT MASK 1 36.326 90.099 36.778 90.159 ;
      RECT MASK 1 37.048 90.099 65.754 90.159 ;
      RECT MASK 1 66.024 90.099 66.476 90.159 ;
      RECT MASK 1 72.716 90.099 73.168 90.159 ;
      RECT MASK 1 73.438 90.099 102.144 90.159 ;
      RECT MASK 1 102.414 90.099 102.866 90.159 ;
      RECT MASK 1 5.984 90.18 7.422 90.36 ;
      RECT MASK 1 2.169 90.19 4.491 90.23 ;
      RECT MASK 1 108.344 90.25 127.654 90.29 ;
      RECT MASK 1 7.617 90.28 22.492 90.38 ;
      RECT MASK 1 2.169 90.43 4.491 90.47 ;
      RECT MASK 1 108.344 90.49 127.654 90.53 ;
      RECT MASK 1 2.169 90.67 4.491 90.71 ;
      RECT MASK 1 6.511 90.73 22.492 90.83 ;
      RECT MASK 1 108.344 90.73 127.654 90.77 ;
      RECT MASK 1 36.326 90.747 66.476 90.807 ;
      RECT MASK 1 72.716 90.747 102.866 90.807 ;
      RECT MASK 1 2.169 90.91 4.491 90.95 ;
      RECT MASK 1 108.344 90.97 127.654 91.01 ;
      RECT MASK 1 36.326 90.999 66.476 91.059 ;
      RECT MASK 1 72.716 90.999 102.866 91.059 ;
      RECT MASK 1 2.169 91.15 4.491 91.19 ;
      RECT MASK 1 7.617 91.18 22.492 91.28 ;
      RECT MASK 1 5.984 91.2 7.422 91.38 ;
      RECT MASK 1 108.344 91.21 127.654 91.25 ;
      RECT MASK 1 2.169 91.39 4.491 91.43 ;
      RECT MASK 1 108.344 91.45 127.654 91.49 ;
      RECT MASK 1 2.169 91.63 4.491 91.67 ;
      RECT MASK 1 36.326 91.647 36.778 91.707 ;
      RECT MASK 1 37.048 91.647 65.754 91.707 ;
      RECT MASK 1 66.024 91.647 66.476 91.707 ;
      RECT MASK 1 72.716 91.647 73.168 91.707 ;
      RECT MASK 1 73.438 91.647 102.144 91.707 ;
      RECT MASK 1 102.414 91.647 102.866 91.707 ;
      RECT MASK 1 108.344 91.69 127.654 91.73 ;
      RECT MASK 1 9.2005 91.765 20.9155 91.825 ;
      RECT MASK 1 2.169 91.87 4.491 91.91 ;
      RECT MASK 1 36.326 91.899 36.778 91.959 ;
      RECT MASK 1 37.048 91.899 65.754 91.959 ;
      RECT MASK 1 66.024 91.899 66.476 91.959 ;
      RECT MASK 1 72.716 91.899 73.168 91.959 ;
      RECT MASK 1 73.438 91.899 102.144 91.959 ;
      RECT MASK 1 102.414 91.899 102.866 91.959 ;
      RECT MASK 1 25.415 91.919 25.475 92.31 ;
      RECT MASK 1 25.685 91.919 25.745 92.31 ;
      RECT MASK 1 25.955 91.919 26.015 92.31 ;
      RECT MASK 1 30.275 91.919 30.335 92.31 ;
      RECT MASK 1 30.545 91.919 30.605 92.31 ;
      RECT MASK 1 30.815 91.919 30.875 92.31 ;
      RECT MASK 1 108.344 91.93 127.654 91.97 ;
      RECT MASK 1 14.6495 92.015 21.734 92.075 ;
      RECT MASK 1 2.169 92.11 4.491 92.15 ;
      RECT MASK 1 108.344 92.17 127.654 92.21 ;
      RECT MASK 1 9.6585 92.33 10.9715 92.41 ;
      RECT MASK 1 14.7065 92.33 15.7025 92.41 ;
      RECT MASK 1 19.0905 92.33 20.7505 92.41 ;
      RECT MASK 1 2.169 92.35 4.491 92.39 ;
      RECT MASK 1 108.344 92.41 127.654 92.45 ;
      RECT MASK 1 36.326 92.547 66.476 92.607 ;
      RECT MASK 1 72.716 92.547 102.866 92.607 ;
      RECT MASK 1 5.984 92.568 7.422 92.748 ;
      RECT MASK 1 2.169 92.59 4.491 92.63 ;
      RECT MASK 1 108.344 92.65 127.654 92.69 ;
      RECT MASK 1 14.6495 92.755 21.734 92.815 ;
      RECT MASK 1 36.326 92.799 66.476 92.859 ;
      RECT MASK 1 72.716 92.799 102.866 92.859 ;
      RECT MASK 1 2.169 92.83 4.491 92.87 ;
      RECT MASK 1 108.344 92.89 127.654 92.93 ;
      RECT MASK 1 2.169 93.07 4.491 93.11 ;
      RECT MASK 1 108.344 93.13 127.654 93.17 ;
      RECT MASK 1 13.4905 93.225 16.956 93.405 ;
      RECT MASK 1 2.169 93.31 4.491 93.35 ;
      RECT MASK 1 108.344 93.37 127.654 93.41 ;
      RECT MASK 1 36.326 93.447 36.778 93.507 ;
      RECT MASK 1 37.048 93.447 65.754 93.507 ;
      RECT MASK 1 66.024 93.447 66.476 93.507 ;
      RECT MASK 1 72.716 93.447 73.168 93.507 ;
      RECT MASK 1 73.438 93.447 102.144 93.507 ;
      RECT MASK 1 102.414 93.447 102.866 93.507 ;
      RECT MASK 1 2.169 93.55 4.491 93.59 ;
      RECT MASK 1 108.344 93.61 127.654 93.65 ;
      RECT MASK 1 36.326 93.699 36.778 93.759 ;
      RECT MASK 1 37.048 93.699 65.754 93.759 ;
      RECT MASK 1 66.024 93.699 66.476 93.759 ;
      RECT MASK 1 72.716 93.699 73.168 93.759 ;
      RECT MASK 1 73.438 93.699 102.144 93.759 ;
      RECT MASK 1 102.414 93.699 102.866 93.759 ;
      RECT MASK 1 2.169 93.79 4.491 93.83 ;
      RECT MASK 1 108.344 93.85 127.654 93.89 ;
      RECT MASK 1 9.68 93.94 24.299 94.04 ;
      RECT MASK 1 2.169 94.03 4.491 94.07 ;
      RECT MASK 1 108.344 94.09 127.654 94.13 ;
      RECT MASK 1 2.169 94.27 4.491 94.31 ;
      RECT MASK 1 108.344 94.33 127.654 94.37 ;
      RECT MASK 1 36.326 94.347 66.476 94.407 ;
      RECT MASK 1 72.716 94.347 102.866 94.407 ;
      RECT MASK 1 14.7225 94.39 24.497 94.49 ;
      RECT MASK 1 2.169 94.51 4.491 94.55 ;
      RECT MASK 1 108.344 94.57 127.654 94.61 ;
      RECT MASK 1 36.326 94.599 66.476 94.659 ;
      RECT MASK 1 72.716 94.599 102.866 94.659 ;
      RECT MASK 1 33.969 94.655 35.302 94.855 ;
      RECT MASK 1 67.52 94.655 68.738 94.855 ;
      RECT MASK 1 70.359 94.745 71.692 94.945 ;
      RECT MASK 1 103.89 94.745 105.223 94.945 ;
      RECT MASK 1 2.169 94.75 4.491 94.79 ;
      RECT MASK 1 108.344 94.81 127.654 94.85 ;
      RECT MASK 1 2.169 94.99 4.491 95.03 ;
      RECT MASK 1 108.344 95.05 127.654 95.09 ;
      RECT MASK 1 33.473 95.105 35.302 95.305 ;
      RECT MASK 1 67.519 95.105 69.163 95.305 ;
      RECT MASK 1 36.1535 95.111 66.6485 95.211 ;
      RECT MASK 1 72.5435 95.111 103.0385 95.211 ;
      RECT MASK 1 69.863 95.195 71.692 95.395 ;
      RECT MASK 1 103.89 95.195 105.719 95.395 ;
      RECT MASK 1 2.169 95.23 4.491 95.27 ;
      RECT MASK 1 108.344 95.29 127.654 95.33 ;
      RECT MASK 1 2.169 95.47 4.491 95.51 ;
      RECT MASK 1 108.344 95.53 127.654 95.57 ;
      RECT MASK 1 2.169 95.71 4.491 95.75 ;
      RECT MASK 1 108.344 95.77 127.654 95.81 ;
      RECT MASK 1 108.344 96.01 127.654 96.05 ;
      RECT MASK 1 108.344 96.25 127.654 96.29 ;
      RECT MASK 1 108.344 96.49 127.654 96.53 ;
      RECT MASK 1 2.303 97.63 43.533 97.67 ;
      RECT MASK 1 45.695 97.63 86.925 97.67 ;
      RECT MASK 1 89.054 97.63 127.544 97.67 ;
      RECT MASK 1 2.303 97.87 43.533 97.91 ;
      RECT MASK 1 45.695 97.87 86.925 97.91 ;
      RECT MASK 1 89.054 97.87 127.544 97.91 ;
      RECT MASK 1 2.303 98.11 43.533 98.15 ;
      RECT MASK 1 45.695 98.11 86.925 98.15 ;
      RECT MASK 1 89.054 98.11 127.544 98.15 ;
      RECT MASK 1 2.303 98.35 43.533 98.39 ;
      RECT MASK 1 45.695 98.35 86.925 98.39 ;
      RECT MASK 1 89.054 98.35 127.544 98.39 ;
      RECT MASK 1 2.303 98.59 43.533 98.63 ;
      RECT MASK 1 45.695 98.59 86.925 98.63 ;
      RECT MASK 1 89.054 98.59 127.544 98.63 ;
      RECT MASK 1 2.303 98.83 43.533 98.87 ;
      RECT MASK 1 45.695 98.83 86.925 98.87 ;
      RECT MASK 1 89.054 98.83 127.544 98.87 ;
      RECT MASK 1 2.303 99.07 43.533 99.11 ;
      RECT MASK 1 45.695 99.07 86.925 99.11 ;
      RECT MASK 1 89.054 99.07 127.544 99.11 ;
      RECT MASK 1 2.303 99.31 43.533 99.35 ;
      RECT MASK 1 45.695 99.31 86.925 99.35 ;
      RECT MASK 1 89.054 99.31 127.544 99.35 ;
      RECT MASK 1 2.303 99.55 43.533 99.59 ;
      RECT MASK 1 45.695 99.55 86.925 99.59 ;
      RECT MASK 1 89.054 99.55 127.544 99.59 ;
      RECT MASK 1 2.303 99.79 43.533 99.83 ;
      RECT MASK 1 45.695 99.79 86.925 99.83 ;
      RECT MASK 1 89.054 99.79 127.544 99.83 ;
      RECT MASK 1 2.303 100.03 43.533 100.07 ;
      RECT MASK 1 45.695 100.03 86.925 100.07 ;
      RECT MASK 1 89.054 100.03 127.544 100.07 ;
      RECT MASK 1 2.303 100.27 43.533 100.31 ;
      RECT MASK 1 45.695 100.27 86.925 100.31 ;
      RECT MASK 1 89.054 100.27 127.544 100.31 ;
      RECT MASK 1 2.303 100.51 43.533 100.55 ;
      RECT MASK 1 45.695 100.51 86.925 100.55 ;
      RECT MASK 1 89.054 100.51 127.544 100.55 ;
      RECT MASK 1 2.303 100.75 43.533 100.79 ;
      RECT MASK 1 45.695 100.75 86.925 100.79 ;
      RECT MASK 1 89.054 100.75 127.544 100.79 ;
      RECT MASK 1 2.303 100.99 43.533 101.03 ;
      RECT MASK 1 45.695 100.99 86.925 101.03 ;
      RECT MASK 1 89.054 100.99 127.544 101.03 ;
      RECT MASK 1 2.303 101.23 43.533 101.27 ;
      RECT MASK 1 45.695 101.23 86.925 101.27 ;
      RECT MASK 1 89.054 101.23 127.544 101.27 ;
      RECT MASK 1 2.303 101.47 43.533 101.51 ;
      RECT MASK 1 45.695 101.47 86.925 101.51 ;
      RECT MASK 1 89.054 101.47 127.544 101.51 ;
      RECT MASK 1 2.303 101.71 43.533 101.75 ;
      RECT MASK 1 45.695 101.71 86.925 101.75 ;
      RECT MASK 1 89.054 101.71 127.544 101.75 ;
      RECT MASK 1 2.303 101.95 43.533 101.99 ;
      RECT MASK 1 45.695 101.95 86.925 101.99 ;
      RECT MASK 1 89.054 101.95 127.544 101.99 ;
      RECT MASK 1 2.303 102.19 43.533 102.23 ;
      RECT MASK 1 45.695 102.19 86.925 102.23 ;
      RECT MASK 1 89.054 102.19 127.544 102.23 ;
      RECT MASK 1 2.303 102.43 43.533 102.47 ;
      RECT MASK 1 45.695 102.43 86.925 102.47 ;
      RECT MASK 1 89.054 102.43 127.544 102.47 ;
      RECT MASK 1 2.303 102.67 43.533 102.71 ;
      RECT MASK 1 45.695 102.67 86.925 102.71 ;
      RECT MASK 1 89.054 102.67 127.544 102.71 ;
      RECT MASK 1 2.303 102.91 43.533 102.95 ;
      RECT MASK 1 45.695 102.91 86.925 102.95 ;
      RECT MASK 1 89.054 102.91 127.544 102.95 ;
      RECT MASK 1 2.303 103.15 43.533 103.19 ;
      RECT MASK 1 45.695 103.15 86.925 103.19 ;
      RECT MASK 1 89.054 103.15 127.544 103.19 ;
      RECT MASK 1 2.303 103.39 43.533 103.43 ;
      RECT MASK 1 45.695 103.39 86.925 103.43 ;
      RECT MASK 1 89.054 103.39 127.544 103.43 ;
      RECT MASK 1 2.303 103.63 43.533 103.67 ;
      RECT MASK 1 45.695 103.63 86.925 103.67 ;
      RECT MASK 1 89.054 103.63 127.544 103.67 ;
      RECT MASK 1 2.303 103.87 43.533 103.91 ;
      RECT MASK 1 45.695 103.87 86.925 103.91 ;
      RECT MASK 1 89.054 103.87 127.544 103.91 ;
      RECT MASK 1 2.303 104.11 43.533 104.15 ;
      RECT MASK 1 45.695 104.11 86.925 104.15 ;
      RECT MASK 1 89.054 104.11 127.544 104.15 ;
      RECT MASK 1 2.303 104.35 43.533 104.39 ;
      RECT MASK 1 45.695 104.35 86.925 104.39 ;
      RECT MASK 1 89.054 104.35 127.544 104.39 ;
      RECT MASK 1 2.303 104.59 43.533 104.63 ;
      RECT MASK 1 45.695 104.59 86.925 104.63 ;
      RECT MASK 1 89.054 104.59 127.544 104.63 ;
      RECT MASK 1 2.303 104.83 43.533 104.87 ;
      RECT MASK 1 45.695 104.83 86.925 104.87 ;
      RECT MASK 1 89.054 104.83 127.544 104.87 ;
      RECT MASK 1 2.303 105.07 43.533 105.11 ;
      RECT MASK 1 45.695 105.07 86.925 105.11 ;
      RECT MASK 1 89.054 105.07 127.544 105.11 ;
      RECT MASK 1 2.303 105.31 43.533 105.35 ;
      RECT MASK 1 45.695 105.31 86.925 105.35 ;
      RECT MASK 1 89.054 105.31 127.544 105.35 ;
      RECT MASK 1 2.303 105.55 43.533 105.59 ;
      RECT MASK 1 45.695 105.55 86.925 105.59 ;
      RECT MASK 1 89.054 105.55 127.544 105.59 ;
      RECT MASK 1 2.303 105.79 43.533 105.83 ;
      RECT MASK 1 45.695 105.79 86.925 105.83 ;
      RECT MASK 1 89.054 105.79 127.544 105.83 ;
      RECT MASK 1 2.303 106.03 43.533 106.07 ;
      RECT MASK 1 45.695 106.03 86.925 106.07 ;
      RECT MASK 1 89.054 106.03 127.544 106.07 ;
      RECT MASK 1 2.303 106.27 43.533 106.31 ;
      RECT MASK 1 45.695 106.27 86.925 106.31 ;
      RECT MASK 1 89.054 106.27 127.544 106.31 ;
      RECT MASK 1 2.303 106.51 43.533 106.55 ;
      RECT MASK 1 45.695 106.51 86.925 106.55 ;
      RECT MASK 1 89.054 106.51 127.544 106.55 ;
      RECT MASK 1 2.303 106.75 43.533 106.79 ;
      RECT MASK 1 45.695 106.75 86.925 106.79 ;
      RECT MASK 1 89.054 106.75 127.544 106.79 ;
      RECT MASK 1 2.303 106.99 43.533 107.03 ;
      RECT MASK 1 45.695 106.99 86.925 107.03 ;
      RECT MASK 1 89.054 106.99 127.544 107.03 ;
      RECT MASK 1 2.303 107.23 43.533 107.27 ;
      RECT MASK 1 45.695 107.23 86.925 107.27 ;
      RECT MASK 1 89.054 107.23 127.544 107.27 ;
      RECT MASK 1 2.303 107.47 43.533 107.51 ;
      RECT MASK 1 45.695 107.47 86.925 107.51 ;
      RECT MASK 1 89.054 107.47 127.544 107.51 ;
    LAYER M3 SPACING 0 ;
      RECT 0 0 130.416 109.44 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 2 23.8135 0.65 48.2385 0.69 ;
      RECT MASK 2 22.8135 0.85 47.6385 0.89 ;
      RECT MASK 2 57.536 0.87 66.237 1.05 ;
      RECT MASK 2 24.2135 1.05 45.9385 1.09 ;
      RECT MASK 2 49.9465 1.13 52.6825 1.17 ;
      RECT MASK 2 23.344 1.25 46.537 1.29 ;
      RECT MASK 2 57.536 1.3 60.453 1.34 ;
      RECT MASK 2 63.778 1.3 66.237 1.34 ;
      RECT MASK 2 49.934 1.33 52.6425 1.37 ;
      RECT MASK 2 61.488 1.54 64.171 1.58 ;
      RECT MASK 2 1.3865 1.8 10.5035 1.98 ;
      RECT MASK 2 11.0835 1.8 12.9405 1.98 ;
      RECT MASK 2 13.6215 1.8 33.3155 1.98 ;
      RECT MASK 2 33.9965 1.8 35.9305 1.98 ;
      RECT MASK 2 36.4335 1.8 45.5505 1.98 ;
      RECT MASK 2 49.3195 1.82 50.2475 1.86 ;
      RECT MASK 2 50.8315 1.82 51.2095 1.86 ;
      RECT MASK 2 51.3895 1.82 51.604 1.86 ;
      RECT MASK 2 52.1595 1.82 52.4375 1.86 ;
      RECT MASK 2 115.3515 1.9 129.1205 1.94 ;
      RECT MASK 2 49.9865 1.98 52.6425 2.02 ;
      RECT MASK 2 61.03 2.02 64.171 2.06 ;
      RECT MASK 2 115.3515 2.14 129.1205 2.18 ;
      RECT MASK 2 1.3865 2.23 21.811 2.27 ;
      RECT MASK 2 22.1665 2.23 24.866 2.31 ;
      RECT MASK 2 25.126 2.23 45.5505 2.27 ;
      RECT MASK 2 58.969 2.26 65.033 2.3 ;
      RECT MASK 2 46.275 2.37 47.156 2.41 ;
      RECT MASK 2 47.5835 2.37 48.4475 2.41 ;
      RECT MASK 2 115.3515 2.38 129.1205 2.42 ;
      RECT MASK 2 2.3125 2.47 9.5875 2.51 ;
      RECT MASK 2 11.0945 2.47 12.9295 2.51 ;
      RECT MASK 2 34.0075 2.47 35.9195 2.51 ;
      RECT MASK 2 37.3495 2.47 44.6245 2.51 ;
      RECT MASK 2 46.6355 2.53 47.4525 2.57 ;
      RECT MASK 2 47.7615 2.53 48.3795 2.57 ;
      RECT MASK 2 115.3515 2.62 129.1205 2.66 ;
      RECT MASK 2 45.873 2.69 49.1005 2.77 ;
      RECT MASK 2 2.3785 2.71 9.6455 2.75 ;
      RECT MASK 2 9.9155 2.71 23.1445 2.75 ;
      RECT MASK 2 23.7925 2.71 37.0215 2.75 ;
      RECT MASK 2 37.2915 2.71 44.5585 2.75 ;
      RECT MASK 2 58.74 2.74 59.308 2.78 ;
      RECT MASK 2 59.656 2.74 60.224 2.78 ;
      RECT MASK 2 63.683 2.74 63.888 2.78 ;
      RECT MASK 2 64.061 2.74 64.804 2.78 ;
      RECT MASK 2 115.3515 2.86 129.1205 2.9 ;
      RECT MASK 2 22.0175 2.87 24.8685 2.95 ;
      RECT MASK 2 8.4845 2.95 13.1245 2.99 ;
      RECT MASK 2 33.8125 2.95 38.4525 2.99 ;
      RECT MASK 2 38.9675 2.95 45.5505 2.99 ;
      RECT MASK 2 45.697 2.95 47.0605 2.99 ;
      RECT MASK 2 47.4305 2.95 48.0485 2.99 ;
      RECT MASK 2 49.9515 2.97 52.6775 3.03 ;
      RECT MASK 2 58.769 2.98 64.801 3.02 ;
      RECT MASK 2 115.3515 3.1 129.1205 3.14 ;
      RECT MASK 2 45.763 3.11 47.2105 3.15 ;
      RECT MASK 2 8.7135 3.19 12.6385 3.23 ;
      RECT MASK 2 12.9125 3.19 21.3145 3.23 ;
      RECT MASK 2 22.0175 3.19 24.8685 3.27 ;
      RECT MASK 2 25.6225 3.19 34.0245 3.23 ;
      RECT MASK 2 34.2985 3.19 38.2235 3.23 ;
      RECT MASK 2 38.9675 3.19 45.5505 3.23 ;
      RECT MASK 2 59.147 3.22 63.659 3.26 ;
      RECT MASK 2 64.007 3.22 64.575 3.26 ;
      RECT MASK 2 47.9205 3.27 48.238 3.31 ;
      RECT MASK 2 115.3515 3.34 129.1205 3.38 ;
      RECT MASK 2 49.9515 3.45 52.6775 3.51 ;
      RECT MASK 2 65.152 3.46 66.8525 3.5 ;
      RECT MASK 2 115.3515 3.58 129.1205 3.62 ;
      RECT MASK 2 49.9515 3.69 52.6775 3.75 ;
      RECT MASK 2 57.536 3.7 60.453 3.74 ;
      RECT MASK 2 61.304 3.7 66.237 3.74 ;
      RECT MASK 2 115.3515 3.82 129.1205 3.86 ;
      RECT MASK 2 46.643 3.91 47.033 3.95 ;
      RECT MASK 2 47.243 3.91 47.664 3.95 ;
      RECT MASK 2 49.9515 3.93 52.6775 3.99 ;
      RECT MASK 2 57.536 3.98 60.453 4.18 ;
      RECT MASK 2 61.304 3.99 66.237 4.17 ;
      RECT MASK 2 115.3515 4.06 129.1205 4.1 ;
      RECT MASK 2 22.0175 4.11 24.8685 4.19 ;
      RECT MASK 2 45.9535 4.13 49.1005 4.21 ;
      RECT MASK 2 8.7135 4.15 12.6385 4.19 ;
      RECT MASK 2 12.9125 4.15 21.3145 4.19 ;
      RECT MASK 2 25.6225 4.15 34.0245 4.19 ;
      RECT MASK 2 34.2985 4.15 38.2235 4.19 ;
      RECT MASK 2 38.9675 4.15 45.5505 4.19 ;
      RECT MASK 2 115.3515 4.3 129.1205 4.34 ;
      RECT MASK 2 8.4845 4.39 13.1245 4.43 ;
      RECT MASK 2 33.8125 4.39 38.4525 4.43 ;
      RECT MASK 2 38.9675 4.39 45.5505 4.43 ;
      RECT MASK 2 72.7145 4.405 113.9905 4.655 ;
      RECT MASK 2 57.536 4.42 60.453 4.46 ;
      RECT MASK 2 61.304 4.42 66.237 4.46 ;
      RECT MASK 2 22.0175 4.43 24.8685 4.51 ;
      RECT MASK 2 115.3515 4.54 129.1205 4.58 ;
      RECT MASK 2 2.3785 4.63 9.6455 4.67 ;
      RECT MASK 2 9.9155 4.63 23.1445 4.67 ;
      RECT MASK 2 23.7925 4.63 37.0215 4.67 ;
      RECT MASK 2 37.2915 4.63 44.5585 4.67 ;
      RECT MASK 2 49.9515 4.65 52.6775 4.71 ;
      RECT MASK 2 56.7835 4.66 65.72 4.7 ;
      RECT MASK 2 115.3515 4.78 129.1205 4.82 ;
      RECT MASK 2 2.3125 4.87 9.5875 4.91 ;
      RECT MASK 2 11.0945 4.87 12.9295 4.91 ;
      RECT MASK 2 34.0075 4.87 35.9195 4.91 ;
      RECT MASK 2 37.3495 4.87 44.6245 4.91 ;
      RECT MASK 2 49.9515 4.89 52.6775 4.95 ;
      RECT MASK 2 59.147 4.9 63.659 4.94 ;
      RECT MASK 2 64.007 4.9 64.575 4.94 ;
      RECT MASK 2 115.3515 5.02 129.1205 5.06 ;
      RECT MASK 2 22.1155 5.07 24.866 5.15 ;
      RECT MASK 2 1.3865 5.11 21.811 5.15 ;
      RECT MASK 2 25.126 5.11 45.5505 5.15 ;
      RECT MASK 2 74.7205 5.125 86.5 5.375 ;
      RECT MASK 2 100.205 5.125 111.9845 5.375 ;
      RECT MASK 2 49.9515 5.13 52.6775 5.19 ;
      RECT MASK 2 58.769 5.14 64.801 5.18 ;
      RECT MASK 2 115.3515 5.26 129.1205 5.3 ;
      RECT MASK 2 58.74 5.38 59.308 5.42 ;
      RECT MASK 2 59.656 5.38 60.224 5.42 ;
      RECT MASK 2 63.683 5.38 63.888 5.42 ;
      RECT MASK 2 64.061 5.38 64.804 5.42 ;
      RECT MASK 2 62.5005 5.3975 63.268 5.4575 ;
      RECT MASK 2 1.3865 5.4 10.5035 5.58 ;
      RECT MASK 2 11.0835 5.4 12.9405 5.58 ;
      RECT MASK 2 13.6215 5.4 33.3155 5.58 ;
      RECT MASK 2 33.9965 5.4 35.9305 5.58 ;
      RECT MASK 2 36.4335 5.4 45.5505 5.58 ;
      RECT MASK 2 115.3515 5.5 129.1205 5.54 ;
      RECT MASK 2 46.09 5.592 49.0705 5.772 ;
      RECT MASK 2 53.499 5.712 56.3975 5.892 ;
      RECT MASK 2 115.3515 5.74 129.1205 5.78 ;
      RECT MASK 2 72.7145 5.845 113.9905 6.095 ;
      RECT MASK 2 58.969 5.86 65.033 5.9 ;
      RECT MASK 2 1.3865 5.88 10.5035 6.06 ;
      RECT MASK 2 11.0835 5.88 12.9405 6.06 ;
      RECT MASK 2 13.6215 5.88 33.3155 6.06 ;
      RECT MASK 2 33.9965 5.88 35.9305 6.06 ;
      RECT MASK 2 36.4335 5.88 45.5505 6.06 ;
      RECT MASK 2 115.3515 5.98 129.1205 6.02 ;
      RECT MASK 2 61.03 6.1 64.171 6.14 ;
      RECT MASK 2 47.2725 6.124 56.4965 6.164 ;
      RECT MASK 2 115.3515 6.22 129.1205 6.26 ;
      RECT MASK 2 49.9865 6.284 52.6745 6.344 ;
      RECT MASK 2 1.3865 6.31 21.811 6.35 ;
      RECT MASK 2 22.1155 6.31 24.866 6.39 ;
      RECT MASK 2 25.126 6.31 45.5505 6.35 ;
      RECT MASK 2 53.054 6.316 55.5915 6.356 ;
      RECT MASK 2 115.3515 6.46 129.1205 6.5 ;
      RECT MASK 2 84.7605 6.5 89.677 6.64 ;
      RECT MASK 2 97.028 6.5 101.9445 6.64 ;
      RECT MASK 2 55.3155 6.518 56.1635 6.558 ;
      RECT MASK 2 2.3125 6.55 9.5875 6.59 ;
      RECT MASK 2 11.0945 6.55 12.9295 6.59 ;
      RECT MASK 2 22.6135 6.55 23.426 6.59 ;
      RECT MASK 2 34.0075 6.55 35.9195 6.59 ;
      RECT MASK 2 37.3495 6.55 44.6245 6.59 ;
      RECT MASK 2 23.7135 6.57 24.3235 6.61 ;
      RECT MASK 2 61.488 6.58 64.171 6.62 ;
      RECT MASK 2 115.3515 6.7 129.1205 6.74 ;
      RECT MASK 2 2.3785 6.79 9.6455 6.83 ;
      RECT MASK 2 9.9155 6.79 23.1445 6.83 ;
      RECT MASK 2 23.7925 6.79 37.0215 6.83 ;
      RECT MASK 2 37.2915 6.79 44.5585 6.83 ;
      RECT MASK 2 49.9515 6.81 52.6775 6.87 ;
      RECT MASK 2 57.536 6.82 60.453 6.86 ;
      RECT MASK 2 63.778 6.82 66.237 6.86 ;
      RECT MASK 2 115.3515 6.94 129.1205 6.98 ;
      RECT MASK 2 22.0175 6.95 24.8685 7.03 ;
      RECT MASK 2 8.4845 7.03 13.1245 7.07 ;
      RECT MASK 2 33.8125 7.03 38.4525 7.07 ;
      RECT MASK 2 57.536 7.11 66.237 7.29 ;
      RECT MASK 2 115.3515 7.18 129.1205 7.22 ;
      RECT MASK 2 54.1575 7.2485 56.96 7.2885 ;
      RECT MASK 2 8.7135 7.27 12.6385 7.31 ;
      RECT MASK 2 12.9125 7.27 21.3145 7.31 ;
      RECT MASK 2 22.0175 7.27 24.8685 7.35 ;
      RECT MASK 2 25.6225 7.27 34.0245 7.31 ;
      RECT MASK 2 34.2985 7.27 38.2235 7.31 ;
      RECT MASK 2 74.7435 7.285 88.0615 7.535 ;
      RECT MASK 2 98.6435 7.285 111.9615 7.535 ;
      RECT MASK 2 49.9515 7.29 52.6775 7.35 ;
      RECT MASK 2 47.6045 7.3445 49.4295 7.3845 ;
      RECT MASK 2 115.3515 7.42 129.1205 7.46 ;
      RECT MASK 2 57.536 7.54 60.453 7.58 ;
      RECT MASK 2 63.778 7.54 66.237 7.58 ;
      RECT MASK 2 46.677 7.559 47.464 7.599 ;
      RECT MASK 2 47.7705 7.559 48.0795 7.599 ;
      RECT MASK 2 115.3515 7.66 129.1205 7.7 ;
      RECT MASK 2 46.9405 7.766 49.4295 7.806 ;
      RECT MASK 2 49.9515 7.77 52.6775 7.83 ;
      RECT MASK 2 61.488 7.78 64.171 7.82 ;
      RECT MASK 2 115.3515 7.9 129.1205 7.94 ;
      RECT MASK 2 79.3245 8.005 91.804 8.2625 ;
      RECT MASK 2 94.901 8.005 107.3805 8.255 ;
      RECT MASK 2 66.513 8.0605 71.2185 8.1005 ;
      RECT MASK 2 46.09 8.088 49.0705 8.268 ;
      RECT MASK 2 115.3515 8.14 129.1205 8.18 ;
      RECT MASK 2 49.9515 8.25 52.6775 8.31 ;
      RECT MASK 2 61.03 8.26 64.171 8.3 ;
      RECT MASK 2 35.4365 8.329 42.2685 8.369 ;
      RECT MASK 2 115.3515 8.38 129.1205 8.42 ;
      RECT MASK 2 46.09 8.472 49.0705 8.652 ;
      RECT MASK 2 58.969 8.5 65.033 8.54 ;
      RECT MASK 2 50.2785 8.53 53.33 8.57 ;
      RECT MASK 2 22.0175 8.61 23.485 8.69 ;
      RECT MASK 2 115.3515 8.62 129.1205 8.66 ;
      RECT MASK 2 8.7135 8.65 12.6385 8.69 ;
      RECT MASK 2 12.9125 8.65 21.3145 8.69 ;
      RECT MASK 2 49.6515 8.69 52.475 8.73 ;
      RECT MASK 2 115.3515 8.86 129.1205 8.9 ;
      RECT MASK 2 8.4845 8.89 13.1245 8.93 ;
      RECT MASK 2 44.048 8.9295 47.949 8.9695 ;
      RECT MASK 2 48.209 8.9295 49.5715 8.9695 ;
      RECT MASK 2 22.0175 8.93 23.485 9.01 ;
      RECT MASK 2 67.346 8.952 71.009 9.132 ;
      RECT MASK 2 58.74 8.98 59.308 9.02 ;
      RECT MASK 2 59.656 8.98 60.224 9.02 ;
      RECT MASK 2 63.683 8.98 63.888 9.02 ;
      RECT MASK 2 64.061 8.98 64.804 9.02 ;
      RECT MASK 2 31.3665 8.982 39.3815 9.162 ;
      RECT MASK 2 53.499 8.982 56.4545 9.162 ;
      RECT MASK 2 115.3515 9.1 129.1205 9.14 ;
      RECT MASK 2 46.9405 9.1215 49.2635 9.1615 ;
      RECT MASK 2 2.3785 9.13 9.6455 9.17 ;
      RECT MASK 2 9.9155 9.13 23.1445 9.17 ;
      RECT MASK 2 50.3835 9.13 53.164 9.17 ;
      RECT MASK 2 105.694 9.202 106.578 9.439 ;
      RECT MASK 2 58.769 9.22 64.801 9.26 ;
      RECT MASK 2 49.9515 9.33 52.6775 9.39 ;
      RECT MASK 2 115.3515 9.34 129.1205 9.38 ;
      RECT MASK 2 21.9785 9.3415 22.319 9.3815 ;
      RECT MASK 2 32.8 9.342 43.3825 9.382 ;
      RECT MASK 2 2.3125 9.37 9.5875 9.41 ;
      RECT MASK 2 11.0945 9.37 12.9295 9.41 ;
      RECT MASK 2 47.2725 9.4095 49.7615 9.4495 ;
      RECT MASK 2 59.147 9.46 63.659 9.5 ;
      RECT MASK 2 64.007 9.46 64.575 9.5 ;
      RECT MASK 2 31.2025 9.514 33.597 9.554 ;
      RECT MASK 2 35.09 9.544 43.2065 9.584 ;
      RECT MASK 2 22.1155 9.57 23.4685 9.65 ;
      RECT MASK 2 115.3515 9.58 129.1205 9.62 ;
      RECT MASK 2 69.824 9.603 95.7725 9.643 ;
      RECT MASK 2 1.3865 9.61 21.811 9.65 ;
      RECT MASK 2 68.528 9.612 69.678 9.652 ;
      RECT MASK 2 65.152 9.7 66.1985 9.74 ;
      RECT MASK 2 30.881 9.716 35.429 9.756 ;
      RECT MASK 2 35.8005 9.716 36.3755 9.756 ;
      RECT MASK 2 37.838 9.717 42.8745 9.757 ;
      RECT MASK 2 115.3515 9.82 129.1205 9.86 ;
      RECT MASK 2 46.667 9.828 56.6305 9.868 ;
      RECT MASK 2 66.667 9.891 69.1475 9.931 ;
      RECT MASK 2 1.3865 9.9 10.5035 10.08 ;
      RECT MASK 2 11.0835 9.9 12.9405 10.08 ;
      RECT MASK 2 13.6215 9.9 23.4685 10.08 ;
      RECT MASK 2 27.187 9.918 32.452 9.958 ;
      RECT MASK 2 34.174 9.918 38.917 9.958 ;
      RECT MASK 2 57.536 9.94 60.453 9.98 ;
      RECT MASK 2 61.658 9.94 66.237 9.98 ;
      RECT MASK 2 49.9515 10.05 52.6775 10.11 ;
      RECT MASK 2 115.3515 10.06 129.1205 10.1 ;
      RECT MASK 2 57.536 10.22 60.453 10.42 ;
      RECT MASK 2 61.304 10.23 66.237 10.41 ;
      RECT MASK 2 23.819 10.298 44.158 10.338 ;
      RECT MASK 2 49.6515 10.298 57.351 10.338 ;
      RECT MASK 2 115.3515 10.3 129.1205 10.34 ;
      RECT MASK 2 5.08 10.506 31.189 10.546 ;
      RECT MASK 2 115.3515 10.54 129.1205 10.58 ;
      RECT MASK 2 49.9515 10.65 52.6775 10.71 ;
      RECT MASK 2 31.87 10.694 44.536 10.734 ;
      RECT MASK 2 4.334 10.708 31.5105 10.748 ;
      RECT MASK 2 115.3515 10.78 129.1205 10.82 ;
      RECT MASK 2 43.0965 10.886 62.323 10.926 ;
      RECT MASK 2 24.1425 11.06 32.0675 11.1 ;
      RECT MASK 2 42.7645 11.078 55.517 11.118 ;
      RECT MASK 2 56.4685 11.078 127.473 11.118 ;
      RECT MASK 2 23.037 11.27 89.713 11.31 ;
      RECT MASK 2 115.3515 11.314 129.1205 11.354 ;
      RECT MASK 2 28.847 11.462 83.903 11.502 ;
      RECT MASK 2 115.3515 11.5 129.1205 11.54 ;
      RECT MASK 2 8.927 11.654 103.823 11.694 ;
      RECT MASK 2 115.3515 11.74 129.1205 11.78 ;
      RECT MASK 2 115.3515 11.98 129.1205 12.02 ;
      RECT MASK 2 56.496 12.056 71.057 12.136 ;
      RECT MASK 2 115.3515 12.22 129.1205 12.26 ;
      RECT MASK 2 115.3515 12.46 129.1205 12.5 ;
      RECT MASK 2 25.693 12.484 73.445 12.524 ;
      RECT MASK 2 24.199 12.58 25.305 12.62 ;
      RECT MASK 2 22.539 12.676 23.645 12.716 ;
      RECT MASK 2 37.313 12.676 38.751 12.716 ;
      RECT MASK 2 38.973 12.676 40.411 12.716 ;
      RECT MASK 2 40.799 12.676 41.075 12.716 ;
      RECT MASK 2 41.516 12.676 41.739 12.716 ;
      RECT MASK 2 42.277 12.676 43.731 12.716 ;
      RECT MASK 2 48.767 12.676 60.663 12.716 ;
      RECT MASK 2 60.885 12.676 65.975 12.716 ;
      RECT MASK 2 66.529 12.676 102.827 12.716 ;
      RECT MASK 2 115.3515 12.7 129.1205 12.74 ;
      RECT MASK 2 25.859 12.864 27.463 12.904 ;
      RECT MASK 2 8.595 12.868 9.369 12.908 ;
      RECT MASK 2 10.255 12.868 11.029 12.908 ;
      RECT MASK 2 32.499 12.868 38.585 12.908 ;
      RECT MASK 2 39.139 12.868 43.565 12.908 ;
      RECT MASK 2 44.451 12.868 53.384 12.908 ;
      RECT MASK 2 54.079 12.868 59.833 12.908 ;
      RECT MASK 2 60.221 12.868 71.287 12.908 ;
      RECT MASK 2 115.3515 12.94 129.1205 12.98 ;
      RECT MASK 2 52.419 13.056 59.335 13.096 ;
      RECT MASK 2 24.033 13.058 25.471 13.098 ;
      RECT MASK 2 26.191 13.058 30.285 13.098 ;
      RECT MASK 2 30.839 13.058 31.945 13.098 ;
      RECT MASK 2 32.831 13.058 33.937 13.098 ;
      RECT MASK 2 34.325 13.058 35.597 13.098 ;
      RECT MASK 2 35.819 13.058 36.925 13.098 ;
      RECT MASK 2 37.811 13.058 40.743 13.098 ;
      RECT MASK 2 40.965 13.058 43.233 13.098 ;
      RECT MASK 2 44.119 13.058 45.5575 13.098 ;
      RECT MASK 2 45.945 13.058 47.266 13.098 ;
      RECT MASK 2 47.439 13.058 48.925 13.098 ;
      RECT MASK 2 49.099 13.058 50.57 13.098 ;
      RECT MASK 2 50.759 13.058 51.865 13.098 ;
      RECT MASK 2 59.723 13.058 62.533 13.098 ;
      RECT MASK 2 63.043 13.058 64.315 13.098 ;
      RECT MASK 2 64.669 13.058 70.83 13.098 ;
      RECT MASK 2 72.007 13.058 73.113 13.098 ;
      RECT MASK 2 73.335 13.058 104.487 13.098 ;
      RECT MASK 2 115.3515 13.18 129.1205 13.22 ;
      RECT MASK 2 4.251 13.278 111.819 13.458 ;
      RECT MASK 2 115.3515 13.42 129.1205 13.46 ;
      RECT MASK 2 115.3515 13.66 129.1205 13.7 ;
      RECT MASK 2 115.3515 13.9 129.1205 13.94 ;
      RECT MASK 2 115.3515 14.14 129.1205 14.18 ;
      RECT MASK 2 4.251 14.142 111.819 14.322 ;
      RECT MASK 2 115.3515 14.38 129.1205 14.42 ;
      RECT MASK 2 26.357 14.502 31.447 14.542 ;
      RECT MASK 2 33.827 14.502 42.237 14.542 ;
      RECT MASK 2 43.123 14.502 56.181 14.542 ;
      RECT MASK 2 56.569 14.502 69.627 14.542 ;
      RECT MASK 2 115.3515 14.62 129.1205 14.66 ;
      RECT MASK 2 6.935 14.692 108.054 14.732 ;
      RECT MASK 2 109.689 14.788 111.127 14.828 ;
      RECT MASK 2 115.3515 14.86 129.1205 14.9 ;
      RECT MASK 2 60.553 14.88 63.153 14.92 ;
      RECT MASK 2 4.943 14.884 16.341 14.924 ;
      RECT MASK 2 16.552 14.884 29.621 14.924 ;
      RECT MASK 2 29.843 14.884 42.901 14.924 ;
      RECT MASK 2 49.597 14.884 59.003 14.924 ;
      RECT MASK 2 66.363 14.884 68.133 14.924 ;
      RECT MASK 2 69.849 14.884 82.907 14.924 ;
      RECT MASK 2 83.129 14.884 96.187 14.924 ;
      RECT MASK 2 96.409 14.884 109.467 14.924 ;
      RECT MASK 2 5.441 15.07 6.746 15.11 ;
      RECT MASK 2 7.101 15.07 7.908 15.11 ;
      RECT MASK 2 8.761 15.07 9.203 15.11 ;
      RECT MASK 2 10.421 15.07 11.832 15.11 ;
      RECT MASK 2 12.081 15.07 13.365 15.11 ;
      RECT MASK 2 13.741 15.07 14.526 15.11 ;
      RECT MASK 2 15.401 15.07 15.843 15.11 ;
      RECT MASK 2 17.061 15.07 18.387 15.11 ;
      RECT MASK 2 18.721 15.07 19.982 15.11 ;
      RECT MASK 2 20.381 15.07 21.144 15.11 ;
      RECT MASK 2 22.041 15.07 22.483 15.11 ;
      RECT MASK 2 23.526 15.07 24.67 15.11 ;
      RECT MASK 2 25.361 15.07 26.6 15.11 ;
      RECT MASK 2 27.021 15.07 27.762 15.11 ;
      RECT MASK 2 28.681 15.07 29.123 15.11 ;
      RECT MASK 2 30.341 15.07 31.447 15.11 ;
      RECT MASK 2 32.001 15.07 33.218 15.11 ;
      RECT MASK 2 33.661 15.07 34.38 15.11 ;
      RECT MASK 2 35.321 15.07 35.763 15.11 ;
      RECT MASK 2 36.981 15.07 37.676 15.11 ;
      RECT MASK 2 38.641 15.07 39.836 15.11 ;
      RECT MASK 2 40.301 15.07 40.998 15.11 ;
      RECT MASK 2 41.961 15.07 42.403 15.11 ;
      RECT MASK 2 43.621 15.07 44.276 15.11 ;
      RECT MASK 2 45.281 15.07 46.454 15.11 ;
      RECT MASK 2 46.941 15.07 47.616 15.11 ;
      RECT MASK 2 48.601 15.07 49.043 15.11 ;
      RECT MASK 2 50.261 15.07 51.114 15.11 ;
      RECT MASK 2 51.921 15.07 52.363 15.11 ;
      RECT MASK 2 53.581 15.07 54.234 15.11 ;
      RECT MASK 2 55.241 15.07 55.683 15.11 ;
      RECT MASK 2 57.067 15.07 58.173 15.11 ;
      RECT MASK 2 58.727 15.07 59.69 15.11 ;
      RECT MASK 2 60.387 15.07 60.852 15.11 ;
      RECT MASK 2 61.886 15.07 62.489 15.11 ;
      RECT MASK 2 63.707 15.07 64.424 15.11 ;
      RECT MASK 2 65.367 15.07 66.474 15.11 ;
      RECT MASK 2 67.027 15.07 67.636 15.11 ;
      RECT MASK 2 68.522 15.07 69.129 15.11 ;
      RECT MASK 2 70.347 15.07 71.453 15.11 ;
      RECT MASK 2 72.007 15.07 72.926 15.11 ;
      RECT MASK 2 73.667 15.07 74.254 15.11 ;
      RECT MASK 2 75.14 15.07 75.769 15.11 ;
      RECT MASK 2 76.987 15.07 78.124 15.11 ;
      RECT MASK 2 78.647 15.07 79.655 15.11 ;
      RECT MASK 2 80.307 15.07 80.749 15.11 ;
      RECT MASK 2 81.758 15.07 82.409 15.11 ;
      RECT MASK 2 83.627 15.07 84.162 15.11 ;
      RECT MASK 2 85.287 15.07 86.162 15.11 ;
      RECT MASK 2 86.947 15.07 87.389 15.11 ;
      RECT MASK 2 88.376 15.07 89.049 15.11 ;
      RECT MASK 2 90.267 15.07 91.0055 15.11 ;
      RECT MASK 2 91.927 15.07 92.78 15.11 ;
      RECT MASK 2 93.587 15.07 94.029 15.11 ;
      RECT MASK 2 94.994 15.07 95.689 15.11 ;
      RECT MASK 2 96.907 15.07 97.698 15.11 ;
      RECT MASK 2 98.567 15.07 99.398 15.11 ;
      RECT MASK 2 100.227 15.07 100.669 15.11 ;
      RECT MASK 2 101.612 15.07 102.329 15.11 ;
      RECT MASK 2 103.547 15.07 104.214 15.11 ;
      RECT MASK 2 105.207 15.07 106.016 15.11 ;
      RECT MASK 2 106.867 15.07 107.333 15.11 ;
      RECT MASK 2 108.23 15.07 108.969 15.11 ;
      RECT MASK 2 110.187 15.07 110.629 15.11 ;
      RECT MASK 2 115.3515 15.1 129.1205 15.14 ;
      RECT MASK 2 115.3515 15.34 129.1205 15.38 ;
      RECT MASK 2 56.407 15.56 61.4555 15.88 ;
      RECT MASK 2 115.3515 15.58 129.1205 15.62 ;
      RECT MASK 2 115.3515 15.82 129.1205 15.86 ;
      RECT MASK 2 115.3515 16.06 129.1205 16.1 ;
      RECT MASK 2 115.3515 16.3 129.1205 16.34 ;
      RECT MASK 2 29.677 16.318 32.277 16.358 ;
      RECT MASK 2 53.274 16.318 60.39 16.358 ;
      RECT MASK 2 42.957 16.324 45.557 16.364 ;
      RECT MASK 2 10.255 16.516 105.483 16.556 ;
      RECT MASK 2 115.3515 16.54 129.1205 16.58 ;
      RECT MASK 2 6.603 16.708 13.353 16.748 ;
      RECT MASK 2 13.552 16.708 14.423 16.748 ;
      RECT MASK 2 14.571 16.708 15.013 16.748 ;
      RECT MASK 2 15.235 16.708 16.009 16.748 ;
      RECT MASK 2 16.231 16.708 16.673 16.748 ;
      RECT MASK 2 16.895 16.708 17.669 16.748 ;
      RECT MASK 2 17.891 16.708 18.333 16.748 ;
      RECT MASK 2 18.887 16.708 19.661 16.748 ;
      RECT MASK 2 19.883 16.708 26.6885 16.748 ;
      RECT MASK 2 26.855 16.708 27.629 16.748 ;
      RECT MASK 2 27.851 16.708 28.293 16.748 ;
      RECT MASK 2 28.515 16.708 29.289 16.748 ;
      RECT MASK 2 29.511 16.708 29.953 16.748 ;
      RECT MASK 2 30.175 16.708 30.949 16.748 ;
      RECT MASK 2 31.171 16.708 32.941 16.748 ;
      RECT MASK 2 33.1035 16.708 39.962 16.748 ;
      RECT MASK 2 40.135 16.708 40.909 16.748 ;
      RECT MASK 2 41.131 16.708 41.573 16.748 ;
      RECT MASK 2 41.795 16.708 42.569 16.748 ;
      RECT MASK 2 42.791 16.708 43.233 16.748 ;
      RECT MASK 2 43.455 16.708 44.229 16.748 ;
      RECT MASK 2 44.451 16.708 46.221 16.748 ;
      RECT MASK 2 46.443 16.708 51.201 16.748 ;
      RECT MASK 2 51.423 16.708 52.861 16.748 ;
      RECT MASK 2 53.0475 16.708 53.229 16.748 ;
      RECT MASK 2 53.415 16.708 54.189 16.748 ;
      RECT MASK 2 54.411 16.708 54.853 16.748 ;
      RECT MASK 2 55.074 16.708 55.849 16.748 ;
      RECT MASK 2 56.071 16.708 56.679 16.748 ;
      RECT MASK 2 56.901 16.708 57.675 16.748 ;
      RECT MASK 2 57.897 16.708 59.667 16.748 ;
      RECT MASK 2 59.853 16.708 66.6895 16.748 ;
      RECT MASK 2 66.861 16.708 67.635 16.748 ;
      RECT MASK 2 67.857 16.708 68.299 16.748 ;
      RECT MASK 2 68.521 16.708 69.295 16.748 ;
      RECT MASK 2 69.517 16.708 69.959 16.748 ;
      RECT MASK 2 70.151 16.708 70.97 16.748 ;
      RECT MASK 2 71.177 16.708 72.977 16.748 ;
      RECT MASK 2 73.169 16.708 79.919 16.748 ;
      RECT MASK 2 80.141 16.708 80.915 16.748 ;
      RECT MASK 2 81.087 16.708 81.312 16.748 ;
      RECT MASK 2 81.4545 16.708 82.907 16.748 ;
      RECT MASK 2 83.0435 16.708 83.2795 16.748 ;
      RECT MASK 2 83.461 16.708 84.235 16.748 ;
      RECT MASK 2 84.457 16.708 86.227 16.748 ;
      RECT MASK 2 86.449 16.708 93.199 16.748 ;
      RECT MASK 2 93.421 16.708 94.195 16.748 ;
      RECT MASK 2 94.417 16.708 94.859 16.748 ;
      RECT MASK 2 95.081 16.708 95.898 16.748 ;
      RECT MASK 2 96.077 16.708 96.519 16.748 ;
      RECT MASK 2 96.741 16.708 97.515 16.748 ;
      RECT MASK 2 97.737 16.708 99.507 16.748 ;
      RECT MASK 2 99.729 16.708 106.495 16.748 ;
      RECT MASK 2 106.701 16.708 107.475 16.748 ;
      RECT MASK 2 107.944 16.708 109.135 16.748 ;
      RECT MASK 2 109.523 16.708 110.795 16.748 ;
      RECT MASK 2 115.3515 16.78 129.1205 16.82 ;
      RECT MASK 2 5.275 16.898 110.463 16.938 ;
      RECT MASK 2 115.3515 17.02 129.1205 17.06 ;
      RECT MASK 2 4.251 17.118 111.819 17.298 ;
      RECT MASK 2 115.3515 17.26 129.1205 17.3 ;
      RECT MASK 2 80.31 17.478 81.084 17.518 ;
      RECT MASK 2 115.3515 17.5 129.1205 17.54 ;
      RECT MASK 2 65.168 17.55 67.728 17.73 ;
      RECT MASK 2 115.3515 17.74 129.1205 17.78 ;
      RECT MASK 2 115.3515 17.98 129.1205 18.02 ;
      RECT MASK 2 115.3515 18.22 129.1205 18.26 ;
      RECT MASK 2 5.031 18.45 109.945 18.63 ;
      RECT MASK 2 115.3515 18.46 129.1205 18.5 ;
      RECT MASK 2 115.3515 18.7 129.1205 18.74 ;
      RECT MASK 2 115.3515 18.94 129.1205 18.98 ;
      RECT MASK 2 115.3515 19.18 129.1205 19.22 ;
      RECT MASK 2 115.3515 19.42 129.1205 19.46 ;
      RECT MASK 2 115.3515 19.66 129.1205 19.7 ;
      RECT MASK 2 1.3325 19.78 4.745 19.82 ;
      RECT MASK 2 5.031 19.818 109.945 20.018 ;
      RECT MASK 2 115.3515 19.9 129.1205 19.94 ;
      RECT MASK 2 1.3325 20.02 4.745 20.06 ;
      RECT MASK 2 115.3515 20.14 129.1205 20.18 ;
      RECT MASK 2 1.3325 20.26 4.745 20.3 ;
      RECT MASK 2 115.3515 20.38 129.1205 20.42 ;
      RECT MASK 2 1.3325 20.5 4.745 20.54 ;
      RECT MASK 2 56.4625 20.54 58.3775 20.6 ;
      RECT MASK 2 115.3515 20.62 129.1205 20.66 ;
      RECT MASK 2 1.3325 20.74 4.745 20.78 ;
      RECT MASK 2 56.4625 20.78 58.3775 20.84 ;
      RECT MASK 2 115.3515 20.86 129.1205 20.9 ;
      RECT MASK 2 1.3325 20.98 4.745 21.02 ;
      RECT MASK 2 115.3515 21.1 129.1205 21.14 ;
      RECT MASK 2 1.3325 21.22 4.745 21.26 ;
      RECT MASK 2 115.3515 21.34 129.1205 21.38 ;
      RECT MASK 2 5.031 21.365 109.945 21.565 ;
      RECT MASK 2 1.3325 21.46 4.745 21.5 ;
      RECT MASK 2 115.3515 21.58 129.1205 21.62 ;
      RECT MASK 2 1.3325 21.7 4.745 21.74 ;
      RECT MASK 2 56.722 21.745 58.9155 21.805 ;
      RECT MASK 2 115.3515 21.82 129.1205 21.86 ;
      RECT MASK 2 1.3325 21.94 4.745 21.98 ;
      RECT MASK 2 115.3515 22.06 129.1205 22.1 ;
      RECT MASK 2 1.3325 22.18 4.745 22.22 ;
      RECT MASK 2 5.779 22.29 6.105 22.35 ;
      RECT MASK 2 6.941 22.29 7.267 22.35 ;
      RECT MASK 2 8.103 22.29 8.429 22.35 ;
      RECT MASK 2 9.265 22.29 9.591 22.35 ;
      RECT MASK 2 12.397 22.29 12.723 22.35 ;
      RECT MASK 2 13.559 22.29 13.885 22.35 ;
      RECT MASK 2 14.721 22.29 15.047 22.35 ;
      RECT MASK 2 15.883 22.29 16.209 22.35 ;
      RECT MASK 2 19.015 22.29 19.341 22.35 ;
      RECT MASK 2 20.177 22.29 20.503 22.35 ;
      RECT MASK 2 21.339 22.29 21.665 22.35 ;
      RECT MASK 2 22.501 22.29 22.827 22.35 ;
      RECT MASK 2 25.633 22.29 25.959 22.35 ;
      RECT MASK 2 26.795 22.29 27.121 22.35 ;
      RECT MASK 2 27.957 22.29 28.283 22.35 ;
      RECT MASK 2 29.119 22.29 29.445 22.35 ;
      RECT MASK 2 32.251 22.29 32.577 22.35 ;
      RECT MASK 2 33.413 22.29 33.739 22.35 ;
      RECT MASK 2 34.575 22.29 34.901 22.35 ;
      RECT MASK 2 35.737 22.29 36.063 22.35 ;
      RECT MASK 2 38.869 22.29 39.195 22.35 ;
      RECT MASK 2 40.031 22.29 40.357 22.35 ;
      RECT MASK 2 41.193 22.29 41.519 22.35 ;
      RECT MASK 2 42.355 22.29 42.681 22.35 ;
      RECT MASK 2 45.487 22.29 45.813 22.35 ;
      RECT MASK 2 46.649 22.29 46.975 22.35 ;
      RECT MASK 2 47.811 22.29 48.137 22.35 ;
      RECT MASK 2 48.973 22.29 49.299 22.35 ;
      RECT MASK 2 52.105 22.29 52.431 22.35 ;
      RECT MASK 2 53.267 22.29 53.593 22.35 ;
      RECT MASK 2 54.429 22.29 54.755 22.35 ;
      RECT MASK 2 55.591 22.29 55.917 22.35 ;
      RECT MASK 2 58.723 22.29 59.049 22.35 ;
      RECT MASK 2 59.885 22.29 60.211 22.35 ;
      RECT MASK 2 61.047 22.29 61.373 22.35 ;
      RECT MASK 2 62.209 22.29 62.535 22.35 ;
      RECT MASK 2 65.341 22.29 65.667 22.35 ;
      RECT MASK 2 66.503 22.29 66.829 22.35 ;
      RECT MASK 2 67.665 22.29 67.991 22.35 ;
      RECT MASK 2 68.827 22.29 69.153 22.35 ;
      RECT MASK 2 71.959 22.29 72.285 22.35 ;
      RECT MASK 2 73.121 22.29 73.447 22.35 ;
      RECT MASK 2 74.283 22.29 74.609 22.35 ;
      RECT MASK 2 75.445 22.29 75.771 22.35 ;
      RECT MASK 2 78.577 22.29 78.903 22.35 ;
      RECT MASK 2 79.739 22.29 80.065 22.35 ;
      RECT MASK 2 80.901 22.29 81.227 22.35 ;
      RECT MASK 2 82.063 22.29 82.389 22.35 ;
      RECT MASK 2 85.195 22.29 85.521 22.35 ;
      RECT MASK 2 86.357 22.29 86.683 22.35 ;
      RECT MASK 2 87.519 22.29 87.845 22.35 ;
      RECT MASK 2 88.681 22.29 89.007 22.35 ;
      RECT MASK 2 91.813 22.29 92.139 22.35 ;
      RECT MASK 2 92.975 22.29 93.301 22.35 ;
      RECT MASK 2 94.137 22.29 94.463 22.35 ;
      RECT MASK 2 95.299 22.29 95.625 22.35 ;
      RECT MASK 2 98.431 22.29 98.757 22.35 ;
      RECT MASK 2 99.593 22.29 99.919 22.35 ;
      RECT MASK 2 100.755 22.29 101.081 22.35 ;
      RECT MASK 2 101.917 22.29 102.243 22.35 ;
      RECT MASK 2 105.049 22.29 105.375 22.35 ;
      RECT MASK 2 106.211 22.29 106.537 22.35 ;
      RECT MASK 2 107.373 22.29 107.699 22.35 ;
      RECT MASK 2 108.535 22.29 108.861 22.35 ;
      RECT MASK 2 115.3515 22.3 129.1205 22.34 ;
      RECT MASK 2 1.3325 22.42 4.745 22.46 ;
      RECT MASK 2 115.3515 22.54 129.1205 22.58 ;
      RECT MASK 2 1.3325 22.66 4.745 22.7 ;
      RECT MASK 2 5.779 22.77 6.105 22.83 ;
      RECT MASK 2 6.941 22.77 7.267 22.83 ;
      RECT MASK 2 8.103 22.77 8.429 22.83 ;
      RECT MASK 2 9.265 22.77 9.591 22.83 ;
      RECT MASK 2 12.397 22.77 12.723 22.83 ;
      RECT MASK 2 13.559 22.77 13.885 22.83 ;
      RECT MASK 2 14.721 22.77 15.047 22.83 ;
      RECT MASK 2 15.883 22.77 16.209 22.83 ;
      RECT MASK 2 19.015 22.77 19.341 22.83 ;
      RECT MASK 2 20.177 22.77 20.503 22.83 ;
      RECT MASK 2 21.339 22.77 21.665 22.83 ;
      RECT MASK 2 22.501 22.77 22.827 22.83 ;
      RECT MASK 2 25.633 22.77 25.959 22.83 ;
      RECT MASK 2 26.795 22.77 27.121 22.83 ;
      RECT MASK 2 27.957 22.77 28.283 22.83 ;
      RECT MASK 2 29.119 22.77 29.445 22.83 ;
      RECT MASK 2 32.251 22.77 32.577 22.83 ;
      RECT MASK 2 33.413 22.77 33.739 22.83 ;
      RECT MASK 2 34.575 22.77 34.901 22.83 ;
      RECT MASK 2 35.737 22.77 36.063 22.83 ;
      RECT MASK 2 38.869 22.77 39.195 22.83 ;
      RECT MASK 2 40.031 22.77 40.357 22.83 ;
      RECT MASK 2 41.193 22.77 41.519 22.83 ;
      RECT MASK 2 42.355 22.77 42.681 22.83 ;
      RECT MASK 2 45.487 22.77 45.813 22.83 ;
      RECT MASK 2 46.649 22.77 46.975 22.83 ;
      RECT MASK 2 47.811 22.77 48.137 22.83 ;
      RECT MASK 2 48.973 22.77 49.299 22.83 ;
      RECT MASK 2 52.105 22.77 52.431 22.83 ;
      RECT MASK 2 53.267 22.77 53.593 22.83 ;
      RECT MASK 2 54.429 22.77 54.755 22.83 ;
      RECT MASK 2 55.591 22.77 55.917 22.83 ;
      RECT MASK 2 58.723 22.77 59.049 22.83 ;
      RECT MASK 2 59.885 22.77 60.211 22.83 ;
      RECT MASK 2 61.047 22.77 61.373 22.83 ;
      RECT MASK 2 62.209 22.77 62.535 22.83 ;
      RECT MASK 2 65.341 22.77 65.667 22.83 ;
      RECT MASK 2 66.503 22.77 66.829 22.83 ;
      RECT MASK 2 67.665 22.77 67.991 22.83 ;
      RECT MASK 2 68.827 22.77 69.153 22.83 ;
      RECT MASK 2 71.959 22.77 72.285 22.83 ;
      RECT MASK 2 73.121 22.77 73.447 22.83 ;
      RECT MASK 2 74.283 22.77 74.609 22.83 ;
      RECT MASK 2 75.445 22.77 75.771 22.83 ;
      RECT MASK 2 78.577 22.77 78.903 22.83 ;
      RECT MASK 2 79.739 22.77 80.065 22.83 ;
      RECT MASK 2 80.901 22.77 81.227 22.83 ;
      RECT MASK 2 82.063 22.77 82.389 22.83 ;
      RECT MASK 2 85.195 22.77 85.521 22.83 ;
      RECT MASK 2 86.357 22.77 86.683 22.83 ;
      RECT MASK 2 87.519 22.77 87.845 22.83 ;
      RECT MASK 2 88.681 22.77 89.007 22.83 ;
      RECT MASK 2 91.813 22.77 92.139 22.83 ;
      RECT MASK 2 92.975 22.77 93.301 22.83 ;
      RECT MASK 2 94.137 22.77 94.463 22.83 ;
      RECT MASK 2 95.299 22.77 95.625 22.83 ;
      RECT MASK 2 98.431 22.77 98.757 22.83 ;
      RECT MASK 2 99.593 22.77 99.919 22.83 ;
      RECT MASK 2 100.755 22.77 101.081 22.83 ;
      RECT MASK 2 101.917 22.77 102.243 22.83 ;
      RECT MASK 2 105.049 22.77 105.375 22.83 ;
      RECT MASK 2 106.211 22.77 106.537 22.83 ;
      RECT MASK 2 107.373 22.77 107.699 22.83 ;
      RECT MASK 2 108.535 22.77 108.861 22.83 ;
      RECT MASK 2 115.3515 22.78 129.1205 22.82 ;
      RECT MASK 2 1.3325 22.9 4.745 22.94 ;
      RECT MASK 2 115.3515 23.02 129.1205 23.06 ;
      RECT MASK 2 1.3325 23.14 4.745 23.18 ;
      RECT MASK 2 115.3515 23.26 129.1205 23.3 ;
      RECT MASK 2 5.319 23.355 10.382 23.475 ;
      RECT MASK 2 11.937 23.355 17 23.475 ;
      RECT MASK 2 18.555 23.355 23.618 23.475 ;
      RECT MASK 2 25.173 23.355 30.236 23.475 ;
      RECT MASK 2 31.791 23.355 36.854 23.475 ;
      RECT MASK 2 38.409 23.355 43.472 23.475 ;
      RECT MASK 2 45.027 23.355 50.09 23.475 ;
      RECT MASK 2 51.645 23.355 56.708 23.475 ;
      RECT MASK 2 58.263 23.355 63.326 23.475 ;
      RECT MASK 2 64.881 23.355 69.944 23.475 ;
      RECT MASK 2 71.499 23.355 76.562 23.475 ;
      RECT MASK 2 78.117 23.355 83.18 23.475 ;
      RECT MASK 2 84.735 23.355 89.798 23.475 ;
      RECT MASK 2 91.353 23.355 96.416 23.475 ;
      RECT MASK 2 97.971 23.355 103.034 23.475 ;
      RECT MASK 2 104.589 23.355 109.652 23.475 ;
      RECT MASK 2 1.3325 23.38 4.745 23.42 ;
      RECT MASK 2 1.3325 23.62 4.745 23.66 ;
      RECT MASK 2 5.319 23.805 10.382 23.925 ;
      RECT MASK 2 11.937 23.805 17 23.925 ;
      RECT MASK 2 18.555 23.805 23.618 23.925 ;
      RECT MASK 2 25.173 23.805 30.236 23.925 ;
      RECT MASK 2 31.791 23.805 36.854 23.925 ;
      RECT MASK 2 38.409 23.805 43.472 23.925 ;
      RECT MASK 2 45.027 23.805 50.09 23.925 ;
      RECT MASK 2 51.645 23.805 56.708 23.925 ;
      RECT MASK 2 58.263 23.805 63.326 23.925 ;
      RECT MASK 2 64.881 23.805 69.944 23.925 ;
      RECT MASK 2 71.499 23.805 76.562 23.925 ;
      RECT MASK 2 78.117 23.805 83.18 23.925 ;
      RECT MASK 2 84.735 23.805 89.798 23.925 ;
      RECT MASK 2 91.353 23.805 96.416 23.925 ;
      RECT MASK 2 97.971 23.805 103.034 23.925 ;
      RECT MASK 2 104.589 23.805 109.652 23.925 ;
      RECT MASK 2 1.3325 23.86 4.745 23.9 ;
      RECT MASK 2 1.3325 24.1 4.745 24.14 ;
      RECT MASK 2 2.327 24.34 3.827 24.38 ;
      RECT MASK 2 5.779 24.689 6.105 24.749 ;
      RECT MASK 2 6.941 24.689 7.267 24.749 ;
      RECT MASK 2 8.103 24.689 8.429 24.749 ;
      RECT MASK 2 9.265 24.689 9.591 24.749 ;
      RECT MASK 2 12.397 24.689 12.723 24.749 ;
      RECT MASK 2 13.559 24.689 13.885 24.749 ;
      RECT MASK 2 14.721 24.689 15.047 24.749 ;
      RECT MASK 2 15.883 24.689 16.209 24.749 ;
      RECT MASK 2 19.015 24.689 19.341 24.749 ;
      RECT MASK 2 20.177 24.689 20.503 24.749 ;
      RECT MASK 2 21.339 24.689 21.665 24.749 ;
      RECT MASK 2 22.501 24.689 22.827 24.749 ;
      RECT MASK 2 25.633 24.689 25.959 24.749 ;
      RECT MASK 2 26.795 24.689 27.121 24.749 ;
      RECT MASK 2 27.957 24.689 28.283 24.749 ;
      RECT MASK 2 29.119 24.689 29.445 24.749 ;
      RECT MASK 2 32.251 24.689 32.577 24.749 ;
      RECT MASK 2 33.413 24.689 33.739 24.749 ;
      RECT MASK 2 34.575 24.689 34.901 24.749 ;
      RECT MASK 2 35.737 24.689 36.063 24.749 ;
      RECT MASK 2 38.869 24.689 39.195 24.749 ;
      RECT MASK 2 40.031 24.689 40.357 24.749 ;
      RECT MASK 2 41.193 24.689 41.519 24.749 ;
      RECT MASK 2 42.355 24.689 42.681 24.749 ;
      RECT MASK 2 45.487 24.689 45.813 24.749 ;
      RECT MASK 2 46.649 24.689 46.975 24.749 ;
      RECT MASK 2 47.811 24.689 48.137 24.749 ;
      RECT MASK 2 48.973 24.689 49.299 24.749 ;
      RECT MASK 2 52.105 24.689 52.431 24.749 ;
      RECT MASK 2 53.267 24.689 53.593 24.749 ;
      RECT MASK 2 54.429 24.689 54.755 24.749 ;
      RECT MASK 2 55.591 24.689 55.917 24.749 ;
      RECT MASK 2 58.723 24.689 59.049 24.749 ;
      RECT MASK 2 59.885 24.689 60.211 24.749 ;
      RECT MASK 2 61.047 24.689 61.373 24.749 ;
      RECT MASK 2 62.209 24.689 62.535 24.749 ;
      RECT MASK 2 65.341 24.689 65.667 24.749 ;
      RECT MASK 2 66.503 24.689 66.829 24.749 ;
      RECT MASK 2 67.665 24.689 67.991 24.749 ;
      RECT MASK 2 68.827 24.689 69.153 24.749 ;
      RECT MASK 2 71.959 24.689 72.285 24.749 ;
      RECT MASK 2 73.121 24.689 73.447 24.749 ;
      RECT MASK 2 74.283 24.689 74.609 24.749 ;
      RECT MASK 2 75.445 24.689 75.771 24.749 ;
      RECT MASK 2 78.577 24.689 78.903 24.749 ;
      RECT MASK 2 79.739 24.689 80.065 24.749 ;
      RECT MASK 2 80.901 24.689 81.227 24.749 ;
      RECT MASK 2 82.063 24.689 82.389 24.749 ;
      RECT MASK 2 85.195 24.689 85.521 24.749 ;
      RECT MASK 2 86.357 24.689 86.683 24.749 ;
      RECT MASK 2 87.519 24.689 87.845 24.749 ;
      RECT MASK 2 88.681 24.689 89.007 24.749 ;
      RECT MASK 2 91.813 24.689 92.139 24.749 ;
      RECT MASK 2 92.975 24.689 93.301 24.749 ;
      RECT MASK 2 94.137 24.689 94.463 24.749 ;
      RECT MASK 2 95.299 24.689 95.625 24.749 ;
      RECT MASK 2 98.431 24.689 98.757 24.749 ;
      RECT MASK 2 99.593 24.689 99.919 24.749 ;
      RECT MASK 2 100.755 24.689 101.081 24.749 ;
      RECT MASK 2 101.917 24.689 102.243 24.749 ;
      RECT MASK 2 105.049 24.689 105.375 24.749 ;
      RECT MASK 2 106.211 24.689 106.537 24.749 ;
      RECT MASK 2 107.373 24.689 107.699 24.749 ;
      RECT MASK 2 108.535 24.689 108.861 24.749 ;
      RECT MASK 2 5.779 25.169 6.0885 25.229 ;
      RECT MASK 2 6.941 25.169 7.2505 25.229 ;
      RECT MASK 2 8.103 25.169 8.4125 25.229 ;
      RECT MASK 2 9.265 25.169 9.5745 25.229 ;
      RECT MASK 2 12.397 25.169 12.7065 25.229 ;
      RECT MASK 2 13.559 25.169 13.8685 25.229 ;
      RECT MASK 2 14.721 25.169 15.0305 25.229 ;
      RECT MASK 2 15.883 25.169 16.1925 25.229 ;
      RECT MASK 2 19.015 25.169 19.3245 25.229 ;
      RECT MASK 2 20.177 25.169 20.4865 25.229 ;
      RECT MASK 2 21.339 25.169 21.6485 25.229 ;
      RECT MASK 2 22.501 25.169 22.8105 25.229 ;
      RECT MASK 2 25.633 25.169 25.9425 25.229 ;
      RECT MASK 2 26.795 25.169 27.1045 25.229 ;
      RECT MASK 2 27.957 25.169 28.2665 25.229 ;
      RECT MASK 2 29.119 25.169 29.4285 25.229 ;
      RECT MASK 2 32.251 25.169 32.5605 25.229 ;
      RECT MASK 2 33.413 25.169 33.7225 25.229 ;
      RECT MASK 2 34.575 25.169 34.8845 25.229 ;
      RECT MASK 2 35.737 25.169 36.0465 25.229 ;
      RECT MASK 2 38.869 25.169 39.1785 25.229 ;
      RECT MASK 2 40.031 25.169 40.3405 25.229 ;
      RECT MASK 2 41.193 25.169 41.5025 25.229 ;
      RECT MASK 2 42.355 25.169 42.6645 25.229 ;
      RECT MASK 2 45.487 25.169 45.7965 25.229 ;
      RECT MASK 2 46.649 25.169 46.9585 25.229 ;
      RECT MASK 2 47.811 25.169 48.1205 25.229 ;
      RECT MASK 2 48.973 25.169 49.2825 25.229 ;
      RECT MASK 2 52.105 25.169 52.4145 25.229 ;
      RECT MASK 2 53.267 25.169 53.5765 25.229 ;
      RECT MASK 2 54.429 25.169 54.7385 25.229 ;
      RECT MASK 2 55.591 25.169 55.9005 25.229 ;
      RECT MASK 2 58.723 25.169 59.0325 25.229 ;
      RECT MASK 2 59.885 25.169 60.1945 25.229 ;
      RECT MASK 2 61.047 25.169 61.3565 25.229 ;
      RECT MASK 2 62.209 25.169 62.5185 25.229 ;
      RECT MASK 2 65.341 25.169 65.6505 25.229 ;
      RECT MASK 2 66.503 25.169 66.8125 25.229 ;
      RECT MASK 2 67.665 25.169 67.9745 25.229 ;
      RECT MASK 2 68.827 25.169 69.1365 25.229 ;
      RECT MASK 2 71.959 25.169 72.2685 25.229 ;
      RECT MASK 2 73.121 25.169 73.4305 25.229 ;
      RECT MASK 2 74.283 25.169 74.5925 25.229 ;
      RECT MASK 2 75.445 25.169 75.7545 25.229 ;
      RECT MASK 2 78.577 25.169 78.8865 25.229 ;
      RECT MASK 2 79.739 25.169 80.0485 25.229 ;
      RECT MASK 2 80.901 25.169 81.2105 25.229 ;
      RECT MASK 2 82.063 25.169 82.3725 25.229 ;
      RECT MASK 2 85.195 25.169 85.5045 25.229 ;
      RECT MASK 2 86.357 25.169 86.6665 25.229 ;
      RECT MASK 2 87.519 25.169 87.8285 25.229 ;
      RECT MASK 2 88.681 25.169 88.9905 25.229 ;
      RECT MASK 2 91.813 25.169 92.1225 25.229 ;
      RECT MASK 2 92.975 25.169 93.2845 25.229 ;
      RECT MASK 2 94.137 25.169 94.4465 25.229 ;
      RECT MASK 2 95.299 25.169 95.6085 25.229 ;
      RECT MASK 2 98.431 25.169 98.7405 25.229 ;
      RECT MASK 2 99.593 25.169 99.9025 25.229 ;
      RECT MASK 2 100.755 25.169 101.0645 25.229 ;
      RECT MASK 2 101.917 25.169 102.2265 25.229 ;
      RECT MASK 2 105.049 25.169 105.3585 25.229 ;
      RECT MASK 2 106.211 25.169 106.5205 25.229 ;
      RECT MASK 2 107.373 25.169 107.6825 25.229 ;
      RECT MASK 2 108.535 25.169 108.8445 25.229 ;
      RECT MASK 2 5.031 25.725 109.945 25.905 ;
      RECT MASK 2 113.368 27.2 126.9585 27.4 ;
      RECT MASK 2 116.318 27.72 126.334 27.92 ;
      RECT MASK 2 116.074 28.32 126.333 28.38 ;
      RECT MASK 2 4.672 28.465 17.578 28.565 ;
      RECT MASK 2 17.908 28.465 30.814 28.565 ;
      RECT MASK 2 31.144 28.465 44.05 28.565 ;
      RECT MASK 2 44.38 28.465 57.286 28.565 ;
      RECT MASK 2 57.616 28.465 70.522 28.565 ;
      RECT MASK 2 70.852 28.465 83.758 28.565 ;
      RECT MASK 2 84.088 28.465 96.994 28.565 ;
      RECT MASK 2 97.324 28.465 110.23 28.565 ;
      RECT MASK 2 116.2095 28.76 126.3345 28.96 ;
      RECT MASK 2 4.656 28.84 17.604 28.94 ;
      RECT MASK 2 17.892 28.84 30.84 28.94 ;
      RECT MASK 2 31.128 28.84 44.076 28.94 ;
      RECT MASK 2 44.364 28.84 57.312 28.94 ;
      RECT MASK 2 57.6 28.84 70.548 28.94 ;
      RECT MASK 2 70.836 28.84 83.784 28.94 ;
      RECT MASK 2 84.072 28.84 97.02 28.94 ;
      RECT MASK 2 97.308 28.84 110.256 28.94 ;
      RECT MASK 2 4.672 29.215 17.578 29.315 ;
      RECT MASK 2 17.908 29.215 30.814 29.315 ;
      RECT MASK 2 31.144 29.215 44.05 29.315 ;
      RECT MASK 2 44.38 29.215 57.286 29.315 ;
      RECT MASK 2 57.616 29.215 70.522 29.315 ;
      RECT MASK 2 70.852 29.215 83.758 29.315 ;
      RECT MASK 2 84.088 29.215 96.994 29.315 ;
      RECT MASK 2 97.324 29.215 110.23 29.315 ;
      RECT MASK 2 116.318 29.28 126.334 29.48 ;
      RECT MASK 2 4.672 29.585 17.578 29.685 ;
      RECT MASK 2 17.908 29.585 30.814 29.685 ;
      RECT MASK 2 31.144 29.585 44.05 29.685 ;
      RECT MASK 2 44.38 29.585 57.286 29.685 ;
      RECT MASK 2 57.616 29.585 70.522 29.685 ;
      RECT MASK 2 70.852 29.585 83.758 29.685 ;
      RECT MASK 2 84.088 29.585 96.994 29.685 ;
      RECT MASK 2 97.324 29.585 110.23 29.685 ;
      RECT MASK 2 4.656 29.96 17.604 30.06 ;
      RECT MASK 2 17.892 29.96 30.84 30.06 ;
      RECT MASK 2 31.128 29.96 44.076 30.06 ;
      RECT MASK 2 44.364 29.96 57.312 30.06 ;
      RECT MASK 2 57.6 29.96 70.548 30.06 ;
      RECT MASK 2 70.836 29.96 83.784 30.06 ;
      RECT MASK 2 84.072 29.96 97.02 30.06 ;
      RECT MASK 2 97.308 29.96 110.256 30.06 ;
      RECT MASK 2 4.672 30.335 17.578 30.435 ;
      RECT MASK 2 17.908 30.335 30.814 30.435 ;
      RECT MASK 2 31.144 30.335 44.05 30.435 ;
      RECT MASK 2 44.38 30.335 57.286 30.435 ;
      RECT MASK 2 57.616 30.335 70.522 30.435 ;
      RECT MASK 2 70.852 30.335 83.758 30.435 ;
      RECT MASK 2 84.088 30.335 96.994 30.435 ;
      RECT MASK 2 97.324 30.335 110.23 30.435 ;
      RECT MASK 2 4.672 30.705 17.578 30.805 ;
      RECT MASK 2 17.908 30.705 30.814 30.805 ;
      RECT MASK 2 31.144 30.705 44.05 30.805 ;
      RECT MASK 2 44.38 30.705 57.286 30.805 ;
      RECT MASK 2 57.616 30.705 70.522 30.805 ;
      RECT MASK 2 70.852 30.705 83.758 30.805 ;
      RECT MASK 2 84.088 30.705 96.994 30.805 ;
      RECT MASK 2 97.324 30.705 110.23 30.805 ;
      RECT MASK 2 4.656 31.08 17.604 31.18 ;
      RECT MASK 2 17.892 31.08 30.84 31.18 ;
      RECT MASK 2 31.128 31.08 44.076 31.18 ;
      RECT MASK 2 44.364 31.08 57.312 31.18 ;
      RECT MASK 2 57.6 31.08 70.548 31.18 ;
      RECT MASK 2 70.836 31.08 83.784 31.18 ;
      RECT MASK 2 84.072 31.08 97.02 31.18 ;
      RECT MASK 2 97.308 31.08 110.256 31.18 ;
      RECT MASK 2 111.0245 31.245 129.1315 31.365 ;
      RECT MASK 2 4.672 31.455 17.578 31.555 ;
      RECT MASK 2 17.908 31.455 30.814 31.555 ;
      RECT MASK 2 31.144 31.455 44.05 31.555 ;
      RECT MASK 2 44.38 31.455 57.286 31.555 ;
      RECT MASK 2 57.616 31.455 70.522 31.555 ;
      RECT MASK 2 70.852 31.455 83.758 31.555 ;
      RECT MASK 2 84.088 31.455 96.994 31.555 ;
      RECT MASK 2 97.324 31.455 110.23 31.555 ;
      RECT MASK 2 4.672 31.825 17.578 31.925 ;
      RECT MASK 2 17.908 31.825 30.814 31.925 ;
      RECT MASK 2 31.144 31.825 44.05 31.925 ;
      RECT MASK 2 44.38 31.825 57.286 31.925 ;
      RECT MASK 2 57.616 31.825 70.522 31.925 ;
      RECT MASK 2 70.852 31.825 83.758 31.925 ;
      RECT MASK 2 84.088 31.825 96.994 31.925 ;
      RECT MASK 2 97.324 31.825 110.23 31.925 ;
      RECT MASK 2 113.0865 32.1375 127.58 32.3875 ;
      RECT MASK 2 4.656 32.2 17.604 32.3 ;
      RECT MASK 2 17.892 32.2 30.84 32.3 ;
      RECT MASK 2 31.128 32.2 44.076 32.3 ;
      RECT MASK 2 44.364 32.2 57.312 32.3 ;
      RECT MASK 2 57.6 32.2 70.548 32.3 ;
      RECT MASK 2 70.836 32.2 83.784 32.3 ;
      RECT MASK 2 84.072 32.2 97.02 32.3 ;
      RECT MASK 2 97.308 32.2 110.256 32.3 ;
      RECT MASK 2 4.672 32.575 17.578 32.675 ;
      RECT MASK 2 17.908 32.575 30.814 32.675 ;
      RECT MASK 2 31.144 32.575 44.05 32.675 ;
      RECT MASK 2 44.38 32.575 57.286 32.675 ;
      RECT MASK 2 57.616 32.575 70.522 32.675 ;
      RECT MASK 2 70.852 32.575 83.758 32.675 ;
      RECT MASK 2 84.088 32.575 96.994 32.675 ;
      RECT MASK 2 97.324 32.575 110.23 32.675 ;
      RECT MASK 2 117.268 32.9125 129.1315 33.1625 ;
      RECT MASK 2 0.567 33.33 115.126 33.45 ;
      RECT MASK 2 117.268 33.6175 129.1315 33.8675 ;
      RECT MASK 2 0.567 33.75 115.126 33.87 ;
      RECT MASK 2 111.044 34.1325 129.1315 34.2325 ;
      RECT MASK 2 4.672 34.555 10.96 34.655 ;
      RECT MASK 2 11.29 34.555 17.578 34.655 ;
      RECT MASK 2 17.908 34.555 24.196 34.655 ;
      RECT MASK 2 24.526 34.555 30.814 34.655 ;
      RECT MASK 2 31.144 34.555 37.432 34.655 ;
      RECT MASK 2 37.762 34.555 44.05 34.655 ;
      RECT MASK 2 44.38 34.555 50.668 34.655 ;
      RECT MASK 2 50.998 34.555 57.286 34.655 ;
      RECT MASK 2 57.616 34.555 63.904 34.655 ;
      RECT MASK 2 64.234 34.555 70.522 34.655 ;
      RECT MASK 2 70.852 34.555 77.14 34.655 ;
      RECT MASK 2 77.47 34.555 83.758 34.655 ;
      RECT MASK 2 84.088 34.555 90.376 34.655 ;
      RECT MASK 2 90.706 34.555 96.994 34.655 ;
      RECT MASK 2 97.324 34.555 103.612 34.655 ;
      RECT MASK 2 103.942 34.555 110.23 34.655 ;
      RECT MASK 2 111.044 34.6475 127.58 34.7475 ;
      RECT MASK 2 4.656 34.93 10.986 35.03 ;
      RECT MASK 2 11.274 34.93 17.604 35.03 ;
      RECT MASK 2 17.892 34.93 24.222 35.03 ;
      RECT MASK 2 24.51 34.93 30.84 35.03 ;
      RECT MASK 2 31.128 34.93 37.458 35.03 ;
      RECT MASK 2 37.746 34.93 44.076 35.03 ;
      RECT MASK 2 44.364 34.93 50.694 35.03 ;
      RECT MASK 2 50.982 34.93 57.312 35.03 ;
      RECT MASK 2 57.6 34.93 63.93 35.03 ;
      RECT MASK 2 64.218 34.93 70.548 35.03 ;
      RECT MASK 2 70.836 34.93 77.166 35.03 ;
      RECT MASK 2 77.454 34.93 83.784 35.03 ;
      RECT MASK 2 84.072 34.93 90.402 35.03 ;
      RECT MASK 2 90.69 34.93 97.02 35.03 ;
      RECT MASK 2 97.308 34.93 103.638 35.03 ;
      RECT MASK 2 103.926 34.93 110.256 35.03 ;
      RECT MASK 2 111.044 34.9675 129.1315 35.2175 ;
      RECT MASK 2 4.672 35.305 10.96 35.405 ;
      RECT MASK 2 11.29 35.305 17.578 35.405 ;
      RECT MASK 2 17.908 35.305 24.196 35.405 ;
      RECT MASK 2 24.526 35.305 30.814 35.405 ;
      RECT MASK 2 31.144 35.305 37.432 35.405 ;
      RECT MASK 2 37.762 35.305 44.05 35.405 ;
      RECT MASK 2 44.38 35.305 50.668 35.405 ;
      RECT MASK 2 50.998 35.305 57.286 35.405 ;
      RECT MASK 2 57.616 35.305 63.904 35.405 ;
      RECT MASK 2 64.234 35.305 70.522 35.405 ;
      RECT MASK 2 70.852 35.305 77.14 35.405 ;
      RECT MASK 2 77.47 35.305 83.758 35.405 ;
      RECT MASK 2 84.088 35.305 90.376 35.405 ;
      RECT MASK 2 90.706 35.305 96.994 35.405 ;
      RECT MASK 2 97.324 35.305 103.612 35.405 ;
      RECT MASK 2 103.942 35.305 110.23 35.405 ;
      RECT MASK 2 111.044 35.4825 129.1315 35.5825 ;
      RECT MASK 2 4.672 35.675 10.96 35.775 ;
      RECT MASK 2 11.29 35.675 17.578 35.775 ;
      RECT MASK 2 17.908 35.675 24.196 35.775 ;
      RECT MASK 2 24.526 35.675 30.814 35.775 ;
      RECT MASK 2 31.144 35.675 37.432 35.775 ;
      RECT MASK 2 37.762 35.675 44.05 35.775 ;
      RECT MASK 2 44.38 35.675 50.668 35.775 ;
      RECT MASK 2 50.998 35.675 57.286 35.775 ;
      RECT MASK 2 57.616 35.675 63.904 35.775 ;
      RECT MASK 2 64.234 35.675 70.522 35.775 ;
      RECT MASK 2 70.852 35.675 77.14 35.775 ;
      RECT MASK 2 77.47 35.675 83.758 35.775 ;
      RECT MASK 2 84.088 35.675 90.376 35.775 ;
      RECT MASK 2 90.706 35.675 96.994 35.775 ;
      RECT MASK 2 97.324 35.675 103.612 35.775 ;
      RECT MASK 2 103.942 35.675 110.23 35.775 ;
      RECT MASK 2 111.044 35.9975 127.58 36.0975 ;
      RECT MASK 2 4.656 36.05 10.986 36.15 ;
      RECT MASK 2 11.274 36.05 17.604 36.15 ;
      RECT MASK 2 17.892 36.05 24.222 36.15 ;
      RECT MASK 2 24.51 36.05 30.84 36.15 ;
      RECT MASK 2 31.128 36.05 37.458 36.15 ;
      RECT MASK 2 37.746 36.05 44.076 36.15 ;
      RECT MASK 2 44.364 36.05 50.694 36.15 ;
      RECT MASK 2 50.982 36.05 57.312 36.15 ;
      RECT MASK 2 57.6 36.05 63.93 36.15 ;
      RECT MASK 2 64.218 36.05 70.548 36.15 ;
      RECT MASK 2 70.836 36.05 77.166 36.15 ;
      RECT MASK 2 77.454 36.05 83.784 36.15 ;
      RECT MASK 2 84.072 36.05 90.402 36.15 ;
      RECT MASK 2 90.69 36.05 97.02 36.15 ;
      RECT MASK 2 97.308 36.05 103.638 36.15 ;
      RECT MASK 2 103.926 36.05 110.256 36.15 ;
      RECT MASK 2 111.044 36.3175 129.1315 36.5675 ;
      RECT MASK 2 4.672 36.425 10.96 36.525 ;
      RECT MASK 2 11.29 36.425 17.578 36.525 ;
      RECT MASK 2 17.908 36.425 24.196 36.525 ;
      RECT MASK 2 24.526 36.425 30.814 36.525 ;
      RECT MASK 2 31.144 36.425 37.432 36.525 ;
      RECT MASK 2 37.762 36.425 44.05 36.525 ;
      RECT MASK 2 44.38 36.425 50.668 36.525 ;
      RECT MASK 2 50.998 36.425 57.286 36.525 ;
      RECT MASK 2 57.616 36.425 63.904 36.525 ;
      RECT MASK 2 64.234 36.425 70.522 36.525 ;
      RECT MASK 2 70.852 36.425 77.14 36.525 ;
      RECT MASK 2 77.47 36.425 83.758 36.525 ;
      RECT MASK 2 84.088 36.425 90.376 36.525 ;
      RECT MASK 2 90.706 36.425 96.994 36.525 ;
      RECT MASK 2 97.324 36.425 103.612 36.525 ;
      RECT MASK 2 103.942 36.425 110.23 36.525 ;
      RECT MASK 2 4.672 36.795 10.96 36.895 ;
      RECT MASK 2 11.29 36.795 17.578 36.895 ;
      RECT MASK 2 17.908 36.795 24.196 36.895 ;
      RECT MASK 2 24.526 36.795 30.814 36.895 ;
      RECT MASK 2 31.144 36.795 37.432 36.895 ;
      RECT MASK 2 37.762 36.795 44.05 36.895 ;
      RECT MASK 2 44.38 36.795 50.668 36.895 ;
      RECT MASK 2 50.998 36.795 57.286 36.895 ;
      RECT MASK 2 57.616 36.795 63.904 36.895 ;
      RECT MASK 2 64.234 36.795 70.522 36.895 ;
      RECT MASK 2 70.852 36.795 77.14 36.895 ;
      RECT MASK 2 77.47 36.795 83.758 36.895 ;
      RECT MASK 2 84.088 36.795 90.376 36.895 ;
      RECT MASK 2 90.706 36.795 96.994 36.895 ;
      RECT MASK 2 97.324 36.795 103.612 36.895 ;
      RECT MASK 2 103.942 36.795 110.23 36.895 ;
      RECT MASK 2 111.044 36.8675 129.1315 36.9675 ;
      RECT MASK 2 4.656 37.17 10.986 37.27 ;
      RECT MASK 2 11.274 37.17 17.604 37.27 ;
      RECT MASK 2 17.892 37.17 24.222 37.27 ;
      RECT MASK 2 24.51 37.17 30.84 37.27 ;
      RECT MASK 2 31.128 37.17 37.458 37.27 ;
      RECT MASK 2 37.746 37.17 44.076 37.27 ;
      RECT MASK 2 44.364 37.17 50.694 37.27 ;
      RECT MASK 2 50.982 37.17 57.312 37.27 ;
      RECT MASK 2 57.6 37.17 63.93 37.27 ;
      RECT MASK 2 64.218 37.17 70.548 37.27 ;
      RECT MASK 2 70.836 37.17 77.166 37.27 ;
      RECT MASK 2 77.454 37.17 83.784 37.27 ;
      RECT MASK 2 84.072 37.17 90.402 37.27 ;
      RECT MASK 2 90.69 37.17 97.02 37.27 ;
      RECT MASK 2 97.308 37.17 103.638 37.27 ;
      RECT MASK 2 103.926 37.17 110.256 37.27 ;
      RECT MASK 2 111.044 37.3475 127.58 37.4475 ;
      RECT MASK 2 4.672 37.545 10.96 37.645 ;
      RECT MASK 2 11.29 37.545 17.578 37.645 ;
      RECT MASK 2 17.908 37.545 24.196 37.645 ;
      RECT MASK 2 24.526 37.545 30.814 37.645 ;
      RECT MASK 2 31.144 37.545 37.432 37.645 ;
      RECT MASK 2 37.762 37.545 44.05 37.645 ;
      RECT MASK 2 44.38 37.545 50.668 37.645 ;
      RECT MASK 2 50.998 37.545 57.286 37.645 ;
      RECT MASK 2 57.616 37.545 63.904 37.645 ;
      RECT MASK 2 64.234 37.545 70.522 37.645 ;
      RECT MASK 2 70.852 37.545 77.14 37.645 ;
      RECT MASK 2 77.47 37.545 83.758 37.645 ;
      RECT MASK 2 84.088 37.545 90.376 37.645 ;
      RECT MASK 2 90.706 37.545 96.994 37.645 ;
      RECT MASK 2 97.324 37.545 103.612 37.645 ;
      RECT MASK 2 103.942 37.545 110.23 37.645 ;
      RECT MASK 2 111.044 37.6675 129.1315 37.9175 ;
      RECT MASK 2 4.672 37.915 10.96 38.015 ;
      RECT MASK 2 11.29 37.915 17.578 38.015 ;
      RECT MASK 2 17.908 37.915 24.196 38.015 ;
      RECT MASK 2 24.526 37.915 30.814 38.015 ;
      RECT MASK 2 31.144 37.915 37.432 38.015 ;
      RECT MASK 2 37.762 37.915 44.05 38.015 ;
      RECT MASK 2 44.38 37.915 50.668 38.015 ;
      RECT MASK 2 50.998 37.915 57.286 38.015 ;
      RECT MASK 2 57.616 37.915 63.904 38.015 ;
      RECT MASK 2 64.234 37.915 70.522 38.015 ;
      RECT MASK 2 70.852 37.915 77.14 38.015 ;
      RECT MASK 2 77.47 37.915 83.758 38.015 ;
      RECT MASK 2 84.088 37.915 90.376 38.015 ;
      RECT MASK 2 90.706 37.915 96.994 38.015 ;
      RECT MASK 2 97.324 37.915 103.612 38.015 ;
      RECT MASK 2 103.942 37.915 110.23 38.015 ;
      RECT MASK 2 111.044 38.1825 129.1315 38.2825 ;
      RECT MASK 2 4.656 38.29 10.986 38.39 ;
      RECT MASK 2 11.274 38.29 17.604 38.39 ;
      RECT MASK 2 17.892 38.29 24.222 38.39 ;
      RECT MASK 2 24.51 38.29 30.84 38.39 ;
      RECT MASK 2 31.128 38.29 37.458 38.39 ;
      RECT MASK 2 37.746 38.29 44.076 38.39 ;
      RECT MASK 2 44.364 38.29 50.694 38.39 ;
      RECT MASK 2 50.982 38.29 57.312 38.39 ;
      RECT MASK 2 57.6 38.29 63.93 38.39 ;
      RECT MASK 2 64.218 38.29 70.548 38.39 ;
      RECT MASK 2 70.836 38.29 77.166 38.39 ;
      RECT MASK 2 77.454 38.29 83.784 38.39 ;
      RECT MASK 2 84.072 38.29 90.402 38.39 ;
      RECT MASK 2 90.69 38.29 97.02 38.39 ;
      RECT MASK 2 97.308 38.29 103.638 38.39 ;
      RECT MASK 2 103.926 38.29 110.256 38.39 ;
      RECT MASK 2 4.672 38.665 10.96 38.765 ;
      RECT MASK 2 11.29 38.665 17.578 38.765 ;
      RECT MASK 2 17.908 38.665 24.196 38.765 ;
      RECT MASK 2 24.526 38.665 30.814 38.765 ;
      RECT MASK 2 31.144 38.665 37.432 38.765 ;
      RECT MASK 2 37.762 38.665 44.05 38.765 ;
      RECT MASK 2 44.38 38.665 50.668 38.765 ;
      RECT MASK 2 50.998 38.665 57.286 38.765 ;
      RECT MASK 2 57.616 38.665 63.904 38.765 ;
      RECT MASK 2 64.234 38.665 70.522 38.765 ;
      RECT MASK 2 70.852 38.665 77.14 38.765 ;
      RECT MASK 2 77.47 38.665 83.758 38.765 ;
      RECT MASK 2 84.088 38.665 90.376 38.765 ;
      RECT MASK 2 90.706 38.665 96.994 38.765 ;
      RECT MASK 2 97.324 38.665 103.612 38.765 ;
      RECT MASK 2 103.942 38.665 110.23 38.765 ;
      RECT MASK 2 111.044 38.6975 127.58 38.7975 ;
      RECT MASK 2 117.268 39.0175 129.1315 39.2675 ;
      RECT MASK 2 0.567 39.42 115.126 39.54 ;
      RECT MASK 2 117.268 39.5325 129.1315 39.6325 ;
      RECT MASK 2 0.567 39.84 115.126 39.96 ;
      RECT MASK 2 111.044 40.1075 127.58 40.2075 ;
      RECT MASK 2 111.044 40.4275 129.1315 40.6775 ;
      RECT MASK 2 4.672 40.675 10.96 40.775 ;
      RECT MASK 2 11.29 40.675 17.578 40.775 ;
      RECT MASK 2 17.908 40.675 24.196 40.775 ;
      RECT MASK 2 24.526 40.675 30.814 40.775 ;
      RECT MASK 2 31.144 40.675 37.432 40.775 ;
      RECT MASK 2 37.762 40.675 44.05 40.775 ;
      RECT MASK 2 44.38 40.675 50.668 40.775 ;
      RECT MASK 2 50.998 40.675 57.286 40.775 ;
      RECT MASK 2 57.616 40.675 63.904 40.775 ;
      RECT MASK 2 64.234 40.675 70.522 40.775 ;
      RECT MASK 2 70.852 40.675 77.14 40.775 ;
      RECT MASK 2 77.47 40.675 83.758 40.775 ;
      RECT MASK 2 84.088 40.675 90.376 40.775 ;
      RECT MASK 2 90.706 40.675 96.994 40.775 ;
      RECT MASK 2 97.324 40.675 103.612 40.775 ;
      RECT MASK 2 103.942 40.675 110.23 40.775 ;
      RECT MASK 2 111.044 40.9425 127.58 41.0425 ;
      RECT MASK 2 4.656 41.05 10.986 41.15 ;
      RECT MASK 2 11.274 41.05 17.604 41.15 ;
      RECT MASK 2 17.892 41.05 24.222 41.15 ;
      RECT MASK 2 24.51 41.05 30.84 41.15 ;
      RECT MASK 2 31.128 41.05 37.458 41.15 ;
      RECT MASK 2 37.746 41.05 44.076 41.15 ;
      RECT MASK 2 44.364 41.05 50.694 41.15 ;
      RECT MASK 2 50.982 41.05 57.312 41.15 ;
      RECT MASK 2 57.6 41.05 63.93 41.15 ;
      RECT MASK 2 64.218 41.05 70.548 41.15 ;
      RECT MASK 2 70.836 41.05 77.166 41.15 ;
      RECT MASK 2 77.454 41.05 83.784 41.15 ;
      RECT MASK 2 84.072 41.05 90.402 41.15 ;
      RECT MASK 2 90.69 41.05 97.02 41.15 ;
      RECT MASK 2 97.308 41.05 103.638 41.15 ;
      RECT MASK 2 103.926 41.05 110.256 41.15 ;
      RECT MASK 2 4.672 41.425 10.96 41.525 ;
      RECT MASK 2 11.29 41.425 17.578 41.525 ;
      RECT MASK 2 17.908 41.425 24.196 41.525 ;
      RECT MASK 2 24.526 41.425 30.814 41.525 ;
      RECT MASK 2 31.144 41.425 37.432 41.525 ;
      RECT MASK 2 37.762 41.425 44.05 41.525 ;
      RECT MASK 2 44.38 41.425 50.668 41.525 ;
      RECT MASK 2 50.998 41.425 57.286 41.525 ;
      RECT MASK 2 57.616 41.425 63.904 41.525 ;
      RECT MASK 2 64.234 41.425 70.522 41.525 ;
      RECT MASK 2 70.852 41.425 77.14 41.525 ;
      RECT MASK 2 77.47 41.425 83.758 41.525 ;
      RECT MASK 2 84.088 41.425 90.376 41.525 ;
      RECT MASK 2 90.706 41.425 96.994 41.525 ;
      RECT MASK 2 97.324 41.425 103.612 41.525 ;
      RECT MASK 2 103.942 41.425 110.23 41.525 ;
      RECT MASK 2 111.044 41.4575 129.1315 41.5575 ;
      RECT MASK 2 111.044 41.7775 129.1315 42.0275 ;
      RECT MASK 2 4.672 41.795 10.96 41.895 ;
      RECT MASK 2 11.29 41.795 17.578 41.895 ;
      RECT MASK 2 17.908 41.795 24.196 41.895 ;
      RECT MASK 2 24.526 41.795 30.814 41.895 ;
      RECT MASK 2 31.144 41.795 37.432 41.895 ;
      RECT MASK 2 37.762 41.795 44.05 41.895 ;
      RECT MASK 2 44.38 41.795 50.668 41.895 ;
      RECT MASK 2 50.998 41.795 57.286 41.895 ;
      RECT MASK 2 57.616 41.795 63.904 41.895 ;
      RECT MASK 2 64.234 41.795 70.522 41.895 ;
      RECT MASK 2 70.852 41.795 77.14 41.895 ;
      RECT MASK 2 77.47 41.795 83.758 41.895 ;
      RECT MASK 2 84.088 41.795 90.376 41.895 ;
      RECT MASK 2 90.706 41.795 96.994 41.895 ;
      RECT MASK 2 97.324 41.795 103.612 41.895 ;
      RECT MASK 2 103.942 41.795 110.23 41.895 ;
      RECT MASK 2 4.656 42.17 10.986 42.27 ;
      RECT MASK 2 11.274 42.17 17.604 42.27 ;
      RECT MASK 2 17.892 42.17 24.222 42.27 ;
      RECT MASK 2 24.51 42.17 30.84 42.27 ;
      RECT MASK 2 31.128 42.17 37.458 42.27 ;
      RECT MASK 2 37.746 42.17 44.076 42.27 ;
      RECT MASK 2 44.364 42.17 50.694 42.27 ;
      RECT MASK 2 50.982 42.17 57.312 42.27 ;
      RECT MASK 2 57.6 42.17 63.93 42.27 ;
      RECT MASK 2 64.218 42.17 70.548 42.27 ;
      RECT MASK 2 70.836 42.17 77.166 42.27 ;
      RECT MASK 2 77.454 42.17 83.784 42.27 ;
      RECT MASK 2 84.072 42.17 90.402 42.27 ;
      RECT MASK 2 90.69 42.17 97.02 42.27 ;
      RECT MASK 2 97.308 42.17 103.638 42.27 ;
      RECT MASK 2 103.926 42.17 110.256 42.27 ;
      RECT MASK 2 111.044 42.2925 127.58 42.3925 ;
      RECT MASK 2 4.672 42.545 10.96 42.645 ;
      RECT MASK 2 11.29 42.545 17.578 42.645 ;
      RECT MASK 2 17.908 42.545 24.196 42.645 ;
      RECT MASK 2 24.526 42.545 30.814 42.645 ;
      RECT MASK 2 31.144 42.545 37.432 42.645 ;
      RECT MASK 2 37.762 42.545 44.05 42.645 ;
      RECT MASK 2 44.38 42.545 50.668 42.645 ;
      RECT MASK 2 50.998 42.545 57.286 42.645 ;
      RECT MASK 2 57.616 42.545 63.904 42.645 ;
      RECT MASK 2 64.234 42.545 70.522 42.645 ;
      RECT MASK 2 70.852 42.545 77.14 42.645 ;
      RECT MASK 2 77.47 42.545 83.758 42.645 ;
      RECT MASK 2 84.088 42.545 90.376 42.645 ;
      RECT MASK 2 90.706 42.545 96.994 42.645 ;
      RECT MASK 2 97.324 42.545 103.612 42.645 ;
      RECT MASK 2 103.942 42.545 110.23 42.645 ;
      RECT MASK 2 111.044 42.8075 127.58 42.9075 ;
      RECT MASK 2 4.672 42.915 10.96 43.015 ;
      RECT MASK 2 11.29 42.915 17.578 43.015 ;
      RECT MASK 2 17.908 42.915 24.196 43.015 ;
      RECT MASK 2 24.526 42.915 30.814 43.015 ;
      RECT MASK 2 31.144 42.915 37.432 43.015 ;
      RECT MASK 2 37.762 42.915 44.05 43.015 ;
      RECT MASK 2 44.38 42.915 50.668 43.015 ;
      RECT MASK 2 50.998 42.915 57.286 43.015 ;
      RECT MASK 2 57.616 42.915 63.904 43.015 ;
      RECT MASK 2 64.234 42.915 70.522 43.015 ;
      RECT MASK 2 70.852 42.915 77.14 43.015 ;
      RECT MASK 2 77.47 42.915 83.758 43.015 ;
      RECT MASK 2 84.088 42.915 90.376 43.015 ;
      RECT MASK 2 90.706 42.915 96.994 43.015 ;
      RECT MASK 2 97.324 42.915 103.612 43.015 ;
      RECT MASK 2 103.942 42.915 110.23 43.015 ;
      RECT MASK 2 111.044 43.1275 129.1315 43.3775 ;
      RECT MASK 2 4.656 43.29 10.986 43.39 ;
      RECT MASK 2 11.274 43.29 17.604 43.39 ;
      RECT MASK 2 17.892 43.29 24.222 43.39 ;
      RECT MASK 2 24.51 43.29 30.84 43.39 ;
      RECT MASK 2 31.128 43.29 37.458 43.39 ;
      RECT MASK 2 37.746 43.29 44.076 43.39 ;
      RECT MASK 2 44.364 43.29 50.694 43.39 ;
      RECT MASK 2 50.982 43.29 57.312 43.39 ;
      RECT MASK 2 57.6 43.29 63.93 43.39 ;
      RECT MASK 2 64.218 43.29 70.548 43.39 ;
      RECT MASK 2 70.836 43.29 77.166 43.39 ;
      RECT MASK 2 77.454 43.29 83.784 43.39 ;
      RECT MASK 2 84.072 43.29 90.402 43.39 ;
      RECT MASK 2 90.69 43.29 97.02 43.39 ;
      RECT MASK 2 97.308 43.29 103.638 43.39 ;
      RECT MASK 2 103.926 43.29 110.256 43.39 ;
      RECT MASK 2 111.044 43.6425 127.58 43.7425 ;
      RECT MASK 2 4.672 43.665 10.96 43.765 ;
      RECT MASK 2 11.29 43.665 17.578 43.765 ;
      RECT MASK 2 17.908 43.665 24.196 43.765 ;
      RECT MASK 2 24.526 43.665 30.814 43.765 ;
      RECT MASK 2 31.144 43.665 37.432 43.765 ;
      RECT MASK 2 37.762 43.665 44.05 43.765 ;
      RECT MASK 2 44.38 43.665 50.668 43.765 ;
      RECT MASK 2 50.998 43.665 57.286 43.765 ;
      RECT MASK 2 57.616 43.665 63.904 43.765 ;
      RECT MASK 2 64.234 43.665 70.522 43.765 ;
      RECT MASK 2 70.852 43.665 77.14 43.765 ;
      RECT MASK 2 77.47 43.665 83.758 43.765 ;
      RECT MASK 2 84.088 43.665 90.376 43.765 ;
      RECT MASK 2 90.706 43.665 96.994 43.765 ;
      RECT MASK 2 97.324 43.665 103.612 43.765 ;
      RECT MASK 2 103.942 43.665 110.23 43.765 ;
      RECT MASK 2 4.672 44.035 10.96 44.135 ;
      RECT MASK 2 11.29 44.035 17.578 44.135 ;
      RECT MASK 2 17.908 44.035 24.196 44.135 ;
      RECT MASK 2 24.526 44.035 30.814 44.135 ;
      RECT MASK 2 31.144 44.035 37.432 44.135 ;
      RECT MASK 2 37.762 44.035 44.05 44.135 ;
      RECT MASK 2 44.38 44.035 50.668 44.135 ;
      RECT MASK 2 50.998 44.035 57.286 44.135 ;
      RECT MASK 2 57.616 44.035 63.904 44.135 ;
      RECT MASK 2 64.234 44.035 70.522 44.135 ;
      RECT MASK 2 70.852 44.035 77.14 44.135 ;
      RECT MASK 2 77.47 44.035 83.758 44.135 ;
      RECT MASK 2 84.088 44.035 90.376 44.135 ;
      RECT MASK 2 90.706 44.035 96.994 44.135 ;
      RECT MASK 2 97.324 44.035 103.612 44.135 ;
      RECT MASK 2 103.942 44.035 110.23 44.135 ;
      RECT MASK 2 111.044 44.1575 127.58 44.2575 ;
      RECT MASK 2 4.656 44.41 10.986 44.51 ;
      RECT MASK 2 11.274 44.41 17.604 44.51 ;
      RECT MASK 2 17.892 44.41 24.222 44.51 ;
      RECT MASK 2 24.51 44.41 30.84 44.51 ;
      RECT MASK 2 31.128 44.41 37.458 44.51 ;
      RECT MASK 2 37.746 44.41 44.076 44.51 ;
      RECT MASK 2 44.364 44.41 50.694 44.51 ;
      RECT MASK 2 50.982 44.41 57.312 44.51 ;
      RECT MASK 2 57.6 44.41 63.93 44.51 ;
      RECT MASK 2 64.218 44.41 70.548 44.51 ;
      RECT MASK 2 70.836 44.41 77.166 44.51 ;
      RECT MASK 2 77.454 44.41 83.784 44.51 ;
      RECT MASK 2 84.072 44.41 90.402 44.51 ;
      RECT MASK 2 90.69 44.41 97.02 44.51 ;
      RECT MASK 2 97.308 44.41 103.638 44.51 ;
      RECT MASK 2 103.926 44.41 110.256 44.51 ;
      RECT MASK 2 111.044 44.4775 129.1315 44.7275 ;
      RECT MASK 2 4.672 44.785 10.96 44.885 ;
      RECT MASK 2 11.29 44.785 17.578 44.885 ;
      RECT MASK 2 17.908 44.785 24.196 44.885 ;
      RECT MASK 2 24.526 44.785 30.814 44.885 ;
      RECT MASK 2 31.144 44.785 37.432 44.885 ;
      RECT MASK 2 37.762 44.785 44.05 44.885 ;
      RECT MASK 2 44.38 44.785 50.668 44.885 ;
      RECT MASK 2 50.998 44.785 57.286 44.885 ;
      RECT MASK 2 57.616 44.785 63.904 44.885 ;
      RECT MASK 2 64.234 44.785 70.522 44.885 ;
      RECT MASK 2 70.852 44.785 77.14 44.885 ;
      RECT MASK 2 77.47 44.785 83.758 44.885 ;
      RECT MASK 2 84.088 44.785 90.376 44.885 ;
      RECT MASK 2 90.706 44.785 96.994 44.885 ;
      RECT MASK 2 97.324 44.785 103.612 44.885 ;
      RECT MASK 2 103.942 44.785 110.23 44.885 ;
      RECT MASK 2 111.044 44.9475 127.58 45.0475 ;
      RECT MASK 2 0.567 45.54 115.126 45.66 ;
      RECT MASK 2 117.268 45.555 129.1315 45.615 ;
      RECT MASK 2 117.181 45.859 129.1315 45.899 ;
      RECT MASK 2 0.567 45.96 115.126 46.08 ;
      RECT MASK 2 117.181 46.019 129.1315 46.059 ;
      RECT MASK 2 117.181 46.179 129.1315 46.219 ;
      RECT MASK 2 117.181 46.339 129.1315 46.379 ;
      RECT MASK 2 4.672 46.795 10.96 46.895 ;
      RECT MASK 2 11.29 46.795 24.196 46.895 ;
      RECT MASK 2 24.526 46.795 37.432 46.895 ;
      RECT MASK 2 37.762 46.795 50.668 46.895 ;
      RECT MASK 2 50.998 46.795 63.904 46.895 ;
      RECT MASK 2 64.234 46.795 77.14 46.895 ;
      RECT MASK 2 77.47 46.795 90.376 46.895 ;
      RECT MASK 2 90.706 46.795 103.612 46.895 ;
      RECT MASK 2 103.942 46.795 126.291 46.895 ;
      RECT MASK 2 4.656 47.17 10.986 47.27 ;
      RECT MASK 2 11.274 47.17 24.222 47.27 ;
      RECT MASK 2 24.51 47.17 37.458 47.27 ;
      RECT MASK 2 37.746 47.17 50.694 47.27 ;
      RECT MASK 2 50.982 47.17 63.93 47.27 ;
      RECT MASK 2 64.218 47.17 77.166 47.27 ;
      RECT MASK 2 77.454 47.17 90.402 47.27 ;
      RECT MASK 2 90.69 47.17 103.638 47.27 ;
      RECT MASK 2 103.926 47.17 126.291 47.27 ;
      RECT MASK 2 4.672 47.545 10.96 47.645 ;
      RECT MASK 2 11.29 47.545 24.196 47.645 ;
      RECT MASK 2 24.526 47.545 37.432 47.645 ;
      RECT MASK 2 37.762 47.545 50.668 47.645 ;
      RECT MASK 2 50.998 47.545 63.904 47.645 ;
      RECT MASK 2 64.234 47.545 77.14 47.645 ;
      RECT MASK 2 77.47 47.545 90.376 47.645 ;
      RECT MASK 2 90.706 47.545 103.612 47.645 ;
      RECT MASK 2 103.942 47.545 126.291 47.645 ;
      RECT MASK 2 4.672 47.915 10.96 48.015 ;
      RECT MASK 2 11.29 47.915 24.196 48.015 ;
      RECT MASK 2 24.526 47.915 37.432 48.015 ;
      RECT MASK 2 37.762 47.915 50.668 48.015 ;
      RECT MASK 2 50.998 47.915 63.904 48.015 ;
      RECT MASK 2 64.234 47.915 77.14 48.015 ;
      RECT MASK 2 77.47 47.915 90.376 48.015 ;
      RECT MASK 2 90.706 47.915 103.612 48.015 ;
      RECT MASK 2 103.942 47.915 126.291 48.015 ;
      RECT MASK 2 4.656 48.29 10.986 48.39 ;
      RECT MASK 2 11.274 48.29 24.222 48.39 ;
      RECT MASK 2 24.51 48.29 37.458 48.39 ;
      RECT MASK 2 37.746 48.29 50.694 48.39 ;
      RECT MASK 2 50.982 48.29 63.93 48.39 ;
      RECT MASK 2 64.218 48.29 77.166 48.39 ;
      RECT MASK 2 77.454 48.29 90.402 48.39 ;
      RECT MASK 2 90.69 48.29 103.638 48.39 ;
      RECT MASK 2 103.926 48.29 126.291 48.39 ;
      RECT MASK 2 4.672 48.665 10.96 48.765 ;
      RECT MASK 2 11.29 48.665 24.196 48.765 ;
      RECT MASK 2 24.526 48.665 37.432 48.765 ;
      RECT MASK 2 37.762 48.665 50.668 48.765 ;
      RECT MASK 2 50.998 48.665 63.904 48.765 ;
      RECT MASK 2 64.234 48.665 77.14 48.765 ;
      RECT MASK 2 77.47 48.665 90.376 48.765 ;
      RECT MASK 2 90.706 48.665 103.612 48.765 ;
      RECT MASK 2 103.942 48.665 126.291 48.765 ;
      RECT MASK 2 4.672 49.035 10.96 49.135 ;
      RECT MASK 2 11.29 49.035 24.196 49.135 ;
      RECT MASK 2 24.526 49.035 37.432 49.135 ;
      RECT MASK 2 37.762 49.035 50.668 49.135 ;
      RECT MASK 2 50.998 49.035 63.904 49.135 ;
      RECT MASK 2 64.234 49.035 77.14 49.135 ;
      RECT MASK 2 77.47 49.035 90.376 49.135 ;
      RECT MASK 2 90.706 49.035 103.612 49.135 ;
      RECT MASK 2 103.942 49.035 126.291 49.135 ;
      RECT MASK 2 4.656 49.41 10.986 49.51 ;
      RECT MASK 2 11.274 49.41 24.222 49.51 ;
      RECT MASK 2 24.51 49.41 37.458 49.51 ;
      RECT MASK 2 37.746 49.41 50.694 49.51 ;
      RECT MASK 2 50.982 49.41 63.93 49.51 ;
      RECT MASK 2 64.218 49.41 77.166 49.51 ;
      RECT MASK 2 77.454 49.41 90.402 49.51 ;
      RECT MASK 2 90.69 49.41 103.638 49.51 ;
      RECT MASK 2 103.926 49.41 126.291 49.51 ;
      RECT MASK 2 4.672 49.785 10.96 49.885 ;
      RECT MASK 2 11.29 49.785 24.196 49.885 ;
      RECT MASK 2 24.526 49.785 37.432 49.885 ;
      RECT MASK 2 37.762 49.785 50.668 49.885 ;
      RECT MASK 2 50.998 49.785 63.904 49.885 ;
      RECT MASK 2 64.234 49.785 77.14 49.885 ;
      RECT MASK 2 77.47 49.785 90.376 49.885 ;
      RECT MASK 2 90.706 49.785 103.612 49.885 ;
      RECT MASK 2 103.942 49.785 126.291 49.885 ;
      RECT MASK 2 4.672 50.155 10.96 50.255 ;
      RECT MASK 2 11.29 50.155 24.196 50.255 ;
      RECT MASK 2 24.526 50.155 37.432 50.255 ;
      RECT MASK 2 37.762 50.155 50.668 50.255 ;
      RECT MASK 2 50.998 50.155 63.904 50.255 ;
      RECT MASK 2 64.234 50.155 77.14 50.255 ;
      RECT MASK 2 77.47 50.155 90.376 50.255 ;
      RECT MASK 2 90.706 50.155 103.612 50.255 ;
      RECT MASK 2 103.942 50.155 126.291 50.255 ;
      RECT MASK 2 4.656 50.53 10.986 50.63 ;
      RECT MASK 2 11.274 50.53 24.222 50.63 ;
      RECT MASK 2 24.51 50.53 37.458 50.63 ;
      RECT MASK 2 37.746 50.53 50.694 50.63 ;
      RECT MASK 2 50.982 50.53 63.93 50.63 ;
      RECT MASK 2 64.218 50.53 77.166 50.63 ;
      RECT MASK 2 77.454 50.53 90.402 50.63 ;
      RECT MASK 2 90.69 50.53 103.638 50.63 ;
      RECT MASK 2 103.926 50.53 126.291 50.63 ;
      RECT MASK 2 4.672 50.905 10.96 51.005 ;
      RECT MASK 2 11.29 50.905 24.196 51.005 ;
      RECT MASK 2 24.526 50.905 37.432 51.005 ;
      RECT MASK 2 37.762 50.905 50.668 51.005 ;
      RECT MASK 2 50.998 50.905 63.904 51.005 ;
      RECT MASK 2 64.234 50.905 77.14 51.005 ;
      RECT MASK 2 77.47 50.905 90.376 51.005 ;
      RECT MASK 2 90.706 50.905 103.612 51.005 ;
      RECT MASK 2 103.942 50.905 126.291 51.005 ;
      RECT MASK 2 117.181 51.42 129.1315 51.46 ;
      RECT MASK 2 117.181 51.58 129.1315 51.62 ;
      RECT MASK 2 0.567 51.66 115.126 51.78 ;
      RECT MASK 2 117.181 51.74 129.1315 51.78 ;
      RECT MASK 2 117.181 51.9 129.1315 51.94 ;
      RECT MASK 2 117.181 52.06 129.1315 52.1 ;
      RECT MASK 2 0.567 52.08 115.126 52.2 ;
      RECT MASK 2 117.181 52.22 129.1315 52.26 ;
      RECT MASK 2 117.181 52.38 129.1315 52.42 ;
      RECT MASK 2 4.672 52.915 10.96 53.015 ;
      RECT MASK 2 11.29 52.915 24.196 53.015 ;
      RECT MASK 2 24.526 52.915 37.432 53.015 ;
      RECT MASK 2 37.762 52.915 50.668 53.015 ;
      RECT MASK 2 50.998 52.915 63.904 53.015 ;
      RECT MASK 2 64.234 52.915 77.14 53.015 ;
      RECT MASK 2 77.47 52.915 90.376 53.015 ;
      RECT MASK 2 90.706 52.915 103.612 53.015 ;
      RECT MASK 2 103.942 52.915 126.291 53.015 ;
      RECT MASK 2 4.656 53.29 10.986 53.39 ;
      RECT MASK 2 11.274 53.29 24.222 53.39 ;
      RECT MASK 2 24.51 53.29 37.458 53.39 ;
      RECT MASK 2 37.746 53.29 50.694 53.39 ;
      RECT MASK 2 50.982 53.29 63.93 53.39 ;
      RECT MASK 2 64.218 53.29 77.166 53.39 ;
      RECT MASK 2 77.454 53.29 90.402 53.39 ;
      RECT MASK 2 90.69 53.29 103.638 53.39 ;
      RECT MASK 2 103.926 53.29 126.291 53.39 ;
      RECT MASK 2 4.672 53.665 10.96 53.765 ;
      RECT MASK 2 11.29 53.665 24.196 53.765 ;
      RECT MASK 2 24.526 53.665 37.432 53.765 ;
      RECT MASK 2 37.762 53.665 50.668 53.765 ;
      RECT MASK 2 50.998 53.665 63.904 53.765 ;
      RECT MASK 2 64.234 53.665 77.14 53.765 ;
      RECT MASK 2 77.47 53.665 90.376 53.765 ;
      RECT MASK 2 90.706 53.665 103.612 53.765 ;
      RECT MASK 2 103.942 53.665 126.291 53.765 ;
      RECT MASK 2 4.672 54.035 10.96 54.135 ;
      RECT MASK 2 11.29 54.035 24.196 54.135 ;
      RECT MASK 2 24.526 54.035 37.432 54.135 ;
      RECT MASK 2 37.762 54.035 50.668 54.135 ;
      RECT MASK 2 50.998 54.035 63.904 54.135 ;
      RECT MASK 2 64.234 54.035 77.14 54.135 ;
      RECT MASK 2 77.47 54.035 90.376 54.135 ;
      RECT MASK 2 90.706 54.035 103.612 54.135 ;
      RECT MASK 2 103.942 54.035 126.291 54.135 ;
      RECT MASK 2 4.656 54.41 10.986 54.51 ;
      RECT MASK 2 11.274 54.41 24.222 54.51 ;
      RECT MASK 2 24.51 54.41 37.458 54.51 ;
      RECT MASK 2 37.746 54.41 50.694 54.51 ;
      RECT MASK 2 50.982 54.41 63.93 54.51 ;
      RECT MASK 2 64.218 54.41 77.166 54.51 ;
      RECT MASK 2 77.454 54.41 90.402 54.51 ;
      RECT MASK 2 90.69 54.41 103.638 54.51 ;
      RECT MASK 2 103.926 54.41 126.291 54.51 ;
      RECT MASK 2 4.672 54.785 10.96 54.885 ;
      RECT MASK 2 11.29 54.785 24.196 54.885 ;
      RECT MASK 2 24.526 54.785 37.432 54.885 ;
      RECT MASK 2 37.762 54.785 50.668 54.885 ;
      RECT MASK 2 50.998 54.785 63.904 54.885 ;
      RECT MASK 2 64.234 54.785 77.14 54.885 ;
      RECT MASK 2 77.47 54.785 90.376 54.885 ;
      RECT MASK 2 90.706 54.785 103.612 54.885 ;
      RECT MASK 2 103.942 54.785 126.291 54.885 ;
      RECT MASK 2 4.672 55.155 10.96 55.255 ;
      RECT MASK 2 11.29 55.155 24.196 55.255 ;
      RECT MASK 2 24.526 55.155 37.432 55.255 ;
      RECT MASK 2 37.762 55.155 50.668 55.255 ;
      RECT MASK 2 50.998 55.155 63.904 55.255 ;
      RECT MASK 2 64.234 55.155 77.14 55.255 ;
      RECT MASK 2 77.47 55.155 90.376 55.255 ;
      RECT MASK 2 90.706 55.155 103.612 55.255 ;
      RECT MASK 2 103.942 55.155 126.291 55.255 ;
      RECT MASK 2 4.656 55.53 10.986 55.63 ;
      RECT MASK 2 11.274 55.53 24.222 55.63 ;
      RECT MASK 2 24.51 55.53 37.458 55.63 ;
      RECT MASK 2 37.746 55.53 50.694 55.63 ;
      RECT MASK 2 50.982 55.53 63.93 55.63 ;
      RECT MASK 2 64.218 55.53 77.166 55.63 ;
      RECT MASK 2 77.454 55.53 90.402 55.63 ;
      RECT MASK 2 90.69 55.53 103.638 55.63 ;
      RECT MASK 2 103.926 55.53 126.291 55.63 ;
      RECT MASK 2 4.672 55.905 10.96 56.005 ;
      RECT MASK 2 11.29 55.905 24.196 56.005 ;
      RECT MASK 2 24.526 55.905 37.432 56.005 ;
      RECT MASK 2 37.762 55.905 50.668 56.005 ;
      RECT MASK 2 50.998 55.905 63.904 56.005 ;
      RECT MASK 2 64.234 55.905 77.14 56.005 ;
      RECT MASK 2 77.47 55.905 90.376 56.005 ;
      RECT MASK 2 90.706 55.905 103.612 56.005 ;
      RECT MASK 2 103.942 55.905 126.291 56.005 ;
      RECT MASK 2 4.672 56.275 10.96 56.375 ;
      RECT MASK 2 11.29 56.275 24.196 56.375 ;
      RECT MASK 2 24.526 56.275 37.432 56.375 ;
      RECT MASK 2 37.762 56.275 50.668 56.375 ;
      RECT MASK 2 50.998 56.275 63.904 56.375 ;
      RECT MASK 2 64.234 56.275 77.14 56.375 ;
      RECT MASK 2 77.47 56.275 90.376 56.375 ;
      RECT MASK 2 90.706 56.275 103.612 56.375 ;
      RECT MASK 2 103.942 56.275 126.291 56.375 ;
      RECT MASK 2 4.656 56.65 10.986 56.75 ;
      RECT MASK 2 11.274 56.65 24.222 56.75 ;
      RECT MASK 2 24.51 56.65 37.458 56.75 ;
      RECT MASK 2 37.746 56.65 50.694 56.75 ;
      RECT MASK 2 50.982 56.65 63.93 56.75 ;
      RECT MASK 2 64.218 56.65 77.166 56.75 ;
      RECT MASK 2 77.454 56.65 90.402 56.75 ;
      RECT MASK 2 90.69 56.65 103.638 56.75 ;
      RECT MASK 2 103.926 56.65 126.291 56.75 ;
      RECT MASK 2 4.672 57.025 10.96 57.125 ;
      RECT MASK 2 11.29 57.025 24.196 57.125 ;
      RECT MASK 2 24.526 57.025 37.432 57.125 ;
      RECT MASK 2 37.762 57.025 50.668 57.125 ;
      RECT MASK 2 50.998 57.025 63.904 57.125 ;
      RECT MASK 2 64.234 57.025 77.14 57.125 ;
      RECT MASK 2 77.47 57.025 90.376 57.125 ;
      RECT MASK 2 90.706 57.025 103.612 57.125 ;
      RECT MASK 2 103.942 57.025 126.291 57.125 ;
      RECT MASK 2 117.181 57.63 129.1315 57.67 ;
      RECT MASK 2 0.567 57.78 115.126 57.9 ;
      RECT MASK 2 117.181 57.79 129.1315 57.83 ;
      RECT MASK 2 117.181 57.95 129.1315 57.99 ;
      RECT MASK 2 0.567 58.2 115.126 58.32 ;
      RECT MASK 2 111.044 58.9075 129.1315 59.1575 ;
      RECT MASK 2 4.672 59.035 10.96 59.135 ;
      RECT MASK 2 11.29 59.035 17.578 59.135 ;
      RECT MASK 2 17.908 59.035 24.196 59.135 ;
      RECT MASK 2 24.526 59.035 30.814 59.135 ;
      RECT MASK 2 31.144 59.035 37.432 59.135 ;
      RECT MASK 2 37.762 59.035 44.05 59.135 ;
      RECT MASK 2 44.38 59.035 50.668 59.135 ;
      RECT MASK 2 50.998 59.035 57.286 59.135 ;
      RECT MASK 2 57.616 59.035 63.904 59.135 ;
      RECT MASK 2 64.234 59.035 70.522 59.135 ;
      RECT MASK 2 70.852 59.035 77.14 59.135 ;
      RECT MASK 2 77.47 59.035 83.758 59.135 ;
      RECT MASK 2 84.088 59.035 90.376 59.135 ;
      RECT MASK 2 90.706 59.035 96.994 59.135 ;
      RECT MASK 2 97.324 59.035 103.612 59.135 ;
      RECT MASK 2 103.942 59.035 110.23 59.135 ;
      RECT MASK 2 4.656 59.41 10.986 59.51 ;
      RECT MASK 2 11.274 59.41 17.604 59.51 ;
      RECT MASK 2 17.892 59.41 24.222 59.51 ;
      RECT MASK 2 24.51 59.41 30.84 59.51 ;
      RECT MASK 2 31.128 59.41 37.458 59.51 ;
      RECT MASK 2 37.746 59.41 44.076 59.51 ;
      RECT MASK 2 44.364 59.41 50.694 59.51 ;
      RECT MASK 2 50.982 59.41 57.312 59.51 ;
      RECT MASK 2 57.6 59.41 63.93 59.51 ;
      RECT MASK 2 64.218 59.41 70.548 59.51 ;
      RECT MASK 2 70.836 59.41 77.166 59.51 ;
      RECT MASK 2 77.454 59.41 83.784 59.51 ;
      RECT MASK 2 84.072 59.41 90.402 59.51 ;
      RECT MASK 2 90.69 59.41 97.02 59.51 ;
      RECT MASK 2 97.308 59.41 103.638 59.51 ;
      RECT MASK 2 103.926 59.41 110.256 59.51 ;
      RECT MASK 2 111.044 59.4225 129.1315 59.5225 ;
      RECT MASK 2 4.672 59.785 10.96 59.885 ;
      RECT MASK 2 11.29 59.785 17.578 59.885 ;
      RECT MASK 2 17.908 59.785 24.196 59.885 ;
      RECT MASK 2 24.526 59.785 30.814 59.885 ;
      RECT MASK 2 31.144 59.785 37.432 59.885 ;
      RECT MASK 2 37.762 59.785 44.05 59.885 ;
      RECT MASK 2 44.38 59.785 50.668 59.885 ;
      RECT MASK 2 50.998 59.785 57.286 59.885 ;
      RECT MASK 2 57.616 59.785 63.904 59.885 ;
      RECT MASK 2 64.234 59.785 70.522 59.885 ;
      RECT MASK 2 70.852 59.785 77.14 59.885 ;
      RECT MASK 2 77.47 59.785 83.758 59.885 ;
      RECT MASK 2 84.088 59.785 90.376 59.885 ;
      RECT MASK 2 90.706 59.785 96.994 59.885 ;
      RECT MASK 2 97.324 59.785 103.612 59.885 ;
      RECT MASK 2 103.942 59.785 110.23 59.885 ;
      RECT MASK 2 111.044 59.9375 127.58 60.0375 ;
      RECT MASK 2 4.672 60.155 10.96 60.255 ;
      RECT MASK 2 11.29 60.155 17.578 60.255 ;
      RECT MASK 2 17.908 60.155 24.196 60.255 ;
      RECT MASK 2 24.526 60.155 30.814 60.255 ;
      RECT MASK 2 31.144 60.155 37.432 60.255 ;
      RECT MASK 2 37.762 60.155 44.05 60.255 ;
      RECT MASK 2 44.38 60.155 50.668 60.255 ;
      RECT MASK 2 50.998 60.155 57.286 60.255 ;
      RECT MASK 2 57.616 60.155 63.904 60.255 ;
      RECT MASK 2 64.234 60.155 70.522 60.255 ;
      RECT MASK 2 70.852 60.155 77.14 60.255 ;
      RECT MASK 2 77.47 60.155 83.758 60.255 ;
      RECT MASK 2 84.088 60.155 90.376 60.255 ;
      RECT MASK 2 90.706 60.155 96.994 60.255 ;
      RECT MASK 2 97.324 60.155 103.612 60.255 ;
      RECT MASK 2 103.942 60.155 110.23 60.255 ;
      RECT MASK 2 111.044 60.2575 129.1315 60.5075 ;
      RECT MASK 2 4.656 60.53 10.986 60.63 ;
      RECT MASK 2 11.274 60.53 17.604 60.63 ;
      RECT MASK 2 17.892 60.53 24.222 60.63 ;
      RECT MASK 2 24.51 60.53 30.84 60.63 ;
      RECT MASK 2 31.128 60.53 37.458 60.63 ;
      RECT MASK 2 37.746 60.53 44.076 60.63 ;
      RECT MASK 2 44.364 60.53 50.694 60.63 ;
      RECT MASK 2 50.982 60.53 57.312 60.63 ;
      RECT MASK 2 57.6 60.53 63.93 60.63 ;
      RECT MASK 2 64.218 60.53 70.548 60.63 ;
      RECT MASK 2 70.836 60.53 77.166 60.63 ;
      RECT MASK 2 77.454 60.53 83.784 60.63 ;
      RECT MASK 2 84.072 60.53 90.402 60.63 ;
      RECT MASK 2 90.69 60.53 97.02 60.63 ;
      RECT MASK 2 97.308 60.53 103.638 60.63 ;
      RECT MASK 2 103.926 60.53 110.256 60.63 ;
      RECT MASK 2 111.044 60.7725 129.1315 60.8725 ;
      RECT MASK 2 4.672 60.905 10.96 61.005 ;
      RECT MASK 2 11.29 60.905 17.578 61.005 ;
      RECT MASK 2 17.908 60.905 24.196 61.005 ;
      RECT MASK 2 24.526 60.905 30.814 61.005 ;
      RECT MASK 2 31.144 60.905 37.432 61.005 ;
      RECT MASK 2 37.762 60.905 44.05 61.005 ;
      RECT MASK 2 44.38 60.905 50.668 61.005 ;
      RECT MASK 2 50.998 60.905 57.286 61.005 ;
      RECT MASK 2 57.616 60.905 63.904 61.005 ;
      RECT MASK 2 64.234 60.905 70.522 61.005 ;
      RECT MASK 2 70.852 60.905 77.14 61.005 ;
      RECT MASK 2 77.47 60.905 83.758 61.005 ;
      RECT MASK 2 84.088 60.905 90.376 61.005 ;
      RECT MASK 2 90.706 60.905 96.994 61.005 ;
      RECT MASK 2 97.324 60.905 103.612 61.005 ;
      RECT MASK 2 103.942 60.905 110.23 61.005 ;
      RECT MASK 2 4.672 61.275 10.96 61.375 ;
      RECT MASK 2 11.29 61.275 17.578 61.375 ;
      RECT MASK 2 17.908 61.275 24.196 61.375 ;
      RECT MASK 2 24.526 61.275 30.814 61.375 ;
      RECT MASK 2 31.144 61.275 37.432 61.375 ;
      RECT MASK 2 37.762 61.275 44.05 61.375 ;
      RECT MASK 2 44.38 61.275 50.668 61.375 ;
      RECT MASK 2 50.998 61.275 57.286 61.375 ;
      RECT MASK 2 57.616 61.275 63.904 61.375 ;
      RECT MASK 2 64.234 61.275 70.522 61.375 ;
      RECT MASK 2 70.852 61.275 77.14 61.375 ;
      RECT MASK 2 77.47 61.275 83.758 61.375 ;
      RECT MASK 2 84.088 61.275 90.376 61.375 ;
      RECT MASK 2 90.706 61.275 96.994 61.375 ;
      RECT MASK 2 97.324 61.275 103.612 61.375 ;
      RECT MASK 2 103.942 61.275 110.23 61.375 ;
      RECT MASK 2 111.044 61.2875 127.58 61.3875 ;
      RECT MASK 2 111.044 61.6075 129.1315 61.8575 ;
      RECT MASK 2 4.656 61.65 10.986 61.75 ;
      RECT MASK 2 11.274 61.65 17.604 61.75 ;
      RECT MASK 2 17.892 61.65 24.222 61.75 ;
      RECT MASK 2 24.51 61.65 30.84 61.75 ;
      RECT MASK 2 31.128 61.65 37.458 61.75 ;
      RECT MASK 2 37.746 61.65 44.076 61.75 ;
      RECT MASK 2 44.364 61.65 50.694 61.75 ;
      RECT MASK 2 50.982 61.65 57.312 61.75 ;
      RECT MASK 2 57.6 61.65 63.93 61.75 ;
      RECT MASK 2 64.218 61.65 70.548 61.75 ;
      RECT MASK 2 70.836 61.65 77.166 61.75 ;
      RECT MASK 2 77.454 61.65 83.784 61.75 ;
      RECT MASK 2 84.072 61.65 90.402 61.75 ;
      RECT MASK 2 90.69 61.65 97.02 61.75 ;
      RECT MASK 2 97.308 61.65 103.638 61.75 ;
      RECT MASK 2 103.926 61.65 110.256 61.75 ;
      RECT MASK 2 4.672 62.025 10.96 62.125 ;
      RECT MASK 2 11.29 62.025 17.578 62.125 ;
      RECT MASK 2 17.908 62.025 24.196 62.125 ;
      RECT MASK 2 24.526 62.025 30.814 62.125 ;
      RECT MASK 2 31.144 62.025 37.432 62.125 ;
      RECT MASK 2 37.762 62.025 44.05 62.125 ;
      RECT MASK 2 44.38 62.025 50.668 62.125 ;
      RECT MASK 2 50.998 62.025 57.286 62.125 ;
      RECT MASK 2 57.616 62.025 63.904 62.125 ;
      RECT MASK 2 64.234 62.025 70.522 62.125 ;
      RECT MASK 2 70.852 62.025 77.14 62.125 ;
      RECT MASK 2 77.47 62.025 83.758 62.125 ;
      RECT MASK 2 84.088 62.025 90.376 62.125 ;
      RECT MASK 2 90.706 62.025 96.994 62.125 ;
      RECT MASK 2 97.324 62.025 103.612 62.125 ;
      RECT MASK 2 103.942 62.025 110.23 62.125 ;
      RECT MASK 2 111.044 62.1225 129.1315 62.2225 ;
      RECT MASK 2 4.672 62.395 10.96 62.495 ;
      RECT MASK 2 11.29 62.395 17.578 62.495 ;
      RECT MASK 2 17.908 62.395 24.196 62.495 ;
      RECT MASK 2 24.526 62.395 30.814 62.495 ;
      RECT MASK 2 31.144 62.395 37.432 62.495 ;
      RECT MASK 2 37.762 62.395 44.05 62.495 ;
      RECT MASK 2 44.38 62.395 50.668 62.495 ;
      RECT MASK 2 50.998 62.395 57.286 62.495 ;
      RECT MASK 2 57.616 62.395 63.904 62.495 ;
      RECT MASK 2 64.234 62.395 70.522 62.495 ;
      RECT MASK 2 70.852 62.395 77.14 62.495 ;
      RECT MASK 2 77.47 62.395 83.758 62.495 ;
      RECT MASK 2 84.088 62.395 90.376 62.495 ;
      RECT MASK 2 90.706 62.395 96.994 62.495 ;
      RECT MASK 2 97.324 62.395 103.612 62.495 ;
      RECT MASK 2 103.942 62.395 110.23 62.495 ;
      RECT MASK 2 111.044 62.6375 127.58 62.7375 ;
      RECT MASK 2 4.656 62.77 10.986 62.87 ;
      RECT MASK 2 11.274 62.77 17.604 62.87 ;
      RECT MASK 2 17.892 62.77 24.222 62.87 ;
      RECT MASK 2 24.51 62.77 30.84 62.87 ;
      RECT MASK 2 31.128 62.77 37.458 62.87 ;
      RECT MASK 2 37.746 62.77 44.076 62.87 ;
      RECT MASK 2 44.364 62.77 50.694 62.87 ;
      RECT MASK 2 50.982 62.77 57.312 62.87 ;
      RECT MASK 2 57.6 62.77 63.93 62.87 ;
      RECT MASK 2 64.218 62.77 70.548 62.87 ;
      RECT MASK 2 70.836 62.77 77.166 62.87 ;
      RECT MASK 2 77.454 62.77 83.784 62.87 ;
      RECT MASK 2 84.072 62.77 90.402 62.87 ;
      RECT MASK 2 90.69 62.77 97.02 62.87 ;
      RECT MASK 2 97.308 62.77 103.638 62.87 ;
      RECT MASK 2 103.926 62.77 110.256 62.87 ;
      RECT MASK 2 111.044 62.9575 129.1315 63.2075 ;
      RECT MASK 2 4.672 63.145 10.96 63.245 ;
      RECT MASK 2 11.29 63.145 17.578 63.245 ;
      RECT MASK 2 17.908 63.145 24.196 63.245 ;
      RECT MASK 2 24.526 63.145 30.814 63.245 ;
      RECT MASK 2 31.144 63.145 37.432 63.245 ;
      RECT MASK 2 37.762 63.145 44.05 63.245 ;
      RECT MASK 2 44.38 63.145 50.668 63.245 ;
      RECT MASK 2 50.998 63.145 57.286 63.245 ;
      RECT MASK 2 57.616 63.145 63.904 63.245 ;
      RECT MASK 2 64.234 63.145 70.522 63.245 ;
      RECT MASK 2 70.852 63.145 77.14 63.245 ;
      RECT MASK 2 77.47 63.145 83.758 63.245 ;
      RECT MASK 2 84.088 63.145 90.376 63.245 ;
      RECT MASK 2 90.706 63.145 96.994 63.245 ;
      RECT MASK 2 97.324 63.145 103.612 63.245 ;
      RECT MASK 2 103.942 63.145 110.23 63.245 ;
      RECT MASK 2 111.044 63.4725 129.1315 63.5725 ;
      RECT MASK 2 0.567 63.9 115.126 64.02 ;
      RECT MASK 2 117.268 64.0175 127.58 64.1175 ;
      RECT MASK 2 0.567 64.32 115.126 64.44 ;
      RECT MASK 2 117.268 64.3375 129.1315 64.5875 ;
      RECT MASK 2 111.044 64.8525 129.1315 64.9525 ;
      RECT MASK 2 4.672 65.155 10.96 65.255 ;
      RECT MASK 2 11.29 65.155 17.578 65.255 ;
      RECT MASK 2 17.908 65.155 24.196 65.255 ;
      RECT MASK 2 24.526 65.155 30.814 65.255 ;
      RECT MASK 2 31.144 65.155 37.432 65.255 ;
      RECT MASK 2 37.762 65.155 44.05 65.255 ;
      RECT MASK 2 44.38 65.155 50.668 65.255 ;
      RECT MASK 2 50.998 65.155 57.286 65.255 ;
      RECT MASK 2 57.616 65.155 63.904 65.255 ;
      RECT MASK 2 64.234 65.155 70.522 65.255 ;
      RECT MASK 2 70.852 65.155 77.14 65.255 ;
      RECT MASK 2 77.47 65.155 83.758 65.255 ;
      RECT MASK 2 84.088 65.155 90.376 65.255 ;
      RECT MASK 2 90.706 65.155 96.994 65.255 ;
      RECT MASK 2 97.324 65.155 103.612 65.255 ;
      RECT MASK 2 103.942 65.155 110.23 65.255 ;
      RECT MASK 2 111.044 65.3675 127.58 65.4675 ;
      RECT MASK 2 4.656 65.53 10.986 65.63 ;
      RECT MASK 2 11.274 65.53 17.604 65.63 ;
      RECT MASK 2 17.892 65.53 24.222 65.63 ;
      RECT MASK 2 24.51 65.53 30.84 65.63 ;
      RECT MASK 2 31.128 65.53 37.458 65.63 ;
      RECT MASK 2 37.746 65.53 44.076 65.63 ;
      RECT MASK 2 44.364 65.53 50.694 65.63 ;
      RECT MASK 2 50.982 65.53 57.312 65.63 ;
      RECT MASK 2 57.6 65.53 63.93 65.63 ;
      RECT MASK 2 64.218 65.53 70.548 65.63 ;
      RECT MASK 2 70.836 65.53 77.166 65.63 ;
      RECT MASK 2 77.454 65.53 83.784 65.63 ;
      RECT MASK 2 84.072 65.53 90.402 65.63 ;
      RECT MASK 2 90.69 65.53 97.02 65.63 ;
      RECT MASK 2 97.308 65.53 103.638 65.63 ;
      RECT MASK 2 103.926 65.53 110.256 65.63 ;
      RECT MASK 2 111.044 65.6875 129.1315 65.9375 ;
      RECT MASK 2 4.672 65.905 10.96 66.005 ;
      RECT MASK 2 11.29 65.905 17.578 66.005 ;
      RECT MASK 2 17.908 65.905 24.196 66.005 ;
      RECT MASK 2 24.526 65.905 30.814 66.005 ;
      RECT MASK 2 31.144 65.905 37.432 66.005 ;
      RECT MASK 2 37.762 65.905 44.05 66.005 ;
      RECT MASK 2 44.38 65.905 50.668 66.005 ;
      RECT MASK 2 50.998 65.905 57.286 66.005 ;
      RECT MASK 2 57.616 65.905 63.904 66.005 ;
      RECT MASK 2 64.234 65.905 70.522 66.005 ;
      RECT MASK 2 70.852 65.905 77.14 66.005 ;
      RECT MASK 2 77.47 65.905 83.758 66.005 ;
      RECT MASK 2 84.088 65.905 90.376 66.005 ;
      RECT MASK 2 90.706 65.905 96.994 66.005 ;
      RECT MASK 2 97.324 65.905 103.612 66.005 ;
      RECT MASK 2 103.942 65.905 110.23 66.005 ;
      RECT MASK 2 111.044 66.2025 129.1315 66.3025 ;
      RECT MASK 2 4.672 66.275 10.96 66.375 ;
      RECT MASK 2 11.29 66.275 17.578 66.375 ;
      RECT MASK 2 17.908 66.275 24.196 66.375 ;
      RECT MASK 2 24.526 66.275 30.814 66.375 ;
      RECT MASK 2 31.144 66.275 37.432 66.375 ;
      RECT MASK 2 37.762 66.275 44.05 66.375 ;
      RECT MASK 2 44.38 66.275 50.668 66.375 ;
      RECT MASK 2 50.998 66.275 57.286 66.375 ;
      RECT MASK 2 57.616 66.275 63.904 66.375 ;
      RECT MASK 2 64.234 66.275 70.522 66.375 ;
      RECT MASK 2 70.852 66.275 77.14 66.375 ;
      RECT MASK 2 77.47 66.275 83.758 66.375 ;
      RECT MASK 2 84.088 66.275 90.376 66.375 ;
      RECT MASK 2 90.706 66.275 96.994 66.375 ;
      RECT MASK 2 97.324 66.275 103.612 66.375 ;
      RECT MASK 2 103.942 66.275 110.23 66.375 ;
      RECT MASK 2 4.656 66.65 10.986 66.75 ;
      RECT MASK 2 11.274 66.65 17.604 66.75 ;
      RECT MASK 2 17.892 66.65 24.222 66.75 ;
      RECT MASK 2 24.51 66.65 30.84 66.75 ;
      RECT MASK 2 31.128 66.65 37.458 66.75 ;
      RECT MASK 2 37.746 66.65 44.076 66.75 ;
      RECT MASK 2 44.364 66.65 50.694 66.75 ;
      RECT MASK 2 50.982 66.65 57.312 66.75 ;
      RECT MASK 2 57.6 66.65 63.93 66.75 ;
      RECT MASK 2 64.218 66.65 70.548 66.75 ;
      RECT MASK 2 70.836 66.65 77.166 66.75 ;
      RECT MASK 2 77.454 66.65 83.784 66.75 ;
      RECT MASK 2 84.072 66.65 90.402 66.75 ;
      RECT MASK 2 90.69 66.65 97.02 66.75 ;
      RECT MASK 2 97.308 66.65 103.638 66.75 ;
      RECT MASK 2 103.926 66.65 110.256 66.75 ;
      RECT MASK 2 111.044 66.7175 127.58 66.8175 ;
      RECT MASK 2 4.672 67.025 10.96 67.125 ;
      RECT MASK 2 11.29 67.025 17.578 67.125 ;
      RECT MASK 2 17.908 67.025 24.196 67.125 ;
      RECT MASK 2 24.526 67.025 30.814 67.125 ;
      RECT MASK 2 31.144 67.025 37.432 67.125 ;
      RECT MASK 2 37.762 67.025 44.05 67.125 ;
      RECT MASK 2 44.38 67.025 50.668 67.125 ;
      RECT MASK 2 50.998 67.025 57.286 67.125 ;
      RECT MASK 2 57.616 67.025 63.904 67.125 ;
      RECT MASK 2 64.234 67.025 70.522 67.125 ;
      RECT MASK 2 70.852 67.025 77.14 67.125 ;
      RECT MASK 2 77.47 67.025 83.758 67.125 ;
      RECT MASK 2 84.088 67.025 90.376 67.125 ;
      RECT MASK 2 90.706 67.025 96.994 67.125 ;
      RECT MASK 2 97.324 67.025 103.612 67.125 ;
      RECT MASK 2 103.942 67.025 110.23 67.125 ;
      RECT MASK 2 111.044 67.0375 129.1315 67.2875 ;
      RECT MASK 2 4.672 67.395 10.96 67.495 ;
      RECT MASK 2 11.29 67.395 17.578 67.495 ;
      RECT MASK 2 17.908 67.395 24.196 67.495 ;
      RECT MASK 2 24.526 67.395 30.814 67.495 ;
      RECT MASK 2 31.144 67.395 37.432 67.495 ;
      RECT MASK 2 37.762 67.395 44.05 67.495 ;
      RECT MASK 2 44.38 67.395 50.668 67.495 ;
      RECT MASK 2 50.998 67.395 57.286 67.495 ;
      RECT MASK 2 57.616 67.395 63.904 67.495 ;
      RECT MASK 2 64.234 67.395 70.522 67.495 ;
      RECT MASK 2 70.852 67.395 77.14 67.495 ;
      RECT MASK 2 77.47 67.395 83.758 67.495 ;
      RECT MASK 2 84.088 67.395 90.376 67.495 ;
      RECT MASK 2 90.706 67.395 96.994 67.495 ;
      RECT MASK 2 97.324 67.395 103.612 67.495 ;
      RECT MASK 2 103.942 67.395 110.23 67.495 ;
      RECT MASK 2 111.044 67.5525 129.1315 67.6525 ;
      RECT MASK 2 4.656 67.77 10.986 67.87 ;
      RECT MASK 2 11.274 67.77 17.604 67.87 ;
      RECT MASK 2 17.892 67.77 24.222 67.87 ;
      RECT MASK 2 24.51 67.77 30.84 67.87 ;
      RECT MASK 2 31.128 67.77 37.458 67.87 ;
      RECT MASK 2 37.746 67.77 44.076 67.87 ;
      RECT MASK 2 44.364 67.77 50.694 67.87 ;
      RECT MASK 2 50.982 67.77 57.312 67.87 ;
      RECT MASK 2 57.6 67.77 63.93 67.87 ;
      RECT MASK 2 64.218 67.77 70.548 67.87 ;
      RECT MASK 2 70.836 67.77 77.166 67.87 ;
      RECT MASK 2 77.454 67.77 83.784 67.87 ;
      RECT MASK 2 84.072 67.77 90.402 67.87 ;
      RECT MASK 2 90.69 67.77 97.02 67.87 ;
      RECT MASK 2 97.308 67.77 103.638 67.87 ;
      RECT MASK 2 103.926 67.77 110.256 67.87 ;
      RECT MASK 2 111.044 68.0675 127.58 68.1675 ;
      RECT MASK 2 4.672 68.145 10.96 68.245 ;
      RECT MASK 2 11.29 68.145 17.578 68.245 ;
      RECT MASK 2 17.908 68.145 24.196 68.245 ;
      RECT MASK 2 24.526 68.145 30.814 68.245 ;
      RECT MASK 2 31.144 68.145 37.432 68.245 ;
      RECT MASK 2 37.762 68.145 44.05 68.245 ;
      RECT MASK 2 44.38 68.145 50.668 68.245 ;
      RECT MASK 2 50.998 68.145 57.286 68.245 ;
      RECT MASK 2 57.616 68.145 63.904 68.245 ;
      RECT MASK 2 64.234 68.145 70.522 68.245 ;
      RECT MASK 2 70.852 68.145 77.14 68.245 ;
      RECT MASK 2 77.47 68.145 83.758 68.245 ;
      RECT MASK 2 84.088 68.145 90.376 68.245 ;
      RECT MASK 2 90.706 68.145 96.994 68.245 ;
      RECT MASK 2 97.324 68.145 103.612 68.245 ;
      RECT MASK 2 103.942 68.145 110.23 68.245 ;
      RECT MASK 2 111.044 68.3875 129.1315 68.6375 ;
      RECT MASK 2 4.672 68.515 10.96 68.615 ;
      RECT MASK 2 11.29 68.515 17.578 68.615 ;
      RECT MASK 2 17.908 68.515 24.196 68.615 ;
      RECT MASK 2 24.526 68.515 30.814 68.615 ;
      RECT MASK 2 31.144 68.515 37.432 68.615 ;
      RECT MASK 2 37.762 68.515 44.05 68.615 ;
      RECT MASK 2 44.38 68.515 50.668 68.615 ;
      RECT MASK 2 50.998 68.515 57.286 68.615 ;
      RECT MASK 2 57.616 68.515 63.904 68.615 ;
      RECT MASK 2 64.234 68.515 70.522 68.615 ;
      RECT MASK 2 70.852 68.515 77.14 68.615 ;
      RECT MASK 2 77.47 68.515 83.758 68.615 ;
      RECT MASK 2 84.088 68.515 90.376 68.615 ;
      RECT MASK 2 90.706 68.515 96.994 68.615 ;
      RECT MASK 2 97.324 68.515 103.612 68.615 ;
      RECT MASK 2 103.942 68.515 110.23 68.615 ;
      RECT MASK 2 4.656 68.89 10.986 68.99 ;
      RECT MASK 2 11.274 68.89 17.604 68.99 ;
      RECT MASK 2 17.892 68.89 24.222 68.99 ;
      RECT MASK 2 24.51 68.89 30.84 68.99 ;
      RECT MASK 2 31.128 68.89 37.458 68.99 ;
      RECT MASK 2 37.746 68.89 44.076 68.99 ;
      RECT MASK 2 44.364 68.89 50.694 68.99 ;
      RECT MASK 2 50.982 68.89 57.312 68.99 ;
      RECT MASK 2 57.6 68.89 63.93 68.99 ;
      RECT MASK 2 64.218 68.89 70.548 68.99 ;
      RECT MASK 2 70.836 68.89 77.166 68.99 ;
      RECT MASK 2 77.454 68.89 83.784 68.99 ;
      RECT MASK 2 84.072 68.89 90.402 68.99 ;
      RECT MASK 2 90.69 68.89 97.02 68.99 ;
      RECT MASK 2 97.308 68.89 103.638 68.99 ;
      RECT MASK 2 103.926 68.89 110.256 68.99 ;
      RECT MASK 2 111.044 68.9025 129.1315 69.0025 ;
      RECT MASK 2 4.672 69.265 10.96 69.365 ;
      RECT MASK 2 11.29 69.265 17.578 69.365 ;
      RECT MASK 2 17.908 69.265 24.196 69.365 ;
      RECT MASK 2 24.526 69.265 30.814 69.365 ;
      RECT MASK 2 31.144 69.265 37.432 69.365 ;
      RECT MASK 2 37.762 69.265 44.05 69.365 ;
      RECT MASK 2 44.38 69.265 50.668 69.365 ;
      RECT MASK 2 50.998 69.265 57.286 69.365 ;
      RECT MASK 2 57.616 69.265 63.904 69.365 ;
      RECT MASK 2 64.234 69.265 70.522 69.365 ;
      RECT MASK 2 70.852 69.265 77.14 69.365 ;
      RECT MASK 2 77.47 69.265 83.758 69.365 ;
      RECT MASK 2 84.088 69.265 90.376 69.365 ;
      RECT MASK 2 90.706 69.265 96.994 69.365 ;
      RECT MASK 2 97.324 69.265 103.612 69.365 ;
      RECT MASK 2 103.942 69.265 110.23 69.365 ;
      RECT MASK 2 111.044 69.4175 127.58 69.5175 ;
      RECT MASK 2 117.268 69.7375 129.1315 69.9875 ;
      RECT MASK 2 0.567 70.02 115.126 70.14 ;
      RECT MASK 2 0.567 70.44 129.1315 70.56 ;
      RECT MASK 2 4.672 71.275 17.578 71.375 ;
      RECT MASK 2 17.908 71.275 30.814 71.375 ;
      RECT MASK 2 31.144 71.275 44.05 71.375 ;
      RECT MASK 2 44.38 71.275 57.286 71.375 ;
      RECT MASK 2 57.616 71.275 70.522 71.375 ;
      RECT MASK 2 70.852 71.275 83.758 71.375 ;
      RECT MASK 2 84.088 71.275 96.994 71.375 ;
      RECT MASK 2 97.324 71.275 110.23 71.375 ;
      RECT MASK 2 4.656 71.65 17.604 71.75 ;
      RECT MASK 2 17.892 71.65 30.84 71.75 ;
      RECT MASK 2 31.128 71.65 44.076 71.75 ;
      RECT MASK 2 44.364 71.65 57.312 71.75 ;
      RECT MASK 2 57.6 71.65 70.548 71.75 ;
      RECT MASK 2 70.836 71.65 83.784 71.75 ;
      RECT MASK 2 84.072 71.65 97.02 71.75 ;
      RECT MASK 2 97.308 71.65 110.256 71.75 ;
      RECT MASK 2 4.672 72.025 17.578 72.125 ;
      RECT MASK 2 17.908 72.025 30.814 72.125 ;
      RECT MASK 2 31.144 72.025 44.05 72.125 ;
      RECT MASK 2 44.38 72.025 57.286 72.125 ;
      RECT MASK 2 57.616 72.025 70.522 72.125 ;
      RECT MASK 2 70.852 72.025 83.758 72.125 ;
      RECT MASK 2 84.088 72.025 96.994 72.125 ;
      RECT MASK 2 97.324 72.025 110.23 72.125 ;
      RECT MASK 2 4.672 72.395 17.578 72.495 ;
      RECT MASK 2 17.908 72.395 30.814 72.495 ;
      RECT MASK 2 31.144 72.395 44.05 72.495 ;
      RECT MASK 2 44.38 72.395 57.286 72.495 ;
      RECT MASK 2 57.616 72.395 70.522 72.495 ;
      RECT MASK 2 70.852 72.395 83.758 72.495 ;
      RECT MASK 2 84.088 72.395 96.994 72.495 ;
      RECT MASK 2 97.324 72.395 110.23 72.495 ;
      RECT MASK 2 4.656 72.77 17.604 72.87 ;
      RECT MASK 2 17.892 72.77 30.84 72.87 ;
      RECT MASK 2 31.128 72.77 44.076 72.87 ;
      RECT MASK 2 44.364 72.77 57.312 72.87 ;
      RECT MASK 2 57.6 72.77 70.548 72.87 ;
      RECT MASK 2 70.836 72.77 83.784 72.87 ;
      RECT MASK 2 84.072 72.77 97.02 72.87 ;
      RECT MASK 2 97.308 72.77 110.256 72.87 ;
      RECT MASK 2 4.672 73.145 17.578 73.245 ;
      RECT MASK 2 17.908 73.145 30.814 73.245 ;
      RECT MASK 2 31.144 73.145 44.05 73.245 ;
      RECT MASK 2 44.38 73.145 57.286 73.245 ;
      RECT MASK 2 57.616 73.145 70.522 73.245 ;
      RECT MASK 2 70.852 73.145 83.758 73.245 ;
      RECT MASK 2 84.088 73.145 96.994 73.245 ;
      RECT MASK 2 97.324 73.145 110.23 73.245 ;
      RECT MASK 2 4.672 73.515 17.578 73.615 ;
      RECT MASK 2 17.908 73.515 30.814 73.615 ;
      RECT MASK 2 31.144 73.515 44.05 73.615 ;
      RECT MASK 2 44.38 73.515 57.286 73.615 ;
      RECT MASK 2 57.616 73.515 70.522 73.615 ;
      RECT MASK 2 70.852 73.515 83.758 73.615 ;
      RECT MASK 2 84.088 73.515 96.994 73.615 ;
      RECT MASK 2 97.324 73.515 110.23 73.615 ;
      RECT MASK 2 116.163 73.74 126.333 73.94 ;
      RECT MASK 2 4.656 73.89 17.604 73.99 ;
      RECT MASK 2 17.892 73.89 30.84 73.99 ;
      RECT MASK 2 31.128 73.89 44.076 73.99 ;
      RECT MASK 2 44.364 73.89 57.312 73.99 ;
      RECT MASK 2 57.6 73.89 70.548 73.99 ;
      RECT MASK 2 70.836 73.89 83.784 73.99 ;
      RECT MASK 2 84.072 73.89 97.02 73.99 ;
      RECT MASK 2 97.308 73.89 110.256 73.99 ;
      RECT MASK 2 4.672 74.265 17.578 74.365 ;
      RECT MASK 2 17.908 74.265 30.814 74.365 ;
      RECT MASK 2 31.144 74.265 44.05 74.365 ;
      RECT MASK 2 44.38 74.265 57.286 74.365 ;
      RECT MASK 2 57.616 74.265 70.522 74.365 ;
      RECT MASK 2 70.852 74.265 83.758 74.365 ;
      RECT MASK 2 84.088 74.265 96.994 74.365 ;
      RECT MASK 2 97.324 74.265 110.23 74.365 ;
      RECT MASK 2 116.218 74.338 126.339 74.398 ;
      RECT MASK 2 4.672 74.635 17.578 74.735 ;
      RECT MASK 2 17.908 74.635 30.814 74.735 ;
      RECT MASK 2 31.144 74.635 44.05 74.735 ;
      RECT MASK 2 44.38 74.635 57.286 74.735 ;
      RECT MASK 2 57.616 74.635 70.522 74.735 ;
      RECT MASK 2 70.852 74.635 83.758 74.735 ;
      RECT MASK 2 84.088 74.635 96.994 74.735 ;
      RECT MASK 2 97.324 74.635 110.23 74.735 ;
      RECT MASK 2 116.163 74.78 126.333 74.98 ;
      RECT MASK 2 4.656 75.01 17.604 75.11 ;
      RECT MASK 2 17.892 75.01 30.84 75.11 ;
      RECT MASK 2 31.128 75.01 44.076 75.11 ;
      RECT MASK 2 44.364 75.01 57.312 75.11 ;
      RECT MASK 2 57.6 75.01 70.548 75.11 ;
      RECT MASK 2 70.836 75.01 83.784 75.11 ;
      RECT MASK 2 84.072 75.01 97.02 75.11 ;
      RECT MASK 2 97.308 75.01 110.256 75.11 ;
      RECT MASK 2 116.162 75.3 126.332 75.5 ;
      RECT MASK 2 4.672 75.385 17.578 75.485 ;
      RECT MASK 2 17.908 75.385 30.814 75.485 ;
      RECT MASK 2 31.144 75.385 44.05 75.485 ;
      RECT MASK 2 44.38 75.385 57.286 75.485 ;
      RECT MASK 2 57.616 75.385 70.522 75.485 ;
      RECT MASK 2 70.852 75.385 83.758 75.485 ;
      RECT MASK 2 84.088 75.385 96.994 75.485 ;
      RECT MASK 2 97.324 75.385 110.23 75.485 ;
      RECT MASK 2 116.218 75.883 126.339 75.943 ;
      RECT MASK 2 116.163 76.34 126.333 76.54 ;
      RECT MASK 2 116.163 76.86 126.333 77.06 ;
      RECT MASK 2 116.218 77.458 126.339 77.518 ;
      RECT MASK 2 115.515 77.9 126.969 78.1 ;
      RECT MASK 2 6.165 78.105 114.086 78.225 ;
      RECT MASK 2 116.163 78.42 126.333 78.62 ;
      RECT MASK 2 6.941 78.751 7.2505 78.811 ;
      RECT MASK 2 8.103 78.751 8.4125 78.811 ;
      RECT MASK 2 9.265 78.751 9.5745 78.811 ;
      RECT MASK 2 12.397 78.751 12.7065 78.811 ;
      RECT MASK 2 13.559 78.751 13.8685 78.811 ;
      RECT MASK 2 14.721 78.751 15.0305 78.811 ;
      RECT MASK 2 15.883 78.751 16.1925 78.811 ;
      RECT MASK 2 19.015 78.751 19.3245 78.811 ;
      RECT MASK 2 20.177 78.751 20.4865 78.811 ;
      RECT MASK 2 21.339 78.751 21.6485 78.811 ;
      RECT MASK 2 22.501 78.751 22.8105 78.811 ;
      RECT MASK 2 25.633 78.751 25.9425 78.811 ;
      RECT MASK 2 26.795 78.751 27.1045 78.811 ;
      RECT MASK 2 27.957 78.751 28.2665 78.811 ;
      RECT MASK 2 29.119 78.751 29.4285 78.811 ;
      RECT MASK 2 32.251 78.751 32.5605 78.811 ;
      RECT MASK 2 33.413 78.751 33.7225 78.811 ;
      RECT MASK 2 34.575 78.751 34.8845 78.811 ;
      RECT MASK 2 35.737 78.751 36.0465 78.811 ;
      RECT MASK 2 38.869 78.751 39.1785 78.811 ;
      RECT MASK 2 40.031 78.751 40.3405 78.811 ;
      RECT MASK 2 41.193 78.751 41.5025 78.811 ;
      RECT MASK 2 42.355 78.751 42.6645 78.811 ;
      RECT MASK 2 45.487 78.751 45.7965 78.811 ;
      RECT MASK 2 46.649 78.751 46.9585 78.811 ;
      RECT MASK 2 47.811 78.751 48.1205 78.811 ;
      RECT MASK 2 48.973 78.751 49.2825 78.811 ;
      RECT MASK 2 52.105 78.751 52.4145 78.811 ;
      RECT MASK 2 53.267 78.751 53.5765 78.811 ;
      RECT MASK 2 54.429 78.751 54.7385 78.811 ;
      RECT MASK 2 55.591 78.751 55.9005 78.811 ;
      RECT MASK 2 58.723 78.751 59.0325 78.811 ;
      RECT MASK 2 59.885 78.751 60.1945 78.811 ;
      RECT MASK 2 61.047 78.751 61.3565 78.811 ;
      RECT MASK 2 62.209 78.751 62.5185 78.811 ;
      RECT MASK 2 65.341 78.751 65.6505 78.811 ;
      RECT MASK 2 66.503 78.751 66.8125 78.811 ;
      RECT MASK 2 67.665 78.751 67.9745 78.811 ;
      RECT MASK 2 68.827 78.751 69.1365 78.811 ;
      RECT MASK 2 71.959 78.751 72.2685 78.811 ;
      RECT MASK 2 73.121 78.751 73.4305 78.811 ;
      RECT MASK 2 74.283 78.751 74.5925 78.811 ;
      RECT MASK 2 75.445 78.751 75.7545 78.811 ;
      RECT MASK 2 78.577 78.751 78.8865 78.811 ;
      RECT MASK 2 79.739 78.751 80.0485 78.811 ;
      RECT MASK 2 80.901 78.751 81.2105 78.811 ;
      RECT MASK 2 82.063 78.751 82.3725 78.811 ;
      RECT MASK 2 85.195 78.751 85.5045 78.811 ;
      RECT MASK 2 86.357 78.751 86.6665 78.811 ;
      RECT MASK 2 87.519 78.751 87.8285 78.811 ;
      RECT MASK 2 88.681 78.751 88.9905 78.811 ;
      RECT MASK 2 91.813 78.751 92.1225 78.811 ;
      RECT MASK 2 92.975 78.751 93.2845 78.811 ;
      RECT MASK 2 94.137 78.751 94.4465 78.811 ;
      RECT MASK 2 95.299 78.751 95.6085 78.811 ;
      RECT MASK 2 98.431 78.751 98.7405 78.811 ;
      RECT MASK 2 99.593 78.751 99.9025 78.811 ;
      RECT MASK 2 100.755 78.751 101.0645 78.811 ;
      RECT MASK 2 101.917 78.751 102.2265 78.811 ;
      RECT MASK 2 105.049 78.751 105.3585 78.811 ;
      RECT MASK 2 106.211 78.751 106.5205 78.811 ;
      RECT MASK 2 107.373 78.751 107.6825 78.811 ;
      RECT MASK 2 108.535 78.751 108.8445 78.811 ;
      RECT MASK 2 116.218 79.012 126.339 79.072 ;
      RECT MASK 2 6.941 79.231 7.267 79.291 ;
      RECT MASK 2 8.103 79.231 8.429 79.291 ;
      RECT MASK 2 9.265 79.231 9.591 79.291 ;
      RECT MASK 2 12.397 79.231 12.723 79.291 ;
      RECT MASK 2 13.559 79.231 13.885 79.291 ;
      RECT MASK 2 14.721 79.231 15.047 79.291 ;
      RECT MASK 2 15.883 79.231 16.209 79.291 ;
      RECT MASK 2 19.015 79.231 19.341 79.291 ;
      RECT MASK 2 20.177 79.231 20.503 79.291 ;
      RECT MASK 2 21.339 79.231 21.665 79.291 ;
      RECT MASK 2 22.501 79.231 22.827 79.291 ;
      RECT MASK 2 25.633 79.231 25.959 79.291 ;
      RECT MASK 2 26.795 79.231 27.121 79.291 ;
      RECT MASK 2 27.957 79.231 28.283 79.291 ;
      RECT MASK 2 29.119 79.231 29.445 79.291 ;
      RECT MASK 2 32.251 79.231 32.577 79.291 ;
      RECT MASK 2 33.413 79.231 33.739 79.291 ;
      RECT MASK 2 34.575 79.231 34.901 79.291 ;
      RECT MASK 2 35.737 79.231 36.063 79.291 ;
      RECT MASK 2 38.869 79.231 39.195 79.291 ;
      RECT MASK 2 40.031 79.231 40.357 79.291 ;
      RECT MASK 2 41.193 79.231 41.519 79.291 ;
      RECT MASK 2 42.355 79.231 42.681 79.291 ;
      RECT MASK 2 45.487 79.231 45.813 79.291 ;
      RECT MASK 2 46.649 79.231 46.975 79.291 ;
      RECT MASK 2 47.811 79.231 48.137 79.291 ;
      RECT MASK 2 48.973 79.231 49.299 79.291 ;
      RECT MASK 2 52.105 79.231 52.431 79.291 ;
      RECT MASK 2 53.267 79.231 53.593 79.291 ;
      RECT MASK 2 54.429 79.231 54.755 79.291 ;
      RECT MASK 2 55.591 79.231 55.917 79.291 ;
      RECT MASK 2 58.723 79.231 59.049 79.291 ;
      RECT MASK 2 59.885 79.231 60.211 79.291 ;
      RECT MASK 2 61.047 79.231 61.373 79.291 ;
      RECT MASK 2 62.209 79.231 62.535 79.291 ;
      RECT MASK 2 65.341 79.231 65.667 79.291 ;
      RECT MASK 2 66.503 79.231 66.829 79.291 ;
      RECT MASK 2 67.665 79.231 67.991 79.291 ;
      RECT MASK 2 68.827 79.231 69.153 79.291 ;
      RECT MASK 2 71.959 79.231 72.285 79.291 ;
      RECT MASK 2 73.121 79.231 73.447 79.291 ;
      RECT MASK 2 74.283 79.231 74.609 79.291 ;
      RECT MASK 2 75.445 79.231 75.771 79.291 ;
      RECT MASK 2 78.577 79.231 78.903 79.291 ;
      RECT MASK 2 79.739 79.231 80.065 79.291 ;
      RECT MASK 2 80.901 79.231 81.227 79.291 ;
      RECT MASK 2 82.063 79.231 82.389 79.291 ;
      RECT MASK 2 85.195 79.231 85.521 79.291 ;
      RECT MASK 2 86.357 79.231 86.683 79.291 ;
      RECT MASK 2 87.519 79.231 87.845 79.291 ;
      RECT MASK 2 88.681 79.231 89.007 79.291 ;
      RECT MASK 2 91.813 79.231 92.139 79.291 ;
      RECT MASK 2 92.975 79.231 93.301 79.291 ;
      RECT MASK 2 94.137 79.231 94.463 79.291 ;
      RECT MASK 2 95.299 79.231 95.625 79.291 ;
      RECT MASK 2 98.431 79.231 98.757 79.291 ;
      RECT MASK 2 99.593 79.231 99.919 79.291 ;
      RECT MASK 2 100.755 79.231 101.081 79.291 ;
      RECT MASK 2 101.917 79.231 102.243 79.291 ;
      RECT MASK 2 105.049 79.231 105.375 79.291 ;
      RECT MASK 2 106.211 79.231 106.537 79.291 ;
      RECT MASK 2 107.373 79.231 107.699 79.291 ;
      RECT MASK 2 108.535 79.231 108.861 79.291 ;
      RECT MASK 2 1.1745 79.27 5.417 79.31 ;
      RECT MASK 2 111.186 79.29 113.365 79.47 ;
      RECT MASK 2 115.515 79.46 126.969 79.66 ;
      RECT MASK 2 1.1745 79.51 5.417 79.55 ;
      RECT MASK 2 1.1745 79.75 5.417 79.79 ;
      RECT MASK 2 1.1745 79.99 5.417 80.03 ;
      RECT MASK 2 6.481 80.055 10.382 80.175 ;
      RECT MASK 2 11.937 80.055 17 80.175 ;
      RECT MASK 2 18.555 80.055 23.618 80.175 ;
      RECT MASK 2 25.173 80.055 30.236 80.175 ;
      RECT MASK 2 31.791 80.055 36.854 80.175 ;
      RECT MASK 2 38.409 80.055 43.472 80.175 ;
      RECT MASK 2 45.027 80.055 50.09 80.175 ;
      RECT MASK 2 51.645 80.055 56.708 80.175 ;
      RECT MASK 2 58.263 80.055 63.326 80.175 ;
      RECT MASK 2 64.881 80.055 69.944 80.175 ;
      RECT MASK 2 71.499 80.055 76.562 80.175 ;
      RECT MASK 2 78.117 80.055 83.18 80.175 ;
      RECT MASK 2 84.735 80.055 89.798 80.175 ;
      RECT MASK 2 91.353 80.055 96.416 80.175 ;
      RECT MASK 2 97.971 80.055 103.034 80.175 ;
      RECT MASK 2 104.589 80.055 109.652 80.175 ;
      RECT MASK 2 1.1745 80.23 5.417 80.27 ;
      RECT MASK 2 57.178 80.465 64.425 80.665 ;
      RECT MASK 2 1.1745 80.47 5.417 80.51 ;
      RECT MASK 2 6.481 80.505 10.382 80.625 ;
      RECT MASK 2 11.937 80.505 17 80.625 ;
      RECT MASK 2 18.555 80.505 23.618 80.625 ;
      RECT MASK 2 25.173 80.505 30.236 80.625 ;
      RECT MASK 2 31.791 80.505 36.854 80.625 ;
      RECT MASK 2 38.409 80.505 43.472 80.625 ;
      RECT MASK 2 45.027 80.505 50.09 80.625 ;
      RECT MASK 2 51.645 80.505 56.708 80.625 ;
      RECT MASK 2 64.881 80.505 69.944 80.625 ;
      RECT MASK 2 71.499 80.505 76.562 80.625 ;
      RECT MASK 2 78.117 80.505 83.18 80.625 ;
      RECT MASK 2 84.735 80.505 89.798 80.625 ;
      RECT MASK 2 91.353 80.505 96.416 80.625 ;
      RECT MASK 2 97.971 80.505 103.034 80.625 ;
      RECT MASK 2 104.589 80.505 109.652 80.625 ;
      RECT MASK 2 111.1115 80.658 113.324 80.838 ;
      RECT MASK 2 1.1745 80.71 5.417 80.75 ;
      RECT MASK 2 57.178 80.91 59.7205 80.97 ;
      RECT MASK 2 63.0635 80.91 64.425 80.97 ;
      RECT MASK 2 1.1745 80.95 5.417 80.99 ;
      RECT MASK 2 6.941 81.15 7.267 81.21 ;
      RECT MASK 2 8.103 81.15 8.429 81.21 ;
      RECT MASK 2 9.265 81.15 9.591 81.21 ;
      RECT MASK 2 12.397 81.15 12.723 81.21 ;
      RECT MASK 2 13.559 81.15 13.885 81.21 ;
      RECT MASK 2 14.721 81.15 15.047 81.21 ;
      RECT MASK 2 15.883 81.15 16.209 81.21 ;
      RECT MASK 2 19.015 81.15 19.341 81.21 ;
      RECT MASK 2 20.177 81.15 20.503 81.21 ;
      RECT MASK 2 21.339 81.15 21.665 81.21 ;
      RECT MASK 2 22.501 81.15 22.827 81.21 ;
      RECT MASK 2 25.633 81.15 25.959 81.21 ;
      RECT MASK 2 26.795 81.15 27.121 81.21 ;
      RECT MASK 2 27.957 81.15 28.283 81.21 ;
      RECT MASK 2 29.119 81.15 29.445 81.21 ;
      RECT MASK 2 32.251 81.15 32.577 81.21 ;
      RECT MASK 2 33.413 81.15 33.739 81.21 ;
      RECT MASK 2 34.575 81.15 34.901 81.21 ;
      RECT MASK 2 35.737 81.15 36.063 81.21 ;
      RECT MASK 2 38.869 81.15 39.195 81.21 ;
      RECT MASK 2 40.031 81.15 40.357 81.21 ;
      RECT MASK 2 41.193 81.15 41.519 81.21 ;
      RECT MASK 2 42.355 81.15 42.681 81.21 ;
      RECT MASK 2 45.487 81.15 45.813 81.21 ;
      RECT MASK 2 46.649 81.15 46.975 81.21 ;
      RECT MASK 2 47.811 81.15 48.137 81.21 ;
      RECT MASK 2 48.973 81.15 49.299 81.21 ;
      RECT MASK 2 52.105 81.15 52.431 81.21 ;
      RECT MASK 2 53.267 81.15 53.593 81.21 ;
      RECT MASK 2 54.429 81.15 54.755 81.21 ;
      RECT MASK 2 55.591 81.15 55.917 81.21 ;
      RECT MASK 2 57.178 81.15 58.3635 81.21 ;
      RECT MASK 2 58.723 81.15 59.049 81.21 ;
      RECT MASK 2 59.885 81.15 60.211 81.21 ;
      RECT MASK 2 61.047 81.15 61.373 81.21 ;
      RECT MASK 2 62.209 81.15 62.535 81.21 ;
      RECT MASK 2 65.341 81.15 65.667 81.21 ;
      RECT MASK 2 66.503 81.15 66.829 81.21 ;
      RECT MASK 2 67.665 81.15 67.991 81.21 ;
      RECT MASK 2 68.827 81.15 69.153 81.21 ;
      RECT MASK 2 71.959 81.15 72.285 81.21 ;
      RECT MASK 2 73.121 81.15 73.447 81.21 ;
      RECT MASK 2 74.283 81.15 74.609 81.21 ;
      RECT MASK 2 75.445 81.15 75.771 81.21 ;
      RECT MASK 2 78.577 81.15 78.903 81.21 ;
      RECT MASK 2 79.739 81.15 80.065 81.21 ;
      RECT MASK 2 80.901 81.15 81.227 81.21 ;
      RECT MASK 2 82.063 81.15 82.389 81.21 ;
      RECT MASK 2 85.195 81.15 85.521 81.21 ;
      RECT MASK 2 86.357 81.15 86.683 81.21 ;
      RECT MASK 2 87.519 81.15 87.845 81.21 ;
      RECT MASK 2 88.681 81.15 89.007 81.21 ;
      RECT MASK 2 91.813 81.15 92.139 81.21 ;
      RECT MASK 2 92.975 81.15 93.301 81.21 ;
      RECT MASK 2 94.137 81.15 94.463 81.21 ;
      RECT MASK 2 95.299 81.15 95.625 81.21 ;
      RECT MASK 2 98.431 81.15 98.757 81.21 ;
      RECT MASK 2 99.593 81.15 99.919 81.21 ;
      RECT MASK 2 100.755 81.15 101.081 81.21 ;
      RECT MASK 2 101.917 81.15 102.243 81.21 ;
      RECT MASK 2 105.049 81.15 105.375 81.21 ;
      RECT MASK 2 106.211 81.15 106.537 81.21 ;
      RECT MASK 2 107.373 81.15 107.699 81.21 ;
      RECT MASK 2 108.535 81.15 108.861 81.21 ;
      RECT MASK 2 1.1745 81.19 5.417 81.23 ;
      RECT MASK 2 63.0635 81.25 64.425 81.31 ;
      RECT MASK 2 1.1745 81.43 5.417 81.47 ;
      RECT MASK 2 6.941 81.63 7.267 81.69 ;
      RECT MASK 2 8.103 81.63 8.429 81.69 ;
      RECT MASK 2 9.265 81.63 9.591 81.69 ;
      RECT MASK 2 12.397 81.63 12.723 81.69 ;
      RECT MASK 2 13.559 81.63 13.885 81.69 ;
      RECT MASK 2 14.721 81.63 15.047 81.69 ;
      RECT MASK 2 15.883 81.63 16.209 81.69 ;
      RECT MASK 2 19.015 81.63 19.341 81.69 ;
      RECT MASK 2 20.177 81.63 20.503 81.69 ;
      RECT MASK 2 21.339 81.63 21.665 81.69 ;
      RECT MASK 2 22.501 81.63 22.827 81.69 ;
      RECT MASK 2 25.633 81.63 25.959 81.69 ;
      RECT MASK 2 26.795 81.63 27.121 81.69 ;
      RECT MASK 2 27.957 81.63 28.283 81.69 ;
      RECT MASK 2 29.119 81.63 29.445 81.69 ;
      RECT MASK 2 32.251 81.63 32.577 81.69 ;
      RECT MASK 2 33.413 81.63 33.739 81.69 ;
      RECT MASK 2 34.575 81.63 34.901 81.69 ;
      RECT MASK 2 35.737 81.63 36.063 81.69 ;
      RECT MASK 2 38.869 81.63 39.195 81.69 ;
      RECT MASK 2 40.031 81.63 40.357 81.69 ;
      RECT MASK 2 41.193 81.63 41.519 81.69 ;
      RECT MASK 2 42.355 81.63 42.681 81.69 ;
      RECT MASK 2 45.487 81.63 45.813 81.69 ;
      RECT MASK 2 46.649 81.63 46.975 81.69 ;
      RECT MASK 2 47.811 81.63 48.137 81.69 ;
      RECT MASK 2 48.973 81.63 49.299 81.69 ;
      RECT MASK 2 52.105 81.63 52.431 81.69 ;
      RECT MASK 2 53.267 81.63 53.593 81.69 ;
      RECT MASK 2 54.429 81.63 54.755 81.69 ;
      RECT MASK 2 55.591 81.63 55.917 81.69 ;
      RECT MASK 2 57.178 81.63 58.386 81.69 ;
      RECT MASK 2 58.723 81.63 59.049 81.69 ;
      RECT MASK 2 59.885 81.63 60.211 81.69 ;
      RECT MASK 2 61.047 81.63 61.373 81.69 ;
      RECT MASK 2 62.209 81.63 62.535 81.69 ;
      RECT MASK 2 63.0635 81.63 64.425 81.69 ;
      RECT MASK 2 65.341 81.63 65.667 81.69 ;
      RECT MASK 2 66.503 81.63 66.829 81.69 ;
      RECT MASK 2 67.665 81.63 67.991 81.69 ;
      RECT MASK 2 68.827 81.63 69.153 81.69 ;
      RECT MASK 2 71.959 81.63 72.285 81.69 ;
      RECT MASK 2 73.121 81.63 73.447 81.69 ;
      RECT MASK 2 74.283 81.63 74.609 81.69 ;
      RECT MASK 2 75.445 81.63 75.771 81.69 ;
      RECT MASK 2 78.577 81.63 78.903 81.69 ;
      RECT MASK 2 79.739 81.63 80.065 81.69 ;
      RECT MASK 2 80.901 81.63 81.227 81.69 ;
      RECT MASK 2 82.063 81.63 82.389 81.69 ;
      RECT MASK 2 85.195 81.63 85.521 81.69 ;
      RECT MASK 2 86.357 81.63 86.683 81.69 ;
      RECT MASK 2 87.519 81.63 87.845 81.69 ;
      RECT MASK 2 88.681 81.63 89.007 81.69 ;
      RECT MASK 2 91.813 81.63 92.139 81.69 ;
      RECT MASK 2 92.975 81.63 93.301 81.69 ;
      RECT MASK 2 94.137 81.63 94.463 81.69 ;
      RECT MASK 2 95.299 81.63 95.625 81.69 ;
      RECT MASK 2 98.431 81.63 98.757 81.69 ;
      RECT MASK 2 99.593 81.63 99.919 81.69 ;
      RECT MASK 2 100.755 81.63 101.081 81.69 ;
      RECT MASK 2 101.917 81.63 102.243 81.69 ;
      RECT MASK 2 105.049 81.63 105.375 81.69 ;
      RECT MASK 2 106.211 81.63 106.537 81.69 ;
      RECT MASK 2 107.373 81.63 107.699 81.69 ;
      RECT MASK 2 108.535 81.63 108.861 81.69 ;
      RECT MASK 2 1.1745 81.67 5.417 81.71 ;
      RECT MASK 2 57.178 81.903 59.7145 81.963 ;
      RECT MASK 2 63.0635 81.903 64.425 81.963 ;
      RECT MASK 2 1.1745 81.91 5.417 81.95 ;
      RECT MASK 2 115.5395 82.06 128.5785 82.1 ;
      RECT MASK 2 57.178 82.143 64.425 82.203 ;
      RECT MASK 2 1.1745 82.15 5.417 82.19 ;
      RECT MASK 2 115.5395 82.3 128.5785 82.34 ;
      RECT MASK 2 1.1745 82.39 5.417 82.43 ;
      RECT MASK 2 6.181 82.415 56.9 82.615 ;
      RECT MASK 2 64.694 82.415 113.11 82.615 ;
      RECT MASK 2 57.174 82.485 64.42 82.545 ;
      RECT MASK 2 115.5395 82.54 128.5785 82.58 ;
      RECT MASK 2 1.1745 82.63 5.417 82.67 ;
      RECT MASK 2 57.178 82.725 64.425 82.785 ;
      RECT MASK 2 115.5395 82.78 128.5785 82.82 ;
      RECT MASK 2 1.1745 82.87 5.417 82.91 ;
      RECT MASK 2 115.5395 83.02 128.5785 83.06 ;
      RECT MASK 2 1.1745 83.11 5.417 83.15 ;
      RECT MASK 2 57.178 83.14 64.425 83.2 ;
      RECT MASK 2 115.5395 83.26 128.5785 83.3 ;
      RECT MASK 2 1.1745 83.35 5.417 83.39 ;
      RECT MASK 2 57.178 83.38 64.425 83.44 ;
      RECT MASK 2 115.5395 83.5 128.5785 83.54 ;
      RECT MASK 2 1.1745 83.59 5.417 83.63 ;
      RECT MASK 2 115.5395 83.74 128.5785 83.78 ;
      RECT MASK 2 1.1745 83.83 5.417 83.87 ;
      RECT MASK 2 6.193 83.962 56.89 84.162 ;
      RECT MASK 2 57.174 83.962 64.42 84.162 ;
      RECT MASK 2 64.694 83.962 113.11 84.162 ;
      RECT MASK 2 115.5395 83.98 128.5785 84.02 ;
      RECT MASK 2 1.1745 84.07 5.417 84.11 ;
      RECT MASK 2 115.5395 84.22 128.5785 84.26 ;
      RECT MASK 2 1.1745 84.31 5.417 84.35 ;
      RECT MASK 2 115.5395 84.46 128.5785 84.5 ;
      RECT MASK 2 1.1745 84.55 5.417 84.59 ;
      RECT MASK 2 115.5395 84.7 128.5785 84.74 ;
      RECT MASK 2 1.1745 84.79 5.417 84.83 ;
      RECT MASK 2 115.5395 84.94 128.5785 84.98 ;
      RECT MASK 2 1.1745 85.03 5.417 85.07 ;
      RECT MASK 2 115.5395 85.18 128.5785 85.22 ;
      RECT MASK 2 1.1745 85.27 5.417 85.31 ;
      RECT MASK 2 6.193 85.35 113.373 85.53 ;
      RECT MASK 2 115.5395 85.42 128.5785 85.46 ;
      RECT MASK 2 1.1745 85.51 5.417 85.55 ;
      RECT MASK 2 115.5395 85.66 128.5785 85.7 ;
      RECT MASK 2 1.1745 85.75 5.417 85.79 ;
      RECT MASK 2 115.5395 85.9 128.5785 85.94 ;
      RECT MASK 2 1.1745 85.99 5.417 86.03 ;
      RECT MASK 2 115.5395 86.14 128.5785 86.18 ;
      RECT MASK 2 1.1745 86.23 5.417 86.27 ;
      RECT MASK 2 115.5395 86.38 128.5785 86.42 ;
      RECT MASK 2 1.1745 86.47 5.417 86.51 ;
      RECT MASK 2 115.5395 86.62 128.5785 86.66 ;
      RECT MASK 2 1.1745 86.71 5.417 86.75 ;
      RECT MASK 2 1.1745 86.95 5.417 86.99 ;
      RECT MASK 2 36.326 87.021 66.476 87.081 ;
      RECT MASK 2 72.716 87.021 102.866 87.081 ;
      RECT MASK 2 25.68 87.096 25.74 88.922 ;
      RECT MASK 2 26.048 87.096 26.108 88.922 ;
      RECT MASK 2 26.36 87.096 26.42 88.922 ;
      RECT MASK 2 26.63 87.096 26.69 88.921 ;
      RECT MASK 2 26.9 87.096 26.96 88.921 ;
      RECT MASK 2 27.17 87.096 27.23 88.921 ;
      RECT MASK 2 27.44 87.096 27.5 88.921 ;
      RECT MASK 2 27.71 87.096 27.77 88.921 ;
      RECT MASK 2 27.98 87.096 28.04 88.921 ;
      RECT MASK 2 28.25 87.096 28.31 88.921 ;
      RECT MASK 2 28.52 87.096 28.58 88.921 ;
      RECT MASK 2 28.79 87.096 28.85 88.921 ;
      RECT MASK 2 29.06 87.096 29.12 88.921 ;
      RECT MASK 2 29.33 87.096 29.39 88.921 ;
      RECT MASK 2 29.6 87.096 29.66 88.921 ;
      RECT MASK 2 29.87 87.096 29.93 88.922 ;
      RECT MASK 2 30.182 87.096 30.242 88.922 ;
      RECT MASK 2 30.55 87.096 30.61 88.922 ;
      RECT MASK 2 1.1745 87.19 5.417 87.23 ;
      RECT MASK 2 36.326 87.273 66.476 87.333 ;
      RECT MASK 2 72.716 87.273 102.866 87.333 ;
      RECT MASK 2 8.1745 87.285 12.804 87.405 ;
      RECT MASK 2 13.2225 87.285 17.188 87.405 ;
      RECT MASK 2 17.6065 87.285 24.05 87.405 ;
      RECT MASK 2 1.1745 87.43 5.417 87.47 ;
      RECT MASK 2 1.1745 87.67 5.417 87.71 ;
      RECT MASK 2 8.195 87.705 22.2565 87.885 ;
      RECT MASK 2 5.984 87.72 7.857 87.9 ;
      RECT MASK 2 22.592 87.87 24.05 87.99 ;
      RECT MASK 2 1.1745 87.91 5.417 87.95 ;
      RECT MASK 2 36.326 87.921 36.778 87.981 ;
      RECT MASK 2 37.048 87.921 65.754 87.981 ;
      RECT MASK 2 66.024 87.921 66.476 87.981 ;
      RECT MASK 2 72.716 87.921 73.168 87.981 ;
      RECT MASK 2 73.438 87.921 102.144 87.981 ;
      RECT MASK 2 102.414 87.921 102.866 87.981 ;
      RECT MASK 2 107.4395 87.97 128.5845 88.01 ;
      RECT MASK 2 1.1745 88.15 5.417 88.19 ;
      RECT MASK 2 36.326 88.173 36.778 88.233 ;
      RECT MASK 2 37.048 88.173 65.754 88.233 ;
      RECT MASK 2 66.024 88.173 66.476 88.233 ;
      RECT MASK 2 72.716 88.173 73.168 88.233 ;
      RECT MASK 2 73.438 88.173 102.144 88.233 ;
      RECT MASK 2 102.414 88.173 102.866 88.233 ;
      RECT MASK 2 107.4395 88.21 128.5845 88.25 ;
      RECT MASK 2 22.592 88.29 24.05 88.41 ;
      RECT MASK 2 1.1745 88.39 5.417 88.43 ;
      RECT MASK 2 9.503 88.44 20.9155 88.5 ;
      RECT MASK 2 107.4395 88.45 128.5845 88.49 ;
      RECT MASK 2 8.2595 88.62 16.9585 88.68 ;
      RECT MASK 2 1.1745 88.63 5.417 88.67 ;
      RECT MASK 2 107.4395 88.69 128.5845 88.73 ;
      RECT MASK 2 22.592 88.71 24.05 88.83 ;
      RECT MASK 2 36.326 88.821 66.476 88.881 ;
      RECT MASK 2 72.716 88.821 102.866 88.881 ;
      RECT MASK 2 1.1745 88.87 5.417 88.91 ;
      RECT MASK 2 107.4395 88.93 128.5845 88.97 ;
      RECT MASK 2 8.9875 89.05 9.4645 89.13 ;
      RECT MASK 2 11.4775 89.05 11.9545 89.13 ;
      RECT MASK 2 14.0355 89.05 14.5125 89.13 ;
      RECT MASK 2 15.8615 89.05 16.3385 89.13 ;
      RECT MASK 2 18.4195 89.05 18.8965 89.13 ;
      RECT MASK 2 20.9095 89.05 21.3865 89.13 ;
      RECT MASK 2 36.326 89.073 66.476 89.133 ;
      RECT MASK 2 72.716 89.073 102.866 89.133 ;
      RECT MASK 2 5.984 89.088 7.09 89.268 ;
      RECT MASK 2 1.1745 89.11 5.417 89.15 ;
      RECT MASK 2 22.592 89.13 24.05 89.25 ;
      RECT MASK 2 107.4395 89.17 128.5845 89.21 ;
      RECT MASK 2 8.9875 89.25 9.4645 89.33 ;
      RECT MASK 2 11.4775 89.25 11.9545 89.33 ;
      RECT MASK 2 14.0355 89.25 14.5125 89.33 ;
      RECT MASK 2 15.8615 89.25 16.3385 89.33 ;
      RECT MASK 2 18.4195 89.25 18.8965 89.33 ;
      RECT MASK 2 20.9095 89.25 21.3865 89.33 ;
      RECT MASK 2 1.1745 89.35 5.417 89.39 ;
      RECT MASK 2 107.4395 89.41 128.5845 89.45 ;
      RECT MASK 2 25.68 89.436 25.74 91.262 ;
      RECT MASK 2 26.048 89.436 26.108 91.262 ;
      RECT MASK 2 26.36 89.436 26.42 91.262 ;
      RECT MASK 2 26.63 89.436 26.69 91.261 ;
      RECT MASK 2 26.9 89.436 26.96 91.261 ;
      RECT MASK 2 27.17 89.436 27.23 91.844 ;
      RECT MASK 2 27.44 89.436 27.5 91.844 ;
      RECT MASK 2 27.71 89.436 27.77 91.844 ;
      RECT MASK 2 27.98 89.436 28.04 91.844 ;
      RECT MASK 2 28.25 89.436 28.31 91.844 ;
      RECT MASK 2 28.52 89.436 28.58 91.844 ;
      RECT MASK 2 28.79 89.436 28.85 91.844 ;
      RECT MASK 2 29.06 89.436 29.12 91.844 ;
      RECT MASK 2 29.33 89.436 29.39 91.844 ;
      RECT MASK 2 29.6 89.436 29.66 91.844 ;
      RECT MASK 2 29.87 89.436 29.93 91.844 ;
      RECT MASK 2 30.182 89.436 30.242 91.262 ;
      RECT MASK 2 30.55 89.436 30.61 91.262 ;
      RECT MASK 2 22.592 89.55 24.05 89.67 ;
      RECT MASK 2 1.1745 89.59 5.417 89.63 ;
      RECT MASK 2 8.2595 89.61 16.9585 89.67 ;
      RECT MASK 2 107.4395 89.65 128.5845 89.69 ;
      RECT MASK 2 36.326 89.721 36.778 89.781 ;
      RECT MASK 2 37.048 89.721 65.754 89.781 ;
      RECT MASK 2 66.024 89.721 66.476 89.781 ;
      RECT MASK 2 72.716 89.721 73.168 89.781 ;
      RECT MASK 2 73.438 89.721 102.144 89.781 ;
      RECT MASK 2 102.414 89.721 102.866 89.781 ;
      RECT MASK 2 1.1745 89.83 5.417 89.87 ;
      RECT MASK 2 107.4395 89.89 128.5845 89.93 ;
      RECT MASK 2 22.924 89.97 24.05 90.09 ;
      RECT MASK 2 36.326 89.973 36.778 90.033 ;
      RECT MASK 2 37.048 89.973 65.754 90.033 ;
      RECT MASK 2 66.024 89.973 66.476 90.033 ;
      RECT MASK 2 72.716 89.973 73.168 90.033 ;
      RECT MASK 2 73.438 89.973 102.144 90.033 ;
      RECT MASK 2 102.414 89.973 102.866 90.033 ;
      RECT MASK 2 8.18 90.015 22.2565 90.195 ;
      RECT MASK 2 1.1745 90.07 5.417 90.11 ;
      RECT MASK 2 107.4395 90.13 128.5845 90.17 ;
      RECT MASK 2 1.1745 90.31 5.417 90.35 ;
      RECT MASK 2 107.4395 90.37 128.5845 90.41 ;
      RECT MASK 2 22.924 90.39 24.05 90.51 ;
      RECT MASK 2 8.1745 90.495 12.804 90.615 ;
      RECT MASK 2 13.2225 90.495 17.188 90.615 ;
      RECT MASK 2 17.6065 90.495 22.236 90.615 ;
      RECT MASK 2 1.1745 90.55 5.417 90.59 ;
      RECT MASK 2 107.4395 90.61 128.5845 90.65 ;
      RECT MASK 2 36.326 90.621 66.476 90.681 ;
      RECT MASK 2 72.716 90.621 102.866 90.681 ;
      RECT MASK 2 1.1745 90.79 5.417 90.83 ;
      RECT MASK 2 22.924 90.81 24.05 90.93 ;
      RECT MASK 2 107.4395 90.85 128.5845 90.89 ;
      RECT MASK 2 36.326 90.873 66.476 90.933 ;
      RECT MASK 2 72.716 90.873 102.866 90.933 ;
      RECT MASK 2 7.6395 90.945 12.804 91.065 ;
      RECT MASK 2 13.2225 90.945 17.188 91.065 ;
      RECT MASK 2 17.6065 90.945 22.236 91.065 ;
      RECT MASK 2 1.1745 91.03 5.417 91.07 ;
      RECT MASK 2 107.4395 91.09 128.5845 91.13 ;
      RECT MASK 2 22.924 91.23 24.05 91.35 ;
      RECT MASK 2 1.1745 91.27 5.417 91.31 ;
      RECT MASK 2 107.4395 91.33 128.5845 91.37 ;
      RECT MASK 2 7.66 91.365 22.2565 91.545 ;
      RECT MASK 2 26.36 91.4615 26.42 92.054 ;
      RECT MASK 2 26.63 91.4615 26.69 92.054 ;
      RECT MASK 2 26.9 91.4615 26.96 92.054 ;
      RECT MASK 2 1.1745 91.51 5.417 91.55 ;
      RECT MASK 2 36.326 91.521 36.778 91.581 ;
      RECT MASK 2 37.048 91.521 65.754 91.581 ;
      RECT MASK 2 66.024 91.521 66.476 91.581 ;
      RECT MASK 2 72.716 91.521 73.168 91.581 ;
      RECT MASK 2 73.438 91.521 102.144 91.581 ;
      RECT MASK 2 102.414 91.521 102.866 91.581 ;
      RECT MASK 2 107.4395 91.57 128.5845 91.61 ;
      RECT MASK 2 22.592 91.65 24.05 91.77 ;
      RECT MASK 2 1.1745 91.75 5.417 91.79 ;
      RECT MASK 2 36.326 91.773 36.778 91.833 ;
      RECT MASK 2 37.048 91.773 65.754 91.833 ;
      RECT MASK 2 66.024 91.773 66.476 91.833 ;
      RECT MASK 2 72.716 91.773 73.168 91.833 ;
      RECT MASK 2 73.438 91.773 102.144 91.833 ;
      RECT MASK 2 102.414 91.773 102.866 91.833 ;
      RECT MASK 2 107.4395 91.81 128.5845 91.85 ;
      RECT MASK 2 8.37 91.89 16.2555 91.95 ;
      RECT MASK 2 1.1745 91.99 5.417 92.03 ;
      RECT MASK 2 107.4395 92.05 128.5845 92.09 ;
      RECT MASK 2 22.592 92.07 24.05 92.19 ;
      RECT MASK 2 1.1745 92.23 5.417 92.27 ;
      RECT MASK 2 8.692 92.23 9.4645 92.31 ;
      RECT MASK 2 11.179 92.23 11.9545 92.31 ;
      RECT MASK 2 14.0355 92.23 14.5125 92.31 ;
      RECT MASK 2 15.8615 92.23 16.3385 92.31 ;
      RECT MASK 2 18.4195 92.23 18.8965 92.31 ;
      RECT MASK 2 20.9095 92.23 21.3865 92.31 ;
      RECT MASK 2 107.4395 92.29 128.5845 92.33 ;
      RECT MASK 2 5.984 92.292 7.09 92.472 ;
      RECT MASK 2 36.326 92.421 66.476 92.481 ;
      RECT MASK 2 72.716 92.421 102.866 92.481 ;
      RECT MASK 2 8.692 92.43 9.4645 92.51 ;
      RECT MASK 2 11.179 92.43 11.9545 92.51 ;
      RECT MASK 2 14.0355 92.43 14.5125 92.51 ;
      RECT MASK 2 15.8615 92.43 16.3385 92.51 ;
      RECT MASK 2 18.4195 92.43 18.8965 92.51 ;
      RECT MASK 2 20.9095 92.43 21.3865 92.51 ;
      RECT MASK 2 1.1745 92.47 5.417 92.51 ;
      RECT MASK 2 22.592 92.49 24.05 92.61 ;
      RECT MASK 2 107.4395 92.53 128.5845 92.57 ;
      RECT MASK 2 36.326 92.673 66.476 92.733 ;
      RECT MASK 2 72.716 92.673 102.866 92.733 ;
      RECT MASK 2 1.1745 92.71 5.417 92.75 ;
      RECT MASK 2 107.4395 92.77 128.5845 92.81 ;
      RECT MASK 2 8.37 92.88 16.2555 92.94 ;
      RECT MASK 2 22.592 92.91 24.05 93.03 ;
      RECT MASK 2 1.1745 92.95 5.417 92.99 ;
      RECT MASK 2 107.4395 93.01 128.5845 93.05 ;
      RECT MASK 2 9.2375 93.06 20.9155 93.12 ;
      RECT MASK 2 8.4375 93.1 8.9945 93.16 ;
      RECT MASK 2 1.1745 93.19 5.417 93.23 ;
      RECT MASK 2 107.4395 93.25 128.5845 93.29 ;
      RECT MASK 2 36.326 93.321 36.778 93.381 ;
      RECT MASK 2 37.048 93.321 65.754 93.381 ;
      RECT MASK 2 66.024 93.321 66.476 93.381 ;
      RECT MASK 2 72.716 93.321 73.168 93.381 ;
      RECT MASK 2 73.438 93.321 102.144 93.381 ;
      RECT MASK 2 102.414 93.321 102.866 93.381 ;
      RECT MASK 2 22.592 93.33 24.05 93.45 ;
      RECT MASK 2 1.1745 93.43 5.417 93.47 ;
      RECT MASK 2 107.4395 93.49 128.5845 93.53 ;
      RECT MASK 2 36.326 93.573 36.778 93.633 ;
      RECT MASK 2 37.048 93.573 65.754 93.633 ;
      RECT MASK 2 66.024 93.573 66.476 93.633 ;
      RECT MASK 2 72.716 93.573 73.168 93.633 ;
      RECT MASK 2 73.438 93.573 102.144 93.633 ;
      RECT MASK 2 102.414 93.573 102.866 93.633 ;
      RECT MASK 2 5.984 93.66 7.3325 93.84 ;
      RECT MASK 2 1.1745 93.67 5.417 93.71 ;
      RECT MASK 2 7.66 93.675 24.05 93.855 ;
      RECT MASK 2 107.4395 93.73 128.5845 93.77 ;
      RECT MASK 2 25.237 93.748 31.053 94.134 ;
      RECT MASK 2 1.1745 93.91 5.417 93.95 ;
      RECT MASK 2 107.4395 93.97 128.5845 94.01 ;
      RECT MASK 2 1.1745 94.15 5.417 94.19 ;
      RECT MASK 2 7.6395 94.155 12.804 94.275 ;
      RECT MASK 2 13.2225 94.155 17.188 94.275 ;
      RECT MASK 2 17.6065 94.155 24.05 94.275 ;
      RECT MASK 2 107.4395 94.21 128.5845 94.25 ;
      RECT MASK 2 36.326 94.221 66.476 94.281 ;
      RECT MASK 2 72.716 94.221 102.866 94.281 ;
      RECT MASK 2 1.1745 94.39 5.417 94.43 ;
      RECT MASK 2 107.4395 94.45 128.5845 94.49 ;
      RECT MASK 2 36.326 94.473 66.476 94.533 ;
      RECT MASK 2 72.716 94.473 102.866 94.533 ;
      RECT MASK 2 22.2955 94.59 31.5535 94.71 ;
      RECT MASK 2 1.1745 94.63 5.417 94.67 ;
      RECT MASK 2 107.4395 94.69 128.5845 94.73 ;
      RECT MASK 2 1.1745 94.87 5.417 94.91 ;
      RECT MASK 2 107.4395 94.93 128.5845 94.97 ;
      RECT MASK 2 22.2955 95.01 31.5535 95.13 ;
      RECT MASK 2 1.1745 95.11 5.417 95.15 ;
      RECT MASK 2 107.4395 95.17 128.5845 95.21 ;
      RECT MASK 2 1.1745 95.35 5.417 95.39 ;
      RECT MASK 2 107.4395 95.41 128.5845 95.45 ;
      RECT MASK 2 22.2955 95.43 31.5535 95.55 ;
      RECT MASK 2 1.1745 95.59 5.417 95.63 ;
      RECT MASK 2 107.4395 95.65 128.5845 95.69 ;
      RECT MASK 2 22.2955 95.85 36.7015 95.97 ;
      RECT MASK 2 107.4395 95.89 128.5845 95.93 ;
      RECT MASK 2 107.4395 96.13 128.5845 96.17 ;
      RECT MASK 2 22.2955 96.27 36.7015 96.39 ;
      RECT MASK 2 107.4395 96.37 128.5845 96.41 ;
      RECT MASK 2 1.439 97.75 128.525 97.79 ;
      RECT MASK 2 1.439 97.99 128.525 98.03 ;
      RECT MASK 2 1.439 98.23 128.525 98.27 ;
      RECT MASK 2 1.439 98.47 128.525 98.51 ;
      RECT MASK 2 1.439 98.71 128.525 98.75 ;
      RECT MASK 2 1.439 98.95 128.525 98.99 ;
      RECT MASK 2 1.439 99.19 128.525 99.23 ;
      RECT MASK 2 1.439 99.43 128.525 99.47 ;
      RECT MASK 2 1.439 99.67 128.525 99.71 ;
      RECT MASK 2 1.439 99.91 128.525 99.95 ;
      RECT MASK 2 1.439 100.15 128.525 100.19 ;
      RECT MASK 2 1.439 100.39 128.525 100.43 ;
      RECT MASK 2 1.439 100.63 128.525 100.67 ;
      RECT MASK 2 1.439 100.87 128.525 100.91 ;
      RECT MASK 2 1.439 101.11 128.525 101.15 ;
      RECT MASK 2 1.439 101.35 128.525 101.39 ;
      RECT MASK 2 1.439 101.59 128.525 101.63 ;
      RECT MASK 2 1.439 101.83 128.525 101.87 ;
      RECT MASK 2 1.439 102.07 128.525 102.11 ;
      RECT MASK 2 1.439 102.31 128.525 102.35 ;
      RECT MASK 2 1.439 102.55 128.525 102.59 ;
      RECT MASK 2 1.439 102.79 128.525 102.83 ;
      RECT MASK 2 1.439 103.03 128.525 103.07 ;
      RECT MASK 2 1.439 103.27 128.525 103.31 ;
      RECT MASK 2 1.439 103.51 128.525 103.55 ;
      RECT MASK 2 1.439 103.75 128.525 103.79 ;
      RECT MASK 2 1.439 103.99 128.525 104.03 ;
      RECT MASK 2 1.439 104.23 128.525 104.27 ;
      RECT MASK 2 1.439 104.47 128.525 104.51 ;
      RECT MASK 2 1.439 104.71 128.525 104.75 ;
      RECT MASK 2 1.439 104.95 128.525 104.99 ;
      RECT MASK 2 1.439 105.19 128.525 105.23 ;
      RECT MASK 2 1.439 105.43 128.525 105.47 ;
      RECT MASK 2 1.439 105.67 128.525 105.71 ;
      RECT MASK 2 1.439 105.91 128.525 105.95 ;
      RECT MASK 2 1.439 106.15 128.525 106.19 ;
      RECT MASK 2 1.439 106.39 128.525 106.43 ;
      RECT MASK 2 1.439 106.63 128.525 106.67 ;
      RECT MASK 2 1.439 106.87 128.525 106.91 ;
      RECT MASK 2 1.439 107.11 128.525 107.15 ;
      RECT MASK 2 1.439 107.35 128.525 107.39 ;
      RECT MASK 2 1.439 107.59 128.525 107.63 ;
    LAYER M3 SPACING 0 ;
      RECT MASK 1 41.7465 0.51 41.8665 8.291 ;
      RECT MASK 1 51.0945 0.51 51.1545 1.875 ;
      RECT MASK 1 51.4145 0.51 51.4745 1.875 ;
      RECT MASK 1 52.2335 0.51 52.2935 1.875 ;
      RECT MASK 1 23.8385 0.635 23.8985 3.0695 ;
      RECT MASK 1 22.6385 0.735 22.6985 6.605 ;
      RECT MASK 1 22.8385 0.83 22.8985 4.793 ;
      RECT MASK 1 24.2385 1.035 24.2985 6.655 ;
      RECT MASK 1 23.369 1.235 23.429 3.2145 ;
      RECT MASK 1 63.036 1.299 63.156 3.0225 ;
      RECT MASK 1 64.3005 1.319 64.3805 3.0225 ;
      RECT MASK 1 65.055 1.319 65.135 3.0225 ;
      RECT MASK 1 63.708 1.405 63.768 3.4 ;
      RECT MASK 1 64.086 1.525 64.146 3.28 ;
      RECT MASK 1 3.2225 1.5365 3.2825 9.065 ;
      RECT MASK 1 43.4535 1.5365 43.5135 9.265 ;
      RECT MASK 1 59.676 1.64 59.736 3.04 ;
      RECT MASK 1 62.448 1.64 62.508 3.16 ;
      RECT MASK 1 64.716 1.64 64.776 3.035 ;
      RECT MASK 1 116.428 1.6565 116.488 23.6505 ;
      RECT MASK 1 116.702 1.6565 116.762 23.6505 ;
      RECT MASK 1 116.976 1.6565 117.036 23.6505 ;
      RECT MASK 1 117.25 1.6565 117.31 23.6505 ;
      RECT MASK 1 117.524 1.6565 117.584 23.6505 ;
      RECT MASK 1 117.798 1.6565 117.858 23.6505 ;
      RECT MASK 1 118.072 1.6565 118.132 23.6505 ;
      RECT MASK 1 118.346 1.6565 118.406 23.6505 ;
      RECT MASK 1 118.62 1.6565 118.68 23.6505 ;
      RECT MASK 1 118.894 1.6565 118.954 23.6505 ;
      RECT MASK 1 119.168 1.6565 119.228 23.6505 ;
      RECT MASK 1 119.442 1.6565 119.502 23.6505 ;
      RECT MASK 1 119.716 1.6565 119.776 23.6505 ;
      RECT MASK 1 119.99 1.6565 120.05 23.6505 ;
      RECT MASK 1 120.264 1.6565 120.324 23.6505 ;
      RECT MASK 1 120.538 1.6565 120.598 23.6505 ;
      RECT MASK 1 120.812 1.6565 120.872 23.6505 ;
      RECT MASK 1 121.086 1.6565 121.146 23.6505 ;
      RECT MASK 1 121.36 1.6565 121.42 23.6505 ;
      RECT MASK 1 121.634 1.6565 121.694 23.6505 ;
      RECT MASK 1 121.908 1.6565 121.968 23.6505 ;
      RECT MASK 1 122.182 1.6565 122.242 23.6505 ;
      RECT MASK 1 122.456 1.6565 122.516 23.6505 ;
      RECT MASK 1 122.73 1.6565 122.79 23.6505 ;
      RECT MASK 1 123.004 1.6565 123.064 23.6505 ;
      RECT MASK 1 123.278 1.6565 123.338 23.6505 ;
      RECT MASK 1 123.552 1.6565 123.612 23.6505 ;
      RECT MASK 1 123.826 1.6565 123.886 23.6505 ;
      RECT MASK 1 124.1 1.6565 124.16 23.6505 ;
      RECT MASK 1 124.374 1.6565 124.434 23.6505 ;
      RECT MASK 1 124.648 1.6565 124.708 23.6505 ;
      RECT MASK 1 124.922 1.6565 124.982 23.6505 ;
      RECT MASK 1 125.196 1.6565 125.256 23.6505 ;
      RECT MASK 1 125.47 1.6565 125.53 23.6505 ;
      RECT MASK 1 125.744 1.6565 125.804 23.6505 ;
      RECT MASK 1 126.018 1.6565 126.078 23.6505 ;
      RECT MASK 1 126.292 1.6565 126.352 23.6505 ;
      RECT MASK 1 126.566 1.6565 126.626 23.6505 ;
      RECT MASK 1 126.84 1.6565 126.9 23.6505 ;
      RECT MASK 1 127.114 1.6565 127.174 10.9675 ;
      RECT MASK 1 127.388 1.6565 127.448 10.737 ;
      RECT MASK 1 127.662 1.6565 127.722 10.9675 ;
      RECT MASK 1 127.936 1.6565 127.996 10.962 ;
      RECT MASK 1 47.881 2.4175 47.941 3.044 ;
      RECT MASK 1 46.734 2.4935 46.794 3.965 ;
      RECT MASK 1 59.172 2.72 59.232 3.875 ;
      RECT MASK 1 60.054 2.72 60.114 3.875 ;
      RECT MASK 1 42.4125 2.811 42.4725 9.498 ;
      RECT MASK 1 4.745 2.815 4.805 10.662 ;
      RECT MASK 1 22.04 2.827 22.12 9.0885 ;
      RECT MASK 1 10.1485 3.03 10.2285 6.634 ;
      RECT MASK 1 10.6685 3.03 10.7485 6.634 ;
      RECT MASK 1 56.911 3.1155 57.011 22.36 ;
      RECT MASK 1 57.289 3.1155 57.389 13.815 ;
      RECT MASK 1 57.667 3.1155 57.767 22.36 ;
      RECT MASK 1 60.257 3.1155 60.377 4.6475 ;
      RECT MASK 1 58.045 3.12 58.145 22.36 ;
      RECT MASK 1 58.423 3.12 58.523 16.675 ;
      RECT MASK 1 47.14 3.175 47.2 3.885 ;
      RECT MASK 1 62.336 3.478 62.456 4.6915 ;
      RECT MASK 1 62.6335 3.478 62.7535 4.6915 ;
      RECT MASK 1 63.887 3.4905 64.007 4.636 ;
      RECT MASK 1 64.1915 3.4905 64.3115 4.6515 ;
      RECT MASK 1 59.736 3.537 59.856 4.6475 ;
      RECT MASK 1 63.5435 3.5425 63.6635 4.636 ;
      RECT MASK 1 64.858 3.5425 64.978 4.636 ;
      RECT MASK 1 23.385 3.744 23.485 10.4515 ;
      RECT MASK 1 23.841 3.744 23.901 9.8925 ;
      RECT MASK 1 59.172 4.285 59.232 5.44 ;
      RECT MASK 1 60.054 4.285 60.114 5.44 ;
      RECT MASK 1 5.5115 4.495 5.5715 10.46 ;
      RECT MASK 1 46.34 4.701 46.4 6.413 ;
      RECT MASK 1 63.708 4.76 63.768 6.755 ;
      RECT MASK 1 62.983 4.765 63.043 10.559 ;
      RECT MASK 1 64.086 4.88 64.146 6.635 ;
      RECT MASK 1 62.448 5 62.508 6.52 ;
      RECT MASK 1 46.702 5.04 46.762 9.883 ;
      RECT MASK 1 47.14 5.04 47.2 9.0805 ;
      RECT MASK 1 47.864 5.0405 47.924 8.9845 ;
      RECT MASK 1 59.676 5.12 59.736 6.52 ;
      RECT MASK 1 64.716 5.125 64.776 6.52 ;
      RECT MASK 1 54.1505 5.16 54.2105 11.355 ;
      RECT MASK 1 55.6725 5.16 55.7325 6.573 ;
      RECT MASK 1 63.5265 5.213 63.5865 10.575 ;
      RECT MASK 1 64.299 5.213 64.379 10.575 ;
      RECT MASK 1 65.051 5.213 65.131 10.575 ;
      RECT MASK 1 62.63 5.2165 62.71 10.575 ;
      RECT MASK 1 90.7905 5.5875 90.8505 6.365 ;
      RECT MASK 1 56.0785 6.493 56.1385 11.229 ;
      RECT MASK 1 24.215 6.833 24.275 9.8925 ;
      RECT MASK 1 22.598 6.8415 22.678 10.9305 ;
      RECT MASK 1 22.966 6.8415 23.046 10.9305 ;
      RECT MASK 1 5.105 6.895 5.165 10.561 ;
      RECT MASK 1 63.708 7.645 63.768 9.64 ;
      RECT MASK 1 64.086 7.765 64.146 9.52 ;
      RECT MASK 1 59.676 7.88 59.736 9.28 ;
      RECT MASK 1 62.448 7.88 62.508 9.4 ;
      RECT MASK 1 64.716 7.88 64.776 9.275 ;
      RECT MASK 1 35.8255 8.213 35.8855 9.771 ;
      RECT MASK 1 35.4615 8.314 35.5215 9.498 ;
      RECT MASK 1 54.9065 8.4295 54.9665 9.395 ;
      RECT MASK 1 55.3055 8.4295 55.3655 9.475 ;
      RECT MASK 1 33.123 8.561 33.203 10.1475 ;
      RECT MASK 1 33.501 8.561 33.581 10.1475 ;
      RECT MASK 1 33.879 8.561 33.959 10.1475 ;
      RECT MASK 1 34.276 8.561 34.356 10.1475 ;
      RECT MASK 1 34.663 8.561 34.743 10.1475 ;
      RECT MASK 1 52.892 8.7785 52.952 11.229 ;
      RECT MASK 1 44.073 8.9145 44.133 10.353 ;
      RECT MASK 1 59.172 8.96 59.232 10.115 ;
      RECT MASK 1 60.054 8.96 60.114 10.115 ;
      RECT MASK 1 4.359 8.995 4.419 10.763 ;
      RECT MASK 1 44.451 9.0105 44.511 10.749 ;
      RECT MASK 1 31.0965 9.583 31.1565 10.5725 ;
      RECT MASK 1 56.511 9.7745 56.571 11.133 ;
      RECT MASK 1 31.418 9.785 31.478 10.7745 ;
      RECT MASK 1 58.801 10.22 58.901 16.662 ;
      RECT MASK 1 59.571 10.22 59.671 14.72 ;
      RECT MASK 1 60.743 10.229 60.823 14.75 ;
      RECT MASK 1 23.824 10.2455 23.924 87.62 ;
      RECT MASK 1 31.9245 10.6455 31.9845 11.12 ;
      RECT MASK 1 59.179 10.745 59.279 17.646 ;
      RECT MASK 1 59.963 10.745 60.083 16.66 ;
      RECT MASK 1 61.135 10.745 61.215 16.7365 ;
      RECT MASK 1 61.513 10.745 61.593 17.646 ;
      RECT MASK 1 61.891 10.745 61.971 14.75 ;
      RECT MASK 1 62.297 10.745 62.377 16.687 ;
      RECT MASK 1 63.539 10.745 63.619 17.646 ;
      RECT MASK 1 63.917 10.745 63.997 17.646 ;
      RECT MASK 1 64.673 10.745 64.753 17.646 ;
      RECT MASK 1 65.429 10.745 65.509 13.821 ;
      RECT MASK 1 65.807 10.745 65.887 13.821 ;
      RECT MASK 1 66.213 10.745 66.293 13.821 ;
      RECT MASK 1 66.591 10.745 66.671 13.821 ;
      RECT MASK 1 66.969 10.745 67.049 13.821 ;
      RECT MASK 1 67.347 10.745 67.427 13.821 ;
      RECT MASK 1 67.753 10.745 67.833 13.821 ;
      RECT MASK 1 68.131 10.745 68.211 13.821 ;
      RECT MASK 1 68.528 10.745 68.608 13.821 ;
      RECT MASK 1 68.915 10.745 68.995 13.821 ;
      RECT MASK 1 69.293 10.745 69.373 13.821 ;
      RECT MASK 1 69.7355 10.745 69.8155 13.821 ;
      RECT MASK 1 70.157 10.745 70.237 13.821 ;
      RECT MASK 1 70.535 10.745 70.615 13.821 ;
      RECT MASK 1 70.913 10.745 70.993 13.821 ;
      RECT MASK 1 71.291 10.745 71.371 13.821 ;
      RECT MASK 1 23.418 10.8535 23.518 87.17 ;
      RECT MASK 1 24.199 10.9275 24.299 94.04 ;
      RECT MASK 1 24.955 11.1105 25.055 85.786 ;
      RECT MASK 1 127.138 11.159 127.258 27.755 ;
      RECT MASK 1 127.578 11.218 127.698 80.021 ;
      RECT MASK 1 22.589 11.354 22.669 14.777 ;
      RECT MASK 1 22.967 11.354 23.047 14.777 ;
      RECT MASK 1 24.587 11.354 24.667 14.777 ;
      RECT MASK 1 25.343 11.354 25.423 14.777 ;
      RECT MASK 1 25.721 11.354 25.801 14.777 ;
      RECT MASK 1 26.099 11.354 26.179 14.777 ;
      RECT MASK 1 26.505 11.354 26.585 14.777 ;
      RECT MASK 1 26.883 11.354 26.963 14.777 ;
      RECT MASK 1 27.261 11.354 27.341 13.773 ;
      RECT MASK 1 27.667 11.354 27.747 14.777 ;
      RECT MASK 1 28.045 11.354 28.125 14.777 ;
      RECT MASK 1 28.423 11.354 28.503 14.783 ;
      RECT MASK 1 56.533 11.384 56.633 22.36 ;
      RECT MASK 1 38.579 11.566 38.659 14.766 ;
      RECT MASK 1 38.957 11.566 39.037 14.766 ;
      RECT MASK 1 39.335 11.566 39.415 14.766 ;
      RECT MASK 1 39.741 11.566 39.821 14.766 ;
      RECT MASK 1 40.119 11.566 40.199 14.766 ;
      RECT MASK 1 40.516 11.566 40.596 13.818 ;
      RECT MASK 1 40.892 11.566 40.972 14.766 ;
      RECT MASK 1 41.318 11.566 41.398 14.766 ;
      RECT MASK 1 41.715 11.566 41.795 14.766 ;
      RECT MASK 1 42.065 11.566 42.145 14.766 ;
      RECT MASK 1 42.443 11.566 42.523 14.766 ;
      RECT MASK 1 42.84 11.566 42.92 14.766 ;
      RECT MASK 1 43.24 11.566 43.32 14.766 ;
      RECT MASK 1 43.685 11.566 43.765 13.771 ;
      RECT MASK 1 44.063 11.566 44.143 14.766 ;
      RECT MASK 1 44.441 11.566 44.521 14.766 ;
      RECT MASK 1 44.819 11.566 44.899 14.766 ;
      RECT MASK 1 45.197 11.566 45.277 14.766 ;
      RECT MASK 1 45.575 11.566 45.655 14.766 ;
      RECT MASK 1 45.953 11.566 46.033 14.766 ;
      RECT MASK 1 46.345 11.566 46.425 14.766 ;
      RECT MASK 1 46.737 11.566 46.817 14.766 ;
      RECT MASK 1 47.115 11.566 47.195 14.766 ;
      RECT MASK 1 47.493 11.566 47.573 14.766 ;
      RECT MASK 1 47.899 11.566 47.979 14.766 ;
      RECT MASK 1 48.277 11.566 48.357 14.766 ;
      RECT MASK 1 48.683 11.566 48.763 14.766 ;
      RECT MASK 1 49.061 11.566 49.141 14.766 ;
      RECT MASK 1 49.439 11.566 49.519 14.766 ;
      RECT MASK 1 49.861 11.566 49.941 14.766 ;
      RECT MASK 1 50.303 11.566 50.383 14.766 ;
      RECT MASK 1 50.681 11.566 50.761 12.857 ;
      RECT MASK 1 51.059 11.566 51.139 14.766 ;
      RECT MASK 1 51.437 11.566 51.517 14.766 ;
      RECT MASK 1 51.815 11.566 51.895 14.766 ;
      RECT MASK 1 52.193 11.566 52.273 14.766 ;
      RECT MASK 1 52.608 11.566 52.688 14.766 ;
      RECT MASK 1 53.754 11.566 53.834 13.836 ;
      RECT MASK 1 54.52 11.566 54.6 14.766 ;
      RECT MASK 1 54.894 11.566 54.974 14.766 ;
      RECT MASK 1 55.302 11.566 55.382 14.766 ;
      RECT MASK 1 55.663 11.566 55.743 14.766 ;
      RECT MASK 1 90.936 11.67 91.056 14.4945 ;
      RECT MASK 1 108.008 11.67 108.128 14.322 ;
      RECT MASK 1 56.058 11.68 56.138 14.766 ;
      RECT MASK 1 54.144 11.685 54.224 14.766 ;
      RECT MASK 1 62.675 11.74 62.755 17.646 ;
      RECT MASK 1 63.161 11.74 63.241 17.646 ;
      RECT MASK 1 64.295 11.74 64.375 14.75 ;
      RECT MASK 1 65.051 11.74 65.131 16.687 ;
      RECT MASK 1 60.351 11.76 60.431 12.72 ;
      RECT MASK 1 38.181 12.848 38.241 14.458 ;
      RECT MASK 1 53.299 12.848 53.359 16.378 ;
      RECT MASK 1 60.305 12.848 60.365 16.378 ;
      RECT MASK 1 50.789 13.136 50.849 14.848 ;
      RECT MASK 1 83.117 13.136 83.177 16.768 ;
      RECT MASK 1 66.959 14.089 67.059 17.82 ;
      RECT MASK 1 17.191 14.576 17.251 16.768 ;
      RECT MASK 1 30.631 14.576 30.691 16.768 ;
      RECT MASK 1 43.831 14.576 43.891 16.768 ;
      RECT MASK 1 57.317 14.576 57.377 16.768 ;
      RECT MASK 1 70.517 14.576 70.577 16.768 ;
      RECT MASK 1 83.837 14.576 83.897 16.768 ;
      RECT MASK 1 97.157 14.576 97.217 16.768 ;
      RECT MASK 1 95.813 14.672 95.873 16.768 ;
      RECT MASK 1 107.969 14.672 108.029 16.768 ;
      RECT MASK 1 27.2785 14.768 27.3385 16.768 ;
      RECT MASK 1 40.5215 14.768 40.5815 16.768 ;
      RECT MASK 1 53.817 14.768 53.877 16.768 ;
      RECT MASK 1 80.575 14.768 80.635 16.768 ;
      RECT MASK 1 82.097 14.864 82.157 16.768 ;
      RECT MASK 1 6.641 15.05 6.741 83.684 ;
      RECT MASK 1 7.803 15.05 7.903 83.684 ;
      RECT MASK 1 8.965 15.05 9.065 83.684 ;
      RECT MASK 1 11.747 15.05 11.807 17.434 ;
      RECT MASK 1 13.259 15.05 13.359 83.684 ;
      RECT MASK 1 14.421 15.05 14.521 83.684 ;
      RECT MASK 1 15.583 15.05 15.683 83.684 ;
      RECT MASK 1 18.271 15.05 18.331 17.434 ;
      RECT MASK 1 19.877 15.05 19.977 83.684 ;
      RECT MASK 1 21.039 15.05 21.139 83.684 ;
      RECT MASK 1 22.201 15.05 22.301 83.684 ;
      RECT MASK 1 24.585 15.05 24.645 17.434 ;
      RECT MASK 1 26.495 15.05 26.595 83.684 ;
      RECT MASK 1 27.657 15.05 27.757 83.684 ;
      RECT MASK 1 28.819 15.05 28.919 83.684 ;
      RECT MASK 1 33.113 15.05 33.213 83.684 ;
      RECT MASK 1 34.275 15.05 34.375 83.684 ;
      RECT MASK 1 35.437 15.05 35.537 83.684 ;
      RECT MASK 1 37.591 15.05 37.651 17.434 ;
      RECT MASK 1 39.731 15.05 39.831 83.684 ;
      RECT MASK 1 40.893 15.05 40.993 83.684 ;
      RECT MASK 1 42.055 15.05 42.155 83.684 ;
      RECT MASK 1 46.349 15.05 46.449 83.684 ;
      RECT MASK 1 47.511 15.05 47.611 83.684 ;
      RECT MASK 1 48.673 15.05 48.773 83.684 ;
      RECT MASK 1 51.029 15.05 51.089 17.434 ;
      RECT MASK 1 52.183 15.05 52.283 20.54 ;
      RECT MASK 1 54.129 15.05 54.229 83.684 ;
      RECT MASK 1 55.291 15.05 55.391 83.684 ;
      RECT MASK 1 59.585 15.05 59.685 83.684 ;
      RECT MASK 1 60.747 15.05 60.847 83.684 ;
      RECT MASK 1 61.909 15.05 62.009 83.684 ;
      RECT MASK 1 64.339 15.05 64.399 17.434 ;
      RECT MASK 1 66.203 15.05 66.303 83.684 ;
      RECT MASK 1 67.365 15.05 67.465 83.684 ;
      RECT MASK 1 68.527 15.05 68.627 83.684 ;
      RECT MASK 1 72.821 15.05 72.921 83.684 ;
      RECT MASK 1 73.983 15.05 74.083 83.684 ;
      RECT MASK 1 75.145 15.05 75.245 83.684 ;
      RECT MASK 1 79.439 15.05 79.539 83.684 ;
      RECT MASK 1 81.763 15.05 81.863 83.684 ;
      RECT MASK 1 84.077 15.05 84.137 17.434 ;
      RECT MASK 1 86.057 15.05 86.157 83.684 ;
      RECT MASK 1 87.219 15.05 87.319 83.684 ;
      RECT MASK 1 88.381 15.05 88.481 83.684 ;
      RECT MASK 1 90.917 15.05 90.977 17.434 ;
      RECT MASK 1 92.675 15.05 92.775 83.684 ;
      RECT MASK 1 93.837 15.05 93.937 83.684 ;
      RECT MASK 1 94.999 15.05 95.099 83.684 ;
      RECT MASK 1 99.293 15.05 99.393 83.684 ;
      RECT MASK 1 100.455 15.05 100.555 83.684 ;
      RECT MASK 1 101.617 15.05 101.717 83.684 ;
      RECT MASK 1 105.911 15.05 106.011 83.684 ;
      RECT MASK 1 107.073 15.05 107.173 83.684 ;
      RECT MASK 1 108.235 15.05 108.335 83.684 ;
      RECT MASK 1 65.807 16.2105 65.887 18.1395 ;
      RECT MASK 1 5.857 16.976 5.957 20.54 ;
      RECT MASK 1 7.019 16.976 7.119 20.54 ;
      RECT MASK 1 8.181 16.976 8.281 20.54 ;
      RECT MASK 1 12.475 16.976 12.575 20.54 ;
      RECT MASK 1 13.637 16.976 13.737 20.54 ;
      RECT MASK 1 14.799 16.976 14.899 20.54 ;
      RECT MASK 1 19.093 16.976 19.193 20.54 ;
      RECT MASK 1 20.255 16.976 20.355 20.54 ;
      RECT MASK 1 25.711 16.976 25.811 20.54 ;
      RECT MASK 1 26.873 16.976 26.973 20.54 ;
      RECT MASK 1 28.035 16.976 28.135 20.54 ;
      RECT MASK 1 32.329 16.976 32.429 20.54 ;
      RECT MASK 1 33.491 16.976 33.591 20.54 ;
      RECT MASK 1 34.653 16.976 34.753 20.54 ;
      RECT MASK 1 38.947 16.976 39.047 20.54 ;
      RECT MASK 1 40.109 16.976 40.209 20.54 ;
      RECT MASK 1 41.271 16.976 41.371 20.54 ;
      RECT MASK 1 45.565 16.976 45.665 20.54 ;
      RECT MASK 1 46.727 16.976 46.827 20.54 ;
      RECT MASK 1 47.889 16.976 47.989 20.54 ;
      RECT MASK 1 52.967 16.976 53.067 83.684 ;
      RECT MASK 1 53.345 16.976 53.445 20.54 ;
      RECT MASK 1 54.507 16.976 54.607 20.54 ;
      RECT MASK 1 58.801 16.976 58.901 20.54 ;
      RECT MASK 1 59.963 16.976 60.063 20.54 ;
      RECT MASK 1 61.125 16.976 61.225 20.54 ;
      RECT MASK 1 65.419 16.976 65.519 20.54 ;
      RECT MASK 1 66.581 16.976 66.681 20.54 ;
      RECT MASK 1 67.743 16.976 67.843 20.54 ;
      RECT MASK 1 72.037 16.976 72.137 20.54 ;
      RECT MASK 1 73.199 16.976 73.299 20.54 ;
      RECT MASK 1 74.361 16.976 74.461 20.54 ;
      RECT MASK 1 78.655 16.976 78.755 20.54 ;
      RECT MASK 1 79.817 16.976 79.917 20.54 ;
      RECT MASK 1 85.273 16.976 85.373 20.54 ;
      RECT MASK 1 86.435 16.976 86.535 20.54 ;
      RECT MASK 1 87.597 16.976 87.697 20.54 ;
      RECT MASK 1 91.891 16.976 91.991 20.54 ;
      RECT MASK 1 93.053 16.976 93.153 20.54 ;
      RECT MASK 1 94.215 16.976 94.315 20.54 ;
      RECT MASK 1 98.509 16.976 98.609 20.54 ;
      RECT MASK 1 99.671 16.976 99.771 20.54 ;
      RECT MASK 1 100.833 16.976 100.933 20.54 ;
      RECT MASK 1 105.127 16.976 105.227 20.54 ;
      RECT MASK 1 106.289 16.976 106.389 20.54 ;
      RECT MASK 1 107.451 16.976 107.551 20.54 ;
      RECT MASK 1 9.343 17.354 9.443 20.54 ;
      RECT MASK 1 12.097 17.354 12.197 83.684 ;
      RECT MASK 1 15.961 17.354 16.061 20.54 ;
      RECT MASK 1 18.715 17.354 18.815 83.684 ;
      RECT MASK 1 21.417 17.354 21.517 20.54 ;
      RECT MASK 1 22.579 17.354 22.679 20.54 ;
      RECT MASK 1 25.333 17.354 25.433 83.684 ;
      RECT MASK 1 29.197 17.354 29.297 20.54 ;
      RECT MASK 1 31.951 17.354 32.051 83.684 ;
      RECT MASK 1 35.815 17.354 35.915 20.54 ;
      RECT MASK 1 38.569 17.354 38.669 83.684 ;
      RECT MASK 1 42.433 17.354 42.533 20.54 ;
      RECT MASK 1 45.187 17.354 45.287 83.684 ;
      RECT MASK 1 49.051 17.354 49.151 20.54 ;
      RECT MASK 1 51.805 17.354 51.905 83.684 ;
      RECT MASK 1 55.669 17.354 55.769 20.54 ;
      RECT MASK 1 58.423 17.354 58.523 83.684 ;
      RECT MASK 1 62.287 17.354 62.387 20.54 ;
      RECT MASK 1 65.041 17.354 65.141 83.684 ;
      RECT MASK 1 68.905 17.354 69.005 20.54 ;
      RECT MASK 1 71.659 17.354 71.759 83.684 ;
      RECT MASK 1 75.523 17.354 75.623 20.54 ;
      RECT MASK 1 78.277 17.354 78.377 83.684 ;
      RECT MASK 1 80.601 17.354 80.701 83.684 ;
      RECT MASK 1 82.141 17.354 82.241 20.54 ;
      RECT MASK 1 84.895 17.354 84.995 83.684 ;
      RECT MASK 1 88.759 17.354 88.859 20.54 ;
      RECT MASK 1 91.513 17.354 91.613 83.684 ;
      RECT MASK 1 95.377 17.354 95.477 20.54 ;
      RECT MASK 1 98.131 17.354 98.231 83.684 ;
      RECT MASK 1 101.995 17.354 102.095 20.54 ;
      RECT MASK 1 104.749 17.354 104.849 83.684 ;
      RECT MASK 1 108.613 17.354 108.713 20.54 ;
      RECT MASK 1 57.289 17.4475 57.389 22.36 ;
      RECT MASK 1 80.979 17.458 81.079 20.54 ;
      RECT MASK 1 2.499 19.63 2.559 24.53 ;
      RECT MASK 1 2.773 19.63 2.833 24.53 ;
      RECT MASK 1 3.047 19.63 3.107 24.53 ;
      RECT MASK 1 3.321 19.63 3.381 24.53 ;
      RECT MASK 1 3.595 19.63 3.655 24.53 ;
      RECT MASK 1 59.179 20.4 59.279 21.679 ;
      RECT MASK 1 60.341 20.4 60.441 21.679 ;
      RECT MASK 1 58.801 20.8 58.901 21.935 ;
      RECT MASK 1 59.963 20.8 60.063 21.92 ;
      RECT MASK 1 7.387 22.0925 7.507 81.8875 ;
      RECT MASK 1 8.549 22.0925 8.669 81.8875 ;
      RECT MASK 1 9.711 22.0925 9.831 81.8875 ;
      RECT MASK 1 12.843 22.0925 12.963 81.8875 ;
      RECT MASK 1 14.005 22.0925 14.125 81.8875 ;
      RECT MASK 1 15.167 22.0925 15.287 81.8875 ;
      RECT MASK 1 16.329 22.0925 16.449 81.8875 ;
      RECT MASK 1 19.461 22.0925 19.581 81.8875 ;
      RECT MASK 1 20.623 22.0925 20.743 81.8875 ;
      RECT MASK 1 21.785 22.0925 21.905 81.8875 ;
      RECT MASK 1 22.947 22.0925 23.067 81.8875 ;
      RECT MASK 1 26.079 22.0925 26.199 81.8875 ;
      RECT MASK 1 27.241 22.0925 27.361 81.8875 ;
      RECT MASK 1 28.403 22.0925 28.523 81.8875 ;
      RECT MASK 1 29.565 22.0925 29.685 81.8875 ;
      RECT MASK 1 32.697 22.0925 32.817 81.8875 ;
      RECT MASK 1 33.859 22.0925 33.979 81.8875 ;
      RECT MASK 1 35.021 22.0925 35.141 81.8875 ;
      RECT MASK 1 36.183 22.0925 36.303 81.8875 ;
      RECT MASK 1 39.315 22.0925 39.435 81.8875 ;
      RECT MASK 1 40.477 22.0925 40.597 81.8875 ;
      RECT MASK 1 41.639 22.0925 41.759 81.8875 ;
      RECT MASK 1 42.801 22.0925 42.921 81.8875 ;
      RECT MASK 1 45.933 22.0925 46.053 81.8875 ;
      RECT MASK 1 47.095 22.0925 47.215 81.8875 ;
      RECT MASK 1 48.257 22.0925 48.377 81.8875 ;
      RECT MASK 1 49.419 22.0925 49.539 81.8875 ;
      RECT MASK 1 52.551 22.0925 52.671 81.8875 ;
      RECT MASK 1 53.713 22.0925 53.833 81.8875 ;
      RECT MASK 1 54.875 22.0925 54.995 81.8875 ;
      RECT MASK 1 56.037 22.0925 56.157 81.8875 ;
      RECT MASK 1 60.331 22.0925 60.451 81.8875 ;
      RECT MASK 1 61.493 22.0925 61.613 81.8875 ;
      RECT MASK 1 62.655 22.0925 62.775 81.8875 ;
      RECT MASK 1 65.787 22.0925 65.907 81.8875 ;
      RECT MASK 1 66.949 22.0925 67.069 81.8875 ;
      RECT MASK 1 68.111 22.0925 68.231 81.8875 ;
      RECT MASK 1 69.273 22.0925 69.393 81.8875 ;
      RECT MASK 1 72.405 22.0925 72.525 81.8875 ;
      RECT MASK 1 73.567 22.0925 73.687 81.8875 ;
      RECT MASK 1 74.729 22.0925 74.849 81.8875 ;
      RECT MASK 1 75.891 22.0925 76.011 81.8875 ;
      RECT MASK 1 79.023 22.0925 79.143 81.8875 ;
      RECT MASK 1 80.185 22.0925 80.305 81.8875 ;
      RECT MASK 1 81.347 22.0925 81.467 81.8875 ;
      RECT MASK 1 82.509 22.0925 82.629 81.8875 ;
      RECT MASK 1 85.641 22.0925 85.761 81.8875 ;
      RECT MASK 1 86.803 22.0925 86.923 81.8875 ;
      RECT MASK 1 87.965 22.0925 88.085 81.8875 ;
      RECT MASK 1 89.127 22.0925 89.247 81.8875 ;
      RECT MASK 1 92.259 22.0925 92.379 81.8875 ;
      RECT MASK 1 93.421 22.0925 93.541 81.8875 ;
      RECT MASK 1 94.583 22.0925 94.703 81.8875 ;
      RECT MASK 1 95.745 22.0925 95.865 81.8875 ;
      RECT MASK 1 98.877 22.0925 98.997 81.8875 ;
      RECT MASK 1 100.039 22.0925 100.159 81.8875 ;
      RECT MASK 1 101.201 22.0925 101.321 81.8875 ;
      RECT MASK 1 102.363 22.0925 102.483 81.8875 ;
      RECT MASK 1 105.495 22.0925 105.615 81.8875 ;
      RECT MASK 1 106.657 22.0925 106.777 81.8875 ;
      RECT MASK 1 107.819 22.0925 107.939 81.8875 ;
      RECT MASK 1 108.981 22.0925 109.101 81.8875 ;
      RECT MASK 1 6.225 22.1225 6.345 25.733 ;
      RECT MASK 1 59.169 22.1225 59.289 81.8875 ;
      RECT MASK 1 5.847 22.234 5.967 57.4415 ;
      RECT MASK 1 7.009 22.234 7.129 51.36 ;
      RECT MASK 1 8.171 22.234 8.291 45.0215 ;
      RECT MASK 1 9.333 22.234 9.453 39.08 ;
      RECT MASK 1 12.465 22.234 12.585 32.729 ;
      RECT MASK 1 13.627 22.234 13.747 39.08 ;
      RECT MASK 1 14.789 22.234 14.909 45.0215 ;
      RECT MASK 1 15.951 22.234 16.071 51.36 ;
      RECT MASK 1 19.083 22.234 19.203 51.4115 ;
      RECT MASK 1 20.245 22.234 20.365 51.36 ;
      RECT MASK 1 21.407 22.234 21.527 45.0215 ;
      RECT MASK 1 22.569 22.234 22.689 39.08 ;
      RECT MASK 1 25.701 22.234 25.821 32.8415 ;
      RECT MASK 1 26.863 22.234 26.983 39.08 ;
      RECT MASK 1 28.025 22.234 28.145 45.0215 ;
      RECT MASK 1 29.187 22.234 29.307 51.36 ;
      RECT MASK 1 32.319 22.234 32.439 51.4115 ;
      RECT MASK 1 33.481 22.234 33.601 51.36 ;
      RECT MASK 1 34.643 22.234 34.763 45.0215 ;
      RECT MASK 1 35.805 22.234 35.925 39.08 ;
      RECT MASK 1 38.937 22.234 39.057 32.8415 ;
      RECT MASK 1 40.099 22.234 40.219 39.08 ;
      RECT MASK 1 41.261 22.234 41.381 45.0215 ;
      RECT MASK 1 42.423 22.234 42.543 51.36 ;
      RECT MASK 1 45.555 22.234 45.675 51.4115 ;
      RECT MASK 1 46.717 22.234 46.837 51.36 ;
      RECT MASK 1 47.879 22.234 47.999 45.0215 ;
      RECT MASK 1 49.041 22.234 49.161 39.08 ;
      RECT MASK 1 52.173 22.234 52.293 32.8415 ;
      RECT MASK 1 53.335 22.234 53.455 39.08 ;
      RECT MASK 1 54.497 22.234 54.617 45.0215 ;
      RECT MASK 1 55.659 22.234 55.779 51.36 ;
      RECT MASK 1 58.791 22.234 58.911 51.4115 ;
      RECT MASK 1 59.953 22.234 60.073 51.36 ;
      RECT MASK 1 61.115 22.234 61.235 45.0215 ;
      RECT MASK 1 62.277 22.234 62.397 39.08 ;
      RECT MASK 1 65.409 22.234 65.529 32.8415 ;
      RECT MASK 1 66.571 22.234 66.691 39.08 ;
      RECT MASK 1 67.733 22.234 67.853 45.0215 ;
      RECT MASK 1 68.895 22.234 69.015 51.36 ;
      RECT MASK 1 72.027 22.234 72.147 51.4115 ;
      RECT MASK 1 73.189 22.234 73.309 51.36 ;
      RECT MASK 1 74.351 22.234 74.471 45.0215 ;
      RECT MASK 1 75.513 22.234 75.633 39.08 ;
      RECT MASK 1 78.645 22.234 78.765 33.0815 ;
      RECT MASK 1 79.807 22.234 79.927 39.08 ;
      RECT MASK 1 80.969 22.234 81.089 45.0215 ;
      RECT MASK 1 82.131 22.234 82.251 51.36 ;
      RECT MASK 1 85.263 22.234 85.383 51.4115 ;
      RECT MASK 1 86.425 22.234 86.545 51.36 ;
      RECT MASK 1 87.587 22.234 87.707 45.0215 ;
      RECT MASK 1 88.749 22.234 88.869 39.08 ;
      RECT MASK 1 91.881 22.234 92.001 33.0815 ;
      RECT MASK 1 93.043 22.234 93.163 39.08 ;
      RECT MASK 1 94.205 22.234 94.325 45.0215 ;
      RECT MASK 1 95.367 22.234 95.487 51.6 ;
      RECT MASK 1 98.499 22.234 98.619 51.4115 ;
      RECT MASK 1 99.661 22.234 99.781 51.36 ;
      RECT MASK 1 100.823 22.234 100.943 45.0215 ;
      RECT MASK 1 101.985 22.234 102.105 39.08 ;
      RECT MASK 1 105.117 22.234 105.237 32.8415 ;
      RECT MASK 1 106.279 22.234 106.399 39.08 ;
      RECT MASK 1 107.441 22.234 107.561 45.0815 ;
      RECT MASK 1 108.603 22.234 108.723 51.45 ;
      RECT MASK 1 1.417 26.1 1.537 77.69 ;
      RECT MASK 1 2.173 26.1 2.293 77.69 ;
      RECT MASK 1 2.929 26.1 3.049 77.69 ;
      RECT MASK 1 3.685 26.1 3.805 77.69 ;
      RECT MASK 1 4.441 26.1 4.561 77.69 ;
      RECT MASK 1 116.323 26.4785 116.463 28.18 ;
      RECT MASK 1 117.079 26.4785 117.219 28.18 ;
      RECT MASK 1 117.835 26.4785 117.975 28.18 ;
      RECT MASK 1 118.591 26.4785 118.731 28.18 ;
      RECT MASK 1 119.347 26.4785 119.487 28.18 ;
      RECT MASK 1 120.103 26.4785 120.243 28.18 ;
      RECT MASK 1 120.859 26.4785 120.999 28.18 ;
      RECT MASK 1 121.615 26.4785 121.755 28.18 ;
      RECT MASK 1 122.371 26.4785 122.511 28.18 ;
      RECT MASK 1 123.127 26.4785 123.267 28.18 ;
      RECT MASK 1 123.883 26.4785 124.023 28.18 ;
      RECT MASK 1 124.639 26.4785 124.779 28.18 ;
      RECT MASK 1 125.395 26.4785 125.535 28.18 ;
      RECT MASK 1 126.151 26.4785 126.291 28.18 ;
      RECT MASK 1 117.457 26.94 117.597 51.3195 ;
      RECT MASK 1 118.213 26.94 118.353 51.3195 ;
      RECT MASK 1 118.969 26.94 119.109 51.3195 ;
      RECT MASK 1 119.725 26.94 119.865 51.3195 ;
      RECT MASK 1 120.481 26.94 120.621 51.3195 ;
      RECT MASK 1 121.237 26.94 121.377 51.3195 ;
      RECT MASK 1 121.993 26.94 122.133 51.3195 ;
      RECT MASK 1 122.749 26.94 122.889 51.3195 ;
      RECT MASK 1 123.505 26.94 123.645 51.3195 ;
      RECT MASK 1 124.261 26.94 124.401 51.3195 ;
      RECT MASK 1 125.017 26.94 125.157 51.3195 ;
      RECT MASK 1 125.773 26.94 125.913 51.3195 ;
      RECT MASK 1 123.883 28.683 124.023 51.3195 ;
      RECT MASK 1 116.323 28.7505 116.463 51.3195 ;
      RECT MASK 1 117.835 28.7505 117.975 51.3195 ;
      RECT MASK 1 118.591 28.7505 118.731 51.3195 ;
      RECT MASK 1 119.347 28.7505 119.487 51.3195 ;
      RECT MASK 1 120.103 28.7505 120.243 51.3195 ;
      RECT MASK 1 120.859 28.7505 120.999 51.3195 ;
      RECT MASK 1 121.615 28.7505 121.755 51.3195 ;
      RECT MASK 1 122.371 28.7505 122.511 51.3195 ;
      RECT MASK 1 123.127 28.7505 123.267 51.3195 ;
      RECT MASK 1 124.639 28.7505 124.779 51.3195 ;
      RECT MASK 1 125.395 28.7505 125.535 51.3195 ;
      RECT MASK 1 126.151 28.7505 126.291 51.3195 ;
      RECT MASK 1 117.079 28.7615 117.219 51.3195 ;
      RECT MASK 1 126.913 30.141 127.033 72.484 ;
      RECT MASK 1 7.009 52.2685 7.129 81.746 ;
      RECT MASK 1 15.951 52.2685 16.071 81.746 ;
      RECT MASK 1 20.245 52.2685 20.365 81.746 ;
      RECT MASK 1 29.187 52.2685 29.307 81.746 ;
      RECT MASK 1 33.481 52.2685 33.601 81.746 ;
      RECT MASK 1 42.423 52.2685 42.543 81.746 ;
      RECT MASK 1 46.717 52.2685 46.837 81.746 ;
      RECT MASK 1 55.659 52.2685 55.779 81.746 ;
      RECT MASK 1 59.953 52.2685 60.073 81.746 ;
      RECT MASK 1 68.895 52.2685 69.015 81.746 ;
      RECT MASK 1 73.189 52.2685 73.309 81.746 ;
      RECT MASK 1 82.131 52.2685 82.251 81.746 ;
      RECT MASK 1 86.425 52.2685 86.545 81.746 ;
      RECT MASK 1 95.367 52.2685 95.487 81.746 ;
      RECT MASK 1 99.661 52.2685 99.781 81.746 ;
      RECT MASK 1 108.603 52.5085 108.723 81.746 ;
      RECT MASK 1 19.083 52.6215 19.203 81.746 ;
      RECT MASK 1 32.319 52.6215 32.439 81.746 ;
      RECT MASK 1 45.555 52.6215 45.675 81.746 ;
      RECT MASK 1 58.791 52.6215 58.911 81.746 ;
      RECT MASK 1 72.027 52.6215 72.147 81.746 ;
      RECT MASK 1 85.263 52.6215 85.383 81.746 ;
      RECT MASK 1 98.499 52.6215 98.619 81.746 ;
      RECT MASK 1 116.323 52.687 116.463 76.57 ;
      RECT MASK 1 117.318 52.687 117.358 69.9575 ;
      RECT MASK 1 117.696 52.687 117.736 69.9575 ;
      RECT MASK 1 118.074 52.687 118.114 69.9575 ;
      RECT MASK 1 118.452 52.687 118.492 69.9575 ;
      RECT MASK 1 118.83 52.687 118.87 69.9575 ;
      RECT MASK 1 119.208 52.687 119.248 69.9575 ;
      RECT MASK 1 119.586 52.687 119.626 69.9575 ;
      RECT MASK 1 119.964 52.687 120.004 69.9575 ;
      RECT MASK 1 120.342 52.687 120.382 69.9575 ;
      RECT MASK 1 120.72 52.687 120.76 69.9575 ;
      RECT MASK 1 121.098 52.687 121.138 69.9575 ;
      RECT MASK 1 121.476 52.687 121.516 69.9575 ;
      RECT MASK 1 121.854 52.687 121.894 69.9575 ;
      RECT MASK 1 122.232 52.687 122.272 69.9575 ;
      RECT MASK 1 122.61 52.687 122.65 69.9575 ;
      RECT MASK 1 122.988 52.687 123.028 69.9575 ;
      RECT MASK 1 123.366 52.687 123.406 69.9575 ;
      RECT MASK 1 123.744 52.687 123.784 69.9575 ;
      RECT MASK 1 124.122 52.687 124.162 69.9575 ;
      RECT MASK 1 124.5 52.687 124.54 69.9575 ;
      RECT MASK 1 124.878 52.687 124.918 69.9575 ;
      RECT MASK 1 125.256 52.687 125.296 69.9575 ;
      RECT MASK 1 125.634 52.687 125.674 69.9575 ;
      RECT MASK 1 126.151 52.687 126.291 76.57 ;
      RECT MASK 1 80.969 58.5875 81.089 81.746 ;
      RECT MASK 1 94.205 58.5875 94.325 81.746 ;
      RECT MASK 1 8.171 58.8275 8.291 81.746 ;
      RECT MASK 1 14.789 58.8275 14.909 81.746 ;
      RECT MASK 1 21.407 58.8275 21.527 81.746 ;
      RECT MASK 1 28.025 58.8275 28.145 81.746 ;
      RECT MASK 1 34.643 58.8275 34.763 81.746 ;
      RECT MASK 1 41.261 58.8275 41.381 81.746 ;
      RECT MASK 1 47.879 58.8275 47.999 81.746 ;
      RECT MASK 1 54.497 58.8275 54.617 81.746 ;
      RECT MASK 1 61.115 58.8275 61.235 81.746 ;
      RECT MASK 1 67.733 58.8275 67.853 81.746 ;
      RECT MASK 1 74.351 58.8275 74.471 81.746 ;
      RECT MASK 1 87.587 58.8275 87.707 81.746 ;
      RECT MASK 1 100.823 58.8275 100.943 81.746 ;
      RECT MASK 1 107.441 58.8275 107.561 81.746 ;
      RECT MASK 1 9.333 64.6885 9.453 81.746 ;
      RECT MASK 1 22.569 64.6885 22.689 81.746 ;
      RECT MASK 1 35.805 64.6885 35.925 81.746 ;
      RECT MASK 1 49.041 64.6885 49.161 81.746 ;
      RECT MASK 1 62.277 64.6885 62.397 81.746 ;
      RECT MASK 1 75.513 64.6885 75.633 81.746 ;
      RECT MASK 1 88.749 64.6885 88.869 81.746 ;
      RECT MASK 1 101.985 64.6885 102.105 81.746 ;
      RECT MASK 1 13.627 64.8465 13.747 81.746 ;
      RECT MASK 1 26.863 64.8465 26.983 81.746 ;
      RECT MASK 1 40.099 64.8465 40.219 81.746 ;
      RECT MASK 1 53.335 64.8465 53.455 81.746 ;
      RECT MASK 1 66.571 64.8465 66.691 81.746 ;
      RECT MASK 1 79.807 64.8465 79.927 81.746 ;
      RECT MASK 1 93.043 64.8465 93.163 81.746 ;
      RECT MASK 1 106.279 64.8465 106.399 81.746 ;
      RECT MASK 1 105.117 70.8115 105.237 81.746 ;
      RECT MASK 1 117.318 70.8925 117.358 76.57 ;
      RECT MASK 1 117.696 70.8925 117.736 76.57 ;
      RECT MASK 1 118.074 70.8925 118.114 76.57 ;
      RECT MASK 1 118.452 70.8925 118.492 76.57 ;
      RECT MASK 1 118.83 70.8925 118.87 76.57 ;
      RECT MASK 1 119.208 70.8925 119.248 76.57 ;
      RECT MASK 1 119.586 70.8925 119.626 76.57 ;
      RECT MASK 1 119.964 70.8925 120.004 76.57 ;
      RECT MASK 1 120.342 70.8925 120.382 76.57 ;
      RECT MASK 1 120.72 70.8925 120.76 76.57 ;
      RECT MASK 1 121.098 70.8925 121.138 76.57 ;
      RECT MASK 1 121.476 70.8925 121.516 76.57 ;
      RECT MASK 1 121.854 70.8925 121.894 76.57 ;
      RECT MASK 1 122.232 70.8925 122.272 76.57 ;
      RECT MASK 1 122.61 70.8925 122.65 76.57 ;
      RECT MASK 1 122.988 70.8925 123.028 76.57 ;
      RECT MASK 1 123.366 70.8925 123.406 76.57 ;
      RECT MASK 1 123.744 70.8925 123.784 76.57 ;
      RECT MASK 1 124.122 70.8925 124.162 76.57 ;
      RECT MASK 1 124.5 70.8925 124.54 76.57 ;
      RECT MASK 1 124.878 70.8925 124.918 76.57 ;
      RECT MASK 1 125.256 70.8925 125.296 76.57 ;
      RECT MASK 1 125.634 70.8925 125.674 76.57 ;
      RECT MASK 1 12.465 71.0515 12.585 81.746 ;
      RECT MASK 1 25.701 71.0515 25.821 81.746 ;
      RECT MASK 1 38.937 71.0515 39.057 81.746 ;
      RECT MASK 1 52.173 71.0515 52.293 81.746 ;
      RECT MASK 1 65.409 71.0515 65.529 81.746 ;
      RECT MASK 1 78.645 71.0515 78.765 81.746 ;
      RECT MASK 1 91.881 71.0515 92.001 81.746 ;
      RECT MASK 1 116.323 77.12 116.463 80.393 ;
      RECT MASK 1 117.318 77.12 117.358 79.4 ;
      RECT MASK 1 117.696 77.12 117.736 79.4 ;
      RECT MASK 1 118.074 77.12 118.114 79.4 ;
      RECT MASK 1 118.452 77.12 118.492 79.4 ;
      RECT MASK 1 118.83 77.12 118.87 79.4 ;
      RECT MASK 1 119.208 77.12 119.248 79.4 ;
      RECT MASK 1 119.586 77.12 119.626 79.4 ;
      RECT MASK 1 119.964 77.12 120.004 79.4 ;
      RECT MASK 1 120.342 77.12 120.382 79.4 ;
      RECT MASK 1 120.72 77.12 120.76 79.4 ;
      RECT MASK 1 121.098 77.12 121.138 79.4 ;
      RECT MASK 1 121.476 77.12 121.516 79.4 ;
      RECT MASK 1 121.854 77.12 121.894 79.4 ;
      RECT MASK 1 122.232 77.12 122.272 79.4 ;
      RECT MASK 1 122.61 77.12 122.65 79.4 ;
      RECT MASK 1 122.988 77.12 123.028 79.4 ;
      RECT MASK 1 123.366 77.12 123.406 79.4 ;
      RECT MASK 1 123.744 77.12 123.784 79.4 ;
      RECT MASK 1 124.122 77.12 124.162 79.4 ;
      RECT MASK 1 124.5 77.12 124.54 79.4 ;
      RECT MASK 1 124.878 77.12 124.918 79.4 ;
      RECT MASK 1 125.256 77.12 125.296 79.4 ;
      RECT MASK 1 125.634 77.12 125.674 79.4 ;
      RECT MASK 1 126.151 77.12 126.291 80.393 ;
      RECT MASK 1 2.341 79.12 2.401 95.78 ;
      RECT MASK 1 2.615 79.12 2.675 95.78 ;
      RECT MASK 1 2.889 79.12 2.949 95.78 ;
      RECT MASK 1 3.163 79.12 3.223 95.78 ;
      RECT MASK 1 3.437 79.12 3.497 95.78 ;
      RECT MASK 1 3.711 79.12 3.771 95.78 ;
      RECT MASK 1 3.985 79.12 4.045 95.78 ;
      RECT MASK 1 4.259 79.12 4.319 95.78 ;
      RECT MASK 1 57.289 80.465 57.409 84.25 ;
      RECT MASK 1 57.667 80.465 57.787 84.25 ;
      RECT MASK 1 58.045 80.465 58.165 84.25 ;
      RECT MASK 1 63.275 80.465 63.395 84.25 ;
      RECT MASK 1 63.653 80.465 63.773 84.25 ;
      RECT MASK 1 64.031 80.465 64.151 84.25 ;
      RECT MASK 1 111.15 80.65 111.27 84.174 ;
      RECT MASK 1 111.793 80.65 111.913 84.174 ;
      RECT MASK 1 112.284 80.65 112.404 84.174 ;
      RECT MASK 1 112.892 80.65 113.012 84.174 ;
      RECT MASK 1 116.736 81.814 116.796 96.653 ;
      RECT MASK 1 117.01 81.814 117.07 96.653 ;
      RECT MASK 1 117.284 81.814 117.344 96.653 ;
      RECT MASK 1 117.558 81.814 117.618 96.653 ;
      RECT MASK 1 117.832 81.814 117.892 96.653 ;
      RECT MASK 1 118.106 81.814 118.166 96.653 ;
      RECT MASK 1 118.38 81.814 118.44 96.653 ;
      RECT MASK 1 118.654 81.814 118.714 96.653 ;
      RECT MASK 1 118.928 81.814 118.988 96.653 ;
      RECT MASK 1 119.202 81.814 119.262 96.653 ;
      RECT MASK 1 119.476 81.814 119.536 96.653 ;
      RECT MASK 1 119.75 81.814 119.81 96.653 ;
      RECT MASK 1 120.024 81.814 120.084 96.653 ;
      RECT MASK 1 120.298 81.814 120.358 96.653 ;
      RECT MASK 1 120.572 81.814 120.632 96.653 ;
      RECT MASK 1 120.846 81.814 120.906 96.653 ;
      RECT MASK 1 121.12 81.814 121.18 96.653 ;
      RECT MASK 1 121.394 81.814 121.454 96.653 ;
      RECT MASK 1 121.668 81.814 121.728 96.653 ;
      RECT MASK 1 121.942 81.814 122.002 96.653 ;
      RECT MASK 1 122.216 81.814 122.276 96.653 ;
      RECT MASK 1 122.49 81.814 122.55 96.653 ;
      RECT MASK 1 122.764 81.814 122.824 96.653 ;
      RECT MASK 1 123.038 81.814 123.098 96.653 ;
      RECT MASK 1 123.312 81.814 123.372 96.653 ;
      RECT MASK 1 123.586 81.814 123.646 96.653 ;
      RECT MASK 1 123.86 81.814 123.92 96.653 ;
      RECT MASK 1 124.134 81.814 124.194 96.653 ;
      RECT MASK 1 124.408 81.814 124.468 96.653 ;
      RECT MASK 1 124.682 81.814 124.742 96.653 ;
      RECT MASK 1 124.956 81.814 125.016 96.653 ;
      RECT MASK 1 125.23 81.814 125.29 96.653 ;
      RECT MASK 1 125.504 81.814 125.564 96.653 ;
      RECT MASK 1 125.778 81.814 125.838 96.653 ;
      RECT MASK 1 126.052 81.814 126.112 96.653 ;
      RECT MASK 1 126.326 81.814 126.386 96.653 ;
      RECT MASK 1 126.6 81.814 126.66 96.653 ;
      RECT MASK 1 126.874 81.814 126.934 96.653 ;
      RECT MASK 1 127.148 81.814 127.208 96.653 ;
      RECT MASK 1 127.422 81.814 127.482 96.653 ;
      RECT MASK 1 58.798 81.95 58.878 84.25 ;
      RECT MASK 1 59.973 81.95 60.053 84.25 ;
      RECT MASK 1 61.135 81.95 61.215 84.25 ;
      RECT MASK 1 62.297 81.95 62.377 84.25 ;
      RECT MASK 1 59.188 82.1185 59.268 84.25 ;
      RECT MASK 1 60.351 82.1185 60.431 84.25 ;
      RECT MASK 1 61.513 82.1185 61.593 84.25 ;
      RECT MASK 1 62.675 82.1185 62.755 84.25 ;
      RECT MASK 1 59.585 83.944 59.685 84.25 ;
      RECT MASK 1 60.747 83.944 60.847 84.25 ;
      RECT MASK 1 61.909 83.944 62.009 84.25 ;
      RECT MASK 1 69.727 86.285 71.692 86.485 ;
      RECT MASK 1 103.89 86.285 106.869 86.485 ;
      RECT MASK 1 35.562 86.35 35.922 95.33 ;
      RECT MASK 1 66.88 86.35 67.24 95.33 ;
      RECT MASK 1 71.952 86.35 72.312 95.33 ;
      RECT MASK 1 103.27 86.35 103.63 95.33 ;
      RECT MASK 1 32.279 86.375 35.302 86.575 ;
      RECT MASK 1 67.5685 86.375 69.467 86.575 ;
      RECT MASK 1 26.225 86.43 26.285 92.31 ;
      RECT MASK 1 26.495 86.43 26.555 92.31 ;
      RECT MASK 1 26.765 86.43 26.825 92.31 ;
      RECT MASK 1 27.035 86.43 27.095 92.31 ;
      RECT MASK 1 27.305 86.43 27.365 92.31 ;
      RECT MASK 1 27.575 86.43 27.635 92.31 ;
      RECT MASK 1 27.845 86.43 27.905 92.31 ;
      RECT MASK 1 28.115 86.43 28.175 92.31 ;
      RECT MASK 1 28.385 86.43 28.445 92.31 ;
      RECT MASK 1 28.655 86.43 28.715 92.31 ;
      RECT MASK 1 28.925 86.43 28.985 92.31 ;
      RECT MASK 1 29.195 86.43 29.255 92.31 ;
      RECT MASK 1 29.465 86.43 29.525 92.31 ;
      RECT MASK 1 29.735 86.43 29.795 92.31 ;
      RECT MASK 1 30.005 86.43 30.065 92.31 ;
      RECT MASK 1 36.2245 86.469 66.5775 86.569 ;
      RECT MASK 1 72.6145 86.469 102.9675 86.569 ;
      RECT MASK 1 69.727 86.735 71.692 86.935 ;
      RECT MASK 1 103.89 86.735 106.869 86.935 ;
      RECT MASK 1 32.279 86.825 35.302 87.025 ;
      RECT MASK 1 67.5715 86.825 69.467 87.025 ;
      RECT MASK 1 14.9155 87.06 14.9955 89.2865 ;
      RECT MASK 1 15.2475 87.06 15.3275 89.2865 ;
      RECT MASK 1 25.864 87.101 25.924 88.982 ;
      RECT MASK 1 30.366 87.101 30.426 88.982 ;
      RECT MASK 1 37.048 87.147 65.754 87.207 ;
      RECT MASK 1 73.438 87.147 102.144 87.207 ;
      RECT MASK 1 17.061 87.19 17.161 94.37 ;
      RECT MASK 1 67.5 87.24 71.692 87.34 ;
      RECT MASK 1 103.89 87.24 106.869 87.34 ;
      RECT MASK 1 8.195 87.244 8.295 94.316 ;
      RECT MASK 1 12.677 87.244 12.777 94.316 ;
      RECT MASK 1 13.243 87.244 13.343 94.316 ;
      RECT MASK 1 17.627 87.244 17.727 94.316 ;
      RECT MASK 1 22.109 87.244 22.209 94.316 ;
      RECT MASK 1 32.279 87.255 35.302 87.355 ;
      RECT MASK 1 37.048 87.399 65.754 87.459 ;
      RECT MASK 1 73.438 87.399 102.144 87.459 ;
      RECT MASK 1 9.7015 87.52 9.7815 89.2865 ;
      RECT MASK 1 10.0335 87.52 10.1135 89.2865 ;
      RECT MASK 1 10.3655 87.52 10.4455 89.2865 ;
      RECT MASK 1 10.6975 87.52 10.7775 89.2865 ;
      RECT MASK 1 11.0295 87.52 11.1095 89.2865 ;
      RECT MASK 1 19.1335 87.52 19.2135 89.2865 ;
      RECT MASK 1 19.4655 87.52 19.5455 89.2865 ;
      RECT MASK 1 19.7975 87.52 19.8775 89.2865 ;
      RECT MASK 1 20.1295 87.52 20.2095 89.2865 ;
      RECT MASK 1 20.4615 87.52 20.5415 89.2865 ;
      RECT MASK 1 67.5 87.592 71.692 87.692 ;
      RECT MASK 1 103.89 87.592 106.869 87.692 ;
      RECT MASK 1 32.279 87.607 35.302 87.707 ;
      RECT MASK 1 13.8265 87.66 13.9265 90.24 ;
      RECT MASK 1 16.4825 87.66 16.5825 90.24 ;
      RECT MASK 1 107.694 87.72 107.754 96.653 ;
      RECT MASK 1 107.968 87.72 108.028 96.653 ;
      RECT MASK 1 108.242 87.72 108.302 96.653 ;
      RECT MASK 1 108.516 87.72 108.576 96.653 ;
      RECT MASK 1 108.79 87.72 108.85 96.653 ;
      RECT MASK 1 109.064 87.72 109.124 96.653 ;
      RECT MASK 1 109.338 87.72 109.398 96.653 ;
      RECT MASK 1 109.612 87.72 109.672 96.653 ;
      RECT MASK 1 109.886 87.72 109.946 96.653 ;
      RECT MASK 1 110.16 87.72 110.22 96.653 ;
      RECT MASK 1 110.434 87.72 110.494 96.653 ;
      RECT MASK 1 110.708 87.72 110.768 96.653 ;
      RECT MASK 1 110.982 87.72 111.042 96.653 ;
      RECT MASK 1 111.256 87.72 111.316 96.653 ;
      RECT MASK 1 111.53 87.72 111.59 96.653 ;
      RECT MASK 1 111.804 87.72 111.864 96.653 ;
      RECT MASK 1 112.078 87.72 112.138 96.653 ;
      RECT MASK 1 112.352 87.72 112.412 96.653 ;
      RECT MASK 1 112.626 87.72 112.686 96.653 ;
      RECT MASK 1 112.9 87.72 112.96 96.653 ;
      RECT MASK 1 113.174 87.72 113.234 96.653 ;
      RECT MASK 1 113.448 87.72 113.508 96.653 ;
      RECT MASK 1 113.722 87.72 113.782 96.653 ;
      RECT MASK 1 113.996 87.72 114.056 96.653 ;
      RECT MASK 1 114.27 87.72 114.33 96.653 ;
      RECT MASK 1 114.544 87.72 114.604 96.653 ;
      RECT MASK 1 114.818 87.72 114.878 96.653 ;
      RECT MASK 1 115.092 87.72 115.152 96.653 ;
      RECT MASK 1 115.366 87.72 115.426 96.653 ;
      RECT MASK 1 115.64 87.72 115.7 96.653 ;
      RECT MASK 1 115.914 87.72 115.974 96.653 ;
      RECT MASK 1 116.188 87.72 116.248 96.653 ;
      RECT MASK 1 116.462 87.72 116.522 96.653 ;
      RECT MASK 1 67.5 87.944 71.692 88.044 ;
      RECT MASK 1 103.89 87.944 106.869 88.044 ;
      RECT MASK 1 32.279 87.959 35.302 88.059 ;
      RECT MASK 1 37.048 88.047 65.754 88.107 ;
      RECT MASK 1 73.438 88.047 102.144 88.107 ;
      RECT MASK 1 8.6115 88.08 8.7315 89.7135 ;
      RECT MASK 1 9.0115 88.08 9.1315 88.7365 ;
      RECT MASK 1 11.8115 88.08 11.9315 88.7365 ;
      RECT MASK 1 12.266 88.08 12.386 89.7135 ;
      RECT MASK 1 14.2115 88.08 14.3315 88.7365 ;
      RECT MASK 1 16.0115 88.08 16.1315 88.7365 ;
      RECT MASK 1 16.7565 88.08 16.8765 89.7135 ;
      RECT MASK 1 67.5 88.296 71.692 88.396 ;
      RECT MASK 1 103.89 88.296 106.869 88.396 ;
      RECT MASK 1 37.048 88.299 65.754 88.359 ;
      RECT MASK 1 73.438 88.299 102.144 88.359 ;
      RECT MASK 1 32.279 88.311 35.302 88.411 ;
      RECT MASK 1 11.3615 88.412 11.4415 89.8155 ;
      RECT MASK 1 20.7935 88.412 20.8735 89.8155 ;
      RECT MASK 1 67.5 88.648 71.692 88.748 ;
      RECT MASK 1 103.89 88.648 106.869 88.748 ;
      RECT MASK 1 32.279 88.663 35.302 88.763 ;
      RECT MASK 1 37.048 88.947 65.754 89.007 ;
      RECT MASK 1 73.438 88.947 102.144 89.007 ;
      RECT MASK 1 67.5 89 71.692 89.1 ;
      RECT MASK 1 103.89 89 106.869 89.1 ;
      RECT MASK 1 32.279 89.015 35.302 89.115 ;
      RECT MASK 1 9.0375 89.025 9.1175 92.535 ;
      RECT MASK 1 9.3695 89.025 9.4495 92.535 ;
      RECT MASK 1 11.6935 89.025 11.7735 92.535 ;
      RECT MASK 1 14.2515 89.025 14.3315 90.39 ;
      RECT MASK 1 15.9115 89.025 15.9915 90.39 ;
      RECT MASK 1 16.2435 89.025 16.3235 90.39 ;
      RECT MASK 1 18.4695 89.025 18.5495 92.535 ;
      RECT MASK 1 18.8015 89.025 18.8815 92.535 ;
      RECT MASK 1 21.1255 89.025 21.2055 92.535 ;
      RECT MASK 1 37.048 89.199 65.754 89.259 ;
      RECT MASK 1 73.438 89.199 102.144 89.259 ;
      RECT MASK 1 67.5 89.352 71.692 89.452 ;
      RECT MASK 1 103.89 89.352 106.869 89.452 ;
      RECT MASK 1 32.279 89.367 35.302 89.467 ;
      RECT MASK 1 25.864 89.441 25.924 91.322 ;
      RECT MASK 1 30.366 89.441 30.426 91.322 ;
      RECT MASK 1 67.5 89.704 71.692 89.804 ;
      RECT MASK 1 103.89 89.704 106.869 89.804 ;
      RECT MASK 1 32.279 89.719 35.302 89.819 ;
      RECT MASK 1 9.8655 89.8275 9.9455 91.7075 ;
      RECT MASK 1 10.1995 89.8275 10.2795 91.7075 ;
      RECT MASK 1 10.5325 89.8275 10.6125 91.7075 ;
      RECT MASK 1 10.8655 89.8275 10.9455 91.7075 ;
      RECT MASK 1 14.581 89.8275 14.661 91.913 ;
      RECT MASK 1 14.911 89.8275 14.991 91.913 ;
      RECT MASK 1 15.244 89.8275 15.324 91.913 ;
      RECT MASK 1 15.577 89.8275 15.657 91.913 ;
      RECT MASK 1 19.2995 89.8275 19.3795 91.665 ;
      RECT MASK 1 19.6335 89.8275 19.7135 91.665 ;
      RECT MASK 1 19.9665 89.8275 20.0465 91.665 ;
      RECT MASK 1 20.2995 89.8275 20.3795 91.665 ;
      RECT MASK 1 37.048 89.847 65.754 89.907 ;
      RECT MASK 1 73.438 89.847 102.144 89.907 ;
      RECT MASK 1 13.4905 90.0145 13.5705 94.3995 ;
      RECT MASK 1 16.8375 90.03 16.9175 94.3995 ;
      RECT MASK 1 67.5 90.056 71.692 90.156 ;
      RECT MASK 1 103.89 90.056 106.869 90.156 ;
      RECT MASK 1 32.279 90.071 35.302 90.171 ;
      RECT MASK 1 37.048 90.099 65.754 90.159 ;
      RECT MASK 1 73.438 90.099 102.144 90.159 ;
      RECT MASK 1 67.5 90.408 71.692 90.508 ;
      RECT MASK 1 103.89 90.408 106.869 90.508 ;
      RECT MASK 1 32.279 90.423 35.302 90.523 ;
      RECT MASK 1 37.048 90.747 65.754 90.807 ;
      RECT MASK 1 73.438 90.747 102.144 90.807 ;
      RECT MASK 1 67.5 90.76 71.692 90.86 ;
      RECT MASK 1 103.89 90.76 106.869 90.86 ;
      RECT MASK 1 32.279 90.775 35.302 90.875 ;
      RECT MASK 1 37.048 90.999 65.754 91.059 ;
      RECT MASK 1 73.438 90.999 102.144 91.059 ;
      RECT MASK 1 67.5 91.112 71.692 91.212 ;
      RECT MASK 1 103.89 91.112 106.869 91.212 ;
      RECT MASK 1 32.279 91.127 35.302 91.227 ;
      RECT MASK 1 14.2515 91.17 14.3315 92.535 ;
      RECT MASK 1 15.9115 91.17 15.9915 92.535 ;
      RECT MASK 1 16.2435 91.17 16.3235 92.535 ;
      RECT MASK 1 13.8265 91.32 13.9265 94.3995 ;
      RECT MASK 1 16.4825 91.32 16.5825 94.3995 ;
      RECT MASK 1 67.5 91.464 71.692 91.564 ;
      RECT MASK 1 103.89 91.464 106.869 91.564 ;
      RECT MASK 1 32.279 91.479 35.302 91.579 ;
      RECT MASK 1 37.048 91.647 65.754 91.707 ;
      RECT MASK 1 73.438 91.647 102.144 91.707 ;
      RECT MASK 1 11.3615 91.7445 11.4415 93.148 ;
      RECT MASK 1 20.7935 91.7445 20.8735 93.148 ;
      RECT MASK 1 67.5 91.816 71.692 91.916 ;
      RECT MASK 1 103.89 91.816 106.869 91.916 ;
      RECT MASK 1 32.279 91.831 35.302 91.931 ;
      RECT MASK 1 37.048 91.899 65.754 91.959 ;
      RECT MASK 1 73.438 91.899 102.144 91.959 ;
      RECT MASK 1 25.415 91.919 25.475 92.31 ;
      RECT MASK 1 25.685 91.919 25.745 92.31 ;
      RECT MASK 1 25.955 91.919 26.015 92.31 ;
      RECT MASK 1 30.275 91.919 30.335 92.31 ;
      RECT MASK 1 30.545 91.919 30.605 92.31 ;
      RECT MASK 1 30.815 91.919 30.875 92.31 ;
      RECT MASK 1 67.5 92.168 71.692 92.268 ;
      RECT MASK 1 103.89 92.168 106.869 92.268 ;
      RECT MASK 1 32.279 92.183 35.302 92.283 ;
      RECT MASK 1 9.7015 92.2735 9.7815 94.04 ;
      RECT MASK 1 10.0335 92.2735 10.1135 94.04 ;
      RECT MASK 1 10.3655 92.2735 10.4455 94.04 ;
      RECT MASK 1 10.6975 92.2735 10.7775 94.04 ;
      RECT MASK 1 14.9155 92.2735 14.9955 94.5 ;
      RECT MASK 1 15.2475 92.2735 15.3275 94.5 ;
      RECT MASK 1 19.1335 92.2735 19.2135 94.04 ;
      RECT MASK 1 19.4655 92.2735 19.5455 94.04 ;
      RECT MASK 1 19.7975 92.2735 19.8775 94.04 ;
      RECT MASK 1 20.1295 92.2735 20.2095 94.04 ;
      RECT MASK 1 20.4615 92.2735 20.5415 94.04 ;
      RECT MASK 1 67.5 92.52 71.692 92.62 ;
      RECT MASK 1 103.89 92.52 106.869 92.62 ;
      RECT MASK 1 32.279 92.535 35.302 92.635 ;
      RECT MASK 1 37.048 92.547 65.754 92.607 ;
      RECT MASK 1 73.438 92.547 102.144 92.607 ;
      RECT MASK 1 14.2515 92.7795 14.3315 94.3995 ;
      RECT MASK 1 14.5835 92.7795 14.6635 94.3995 ;
      RECT MASK 1 15.5795 92.7795 15.6595 94.3995 ;
      RECT MASK 1 15.9115 92.7795 15.9915 94.3995 ;
      RECT MASK 1 16.2445 92.7795 16.3245 94.3995 ;
      RECT MASK 1 37.048 92.799 65.754 92.859 ;
      RECT MASK 1 73.438 92.799 102.144 92.859 ;
      RECT MASK 1 67.5 92.872 71.692 92.972 ;
      RECT MASK 1 103.89 92.872 106.869 92.972 ;
      RECT MASK 1 32.279 92.887 35.302 92.987 ;
      RECT MASK 1 67.5 93.224 71.692 93.324 ;
      RECT MASK 1 103.89 93.224 106.869 93.324 ;
      RECT MASK 1 32.279 93.239 35.302 93.339 ;
      RECT MASK 1 37.048 93.447 65.754 93.507 ;
      RECT MASK 1 73.438 93.447 102.144 93.507 ;
      RECT MASK 1 67.5 93.576 71.692 93.676 ;
      RECT MASK 1 103.89 93.576 106.869 93.676 ;
      RECT MASK 1 32.279 93.591 35.302 93.691 ;
      RECT MASK 1 37.048 93.699 65.754 93.759 ;
      RECT MASK 1 73.438 93.699 102.144 93.759 ;
      RECT MASK 1 67.5 93.928 71.692 94.028 ;
      RECT MASK 1 103.89 93.928 106.869 94.028 ;
      RECT MASK 1 32.279 93.943 35.302 94.043 ;
      RECT MASK 1 67.5 94.28 71.692 94.38 ;
      RECT MASK 1 103.89 94.28 106.869 94.38 ;
      RECT MASK 1 32.279 94.295 35.302 94.395 ;
      RECT MASK 1 37.048 94.347 65.754 94.407 ;
      RECT MASK 1 73.438 94.347 102.144 94.407 ;
      RECT MASK 1 37.048 94.599 65.754 94.659 ;
      RECT MASK 1 73.438 94.599 102.144 94.659 ;
      RECT MASK 1 32.279 94.655 35.302 94.855 ;
      RECT MASK 1 67.5 94.655 69.471 94.855 ;
      RECT MASK 1 69.731 94.745 71.692 94.945 ;
      RECT MASK 1 103.89 94.745 106.869 94.945 ;
      RECT MASK 1 32.279 95.105 35.302 95.305 ;
      RECT MASK 1 67.5 95.105 69.471 95.305 ;
      RECT MASK 1 36.2245 95.111 66.5775 95.211 ;
      RECT MASK 1 72.6145 95.111 102.9675 95.211 ;
      RECT MASK 1 69.731 95.195 71.692 95.395 ;
      RECT MASK 1 103.89 95.195 106.869 95.395 ;
      RECT MASK 1 2.475 97.41 2.535 108.838 ;
      RECT MASK 1 2.749 97.41 2.809 108.838 ;
      RECT MASK 1 3.023 97.41 3.083 108.838 ;
      RECT MASK 1 3.297 97.41 3.357 108.838 ;
      RECT MASK 1 3.571 97.41 3.631 108.838 ;
      RECT MASK 1 3.845 97.41 3.905 108.838 ;
      RECT MASK 1 4.119 97.41 4.179 108.838 ;
      RECT MASK 1 4.393 97.41 4.453 108.838 ;
      RECT MASK 1 4.667 97.41 4.727 108.838 ;
      RECT MASK 1 4.941 97.41 5.001 108.838 ;
      RECT MASK 1 5.215 97.41 5.275 108.838 ;
      RECT MASK 1 5.489 97.41 5.549 108.838 ;
      RECT MASK 1 5.763 97.41 5.823 108.838 ;
      RECT MASK 1 6.037 97.41 6.097 108.838 ;
      RECT MASK 1 6.311 97.41 6.371 108.838 ;
      RECT MASK 1 6.585 97.41 6.645 108.838 ;
      RECT MASK 1 6.859 97.41 6.919 108.838 ;
      RECT MASK 1 7.133 97.41 7.193 108.838 ;
      RECT MASK 1 7.407 97.41 7.467 108.838 ;
      RECT MASK 1 7.681 97.41 7.741 108.838 ;
      RECT MASK 1 7.955 97.41 8.015 108.838 ;
      RECT MASK 1 8.229 97.41 8.289 108.838 ;
      RECT MASK 1 8.503 97.41 8.563 108.838 ;
      RECT MASK 1 8.777 97.41 8.837 108.838 ;
      RECT MASK 1 9.051 97.41 9.111 108.838 ;
      RECT MASK 1 9.325 97.41 9.385 108.838 ;
      RECT MASK 1 9.599 97.41 9.659 108.838 ;
      RECT MASK 1 9.873 97.41 9.933 108.838 ;
      RECT MASK 1 10.147 97.41 10.207 108.838 ;
      RECT MASK 1 10.421 97.41 10.481 108.838 ;
      RECT MASK 1 10.695 97.41 10.755 108.838 ;
      RECT MASK 1 10.969 97.41 11.029 108.838 ;
      RECT MASK 1 11.243 97.41 11.303 108.838 ;
      RECT MASK 1 11.517 97.41 11.577 108.838 ;
      RECT MASK 1 11.791 97.41 11.851 108.838 ;
      RECT MASK 1 12.065 97.41 12.125 108.838 ;
      RECT MASK 1 12.339 97.41 12.399 108.838 ;
      RECT MASK 1 12.613 97.41 12.673 108.838 ;
      RECT MASK 1 12.887 97.41 12.947 108.838 ;
      RECT MASK 1 13.161 97.41 13.221 108.838 ;
      RECT MASK 1 13.435 97.41 13.495 108.838 ;
      RECT MASK 1 13.709 97.41 13.769 108.838 ;
      RECT MASK 1 13.983 97.41 14.043 108.838 ;
      RECT MASK 1 14.257 97.41 14.317 108.838 ;
      RECT MASK 1 14.531 97.41 14.591 108.838 ;
      RECT MASK 1 14.805 97.41 14.865 108.838 ;
      RECT MASK 1 15.079 97.41 15.139 108.838 ;
      RECT MASK 1 15.353 97.41 15.413 108.838 ;
      RECT MASK 1 15.627 97.41 15.687 108.838 ;
      RECT MASK 1 15.901 97.41 15.961 108.838 ;
      RECT MASK 1 16.175 97.41 16.235 108.838 ;
      RECT MASK 1 16.449 97.41 16.509 108.838 ;
      RECT MASK 1 16.723 97.41 16.783 108.838 ;
      RECT MASK 1 16.997 97.41 17.057 108.838 ;
      RECT MASK 1 17.271 97.41 17.331 108.838 ;
      RECT MASK 1 17.545 97.41 17.605 108.838 ;
      RECT MASK 1 17.819 97.41 17.879 108.838 ;
      RECT MASK 1 18.093 97.41 18.153 108.838 ;
      RECT MASK 1 18.367 97.41 18.427 108.838 ;
      RECT MASK 1 18.641 97.41 18.701 108.838 ;
      RECT MASK 1 18.915 97.41 18.975 108.838 ;
      RECT MASK 1 19.189 97.41 19.249 108.838 ;
      RECT MASK 1 19.463 97.41 19.523 108.838 ;
      RECT MASK 1 19.737 97.41 19.797 108.838 ;
      RECT MASK 1 20.011 97.41 20.071 108.838 ;
      RECT MASK 1 20.285 97.41 20.345 108.838 ;
      RECT MASK 1 20.559 97.41 20.619 108.838 ;
      RECT MASK 1 20.833 97.41 20.893 108.838 ;
      RECT MASK 1 21.107 97.41 21.167 108.838 ;
      RECT MASK 1 21.381 97.41 21.441 108.838 ;
      RECT MASK 1 21.655 97.41 21.715 108.838 ;
      RECT MASK 1 21.929 97.41 21.989 108.838 ;
      RECT MASK 1 22.203 97.41 22.263 108.838 ;
      RECT MASK 1 22.477 97.41 22.537 108.838 ;
      RECT MASK 1 22.751 97.41 22.811 108.838 ;
      RECT MASK 1 23.025 97.41 23.085 108.838 ;
      RECT MASK 1 23.299 97.41 23.359 108.838 ;
      RECT MASK 1 23.573 97.41 23.633 108.838 ;
      RECT MASK 1 23.847 97.41 23.907 108.838 ;
      RECT MASK 1 24.121 97.41 24.181 108.838 ;
      RECT MASK 1 24.395 97.41 24.455 108.838 ;
      RECT MASK 1 24.669 97.41 24.729 108.838 ;
      RECT MASK 1 24.943 97.41 25.003 108.838 ;
      RECT MASK 1 25.217 97.41 25.277 108.838 ;
      RECT MASK 1 25.491 97.41 25.551 108.838 ;
      RECT MASK 1 25.765 97.41 25.825 108.838 ;
      RECT MASK 1 26.039 97.41 26.099 108.838 ;
      RECT MASK 1 26.313 97.41 26.373 108.838 ;
      RECT MASK 1 26.587 97.41 26.647 108.838 ;
      RECT MASK 1 26.861 97.41 26.921 108.838 ;
      RECT MASK 1 27.135 97.41 27.195 108.838 ;
      RECT MASK 1 27.409 97.41 27.469 108.838 ;
      RECT MASK 1 27.683 97.41 27.743 108.838 ;
      RECT MASK 1 27.957 97.41 28.017 108.838 ;
      RECT MASK 1 28.231 97.41 28.291 108.838 ;
      RECT MASK 1 28.505 97.41 28.565 108.838 ;
      RECT MASK 1 28.779 97.41 28.839 108.838 ;
      RECT MASK 1 29.053 97.41 29.113 108.838 ;
      RECT MASK 1 29.327 97.41 29.387 108.838 ;
      RECT MASK 1 29.601 97.41 29.661 108.838 ;
      RECT MASK 1 29.875 97.41 29.935 108.838 ;
      RECT MASK 1 30.149 97.41 30.209 108.838 ;
      RECT MASK 1 30.423 97.41 30.483 108.838 ;
      RECT MASK 1 30.697 97.41 30.757 108.838 ;
      RECT MASK 1 30.971 97.41 31.031 108.838 ;
      RECT MASK 1 31.245 97.41 31.305 108.838 ;
      RECT MASK 1 31.519 97.41 31.579 108.838 ;
      RECT MASK 1 31.793 97.41 31.853 108.838 ;
      RECT MASK 1 32.067 97.41 32.127 108.838 ;
      RECT MASK 1 32.341 97.41 32.401 108.838 ;
      RECT MASK 1 32.615 97.41 32.675 108.838 ;
      RECT MASK 1 32.889 97.41 32.949 108.838 ;
      RECT MASK 1 33.163 97.41 33.223 108.838 ;
      RECT MASK 1 33.437 97.41 33.497 108.838 ;
      RECT MASK 1 33.711 97.41 33.771 108.838 ;
      RECT MASK 1 33.985 97.41 34.045 108.838 ;
      RECT MASK 1 34.259 97.41 34.319 108.838 ;
      RECT MASK 1 34.533 97.41 34.593 108.838 ;
      RECT MASK 1 34.807 97.41 34.867 108.838 ;
      RECT MASK 1 35.081 97.41 35.141 108.838 ;
      RECT MASK 1 35.355 97.41 35.415 108.838 ;
      RECT MASK 1 35.629 97.41 35.689 108.838 ;
      RECT MASK 1 35.903 97.41 35.963 108.838 ;
      RECT MASK 1 36.177 97.41 36.237 108.838 ;
      RECT MASK 1 36.451 97.41 36.511 108.838 ;
      RECT MASK 1 36.725 97.41 36.785 108.838 ;
      RECT MASK 1 36.999 97.41 37.059 108.838 ;
      RECT MASK 1 37.273 97.41 37.333 108.838 ;
      RECT MASK 1 37.547 97.41 37.607 108.838 ;
      RECT MASK 1 37.821 97.41 37.881 108.838 ;
      RECT MASK 1 38.095 97.41 38.155 108.838 ;
      RECT MASK 1 38.369 97.41 38.429 108.838 ;
      RECT MASK 1 38.643 97.41 38.703 108.838 ;
      RECT MASK 1 38.917 97.41 38.977 108.838 ;
      RECT MASK 1 39.191 97.41 39.251 108.838 ;
      RECT MASK 1 39.465 97.41 39.525 108.838 ;
      RECT MASK 1 39.739 97.41 39.799 108.838 ;
      RECT MASK 1 40.013 97.41 40.073 108.838 ;
      RECT MASK 1 40.287 97.41 40.347 108.838 ;
      RECT MASK 1 40.561 97.41 40.621 108.838 ;
      RECT MASK 1 40.835 97.41 40.895 108.838 ;
      RECT MASK 1 41.109 97.41 41.169 108.838 ;
      RECT MASK 1 41.383 97.41 41.443 108.838 ;
      RECT MASK 1 41.657 97.41 41.717 108.838 ;
      RECT MASK 1 41.931 97.41 41.991 108.838 ;
      RECT MASK 1 42.205 97.41 42.265 108.838 ;
      RECT MASK 1 42.479 97.41 42.539 108.838 ;
      RECT MASK 1 42.753 97.41 42.813 108.838 ;
      RECT MASK 1 43.027 97.41 43.087 108.838 ;
      RECT MASK 1 43.301 97.41 43.361 108.838 ;
      RECT MASK 1 45.867 97.41 45.927 108.838 ;
      RECT MASK 1 46.141 97.41 46.201 108.838 ;
      RECT MASK 1 46.415 97.41 46.475 108.838 ;
      RECT MASK 1 46.689 97.41 46.749 108.838 ;
      RECT MASK 1 46.963 97.41 47.023 108.838 ;
      RECT MASK 1 47.237 97.41 47.297 108.838 ;
      RECT MASK 1 47.511 97.41 47.571 108.838 ;
      RECT MASK 1 47.785 97.41 47.845 108.838 ;
      RECT MASK 1 48.059 97.41 48.119 108.838 ;
      RECT MASK 1 48.333 97.41 48.393 108.838 ;
      RECT MASK 1 48.607 97.41 48.667 108.838 ;
      RECT MASK 1 48.881 97.41 48.941 108.838 ;
      RECT MASK 1 49.155 97.41 49.215 108.838 ;
      RECT MASK 1 49.429 97.41 49.489 108.838 ;
      RECT MASK 1 49.703 97.41 49.763 108.838 ;
      RECT MASK 1 49.977 97.41 50.037 108.838 ;
      RECT MASK 1 50.251 97.41 50.311 108.838 ;
      RECT MASK 1 50.525 97.41 50.585 108.838 ;
      RECT MASK 1 50.799 97.41 50.859 108.838 ;
      RECT MASK 1 51.073 97.41 51.133 108.838 ;
      RECT MASK 1 51.347 97.41 51.407 108.838 ;
      RECT MASK 1 51.621 97.41 51.681 108.838 ;
      RECT MASK 1 51.895 97.41 51.955 108.838 ;
      RECT MASK 1 52.169 97.41 52.229 108.838 ;
      RECT MASK 1 52.443 97.41 52.503 108.838 ;
      RECT MASK 1 52.717 97.41 52.777 108.838 ;
      RECT MASK 1 52.991 97.41 53.051 108.838 ;
      RECT MASK 1 53.265 97.41 53.325 108.838 ;
      RECT MASK 1 53.539 97.41 53.599 108.838 ;
      RECT MASK 1 53.813 97.41 53.873 108.838 ;
      RECT MASK 1 54.087 97.41 54.147 108.838 ;
      RECT MASK 1 54.361 97.41 54.421 108.838 ;
      RECT MASK 1 54.635 97.41 54.695 108.838 ;
      RECT MASK 1 54.909 97.41 54.969 108.838 ;
      RECT MASK 1 55.183 97.41 55.243 108.838 ;
      RECT MASK 1 55.457 97.41 55.517 108.838 ;
      RECT MASK 1 55.731 97.41 55.791 108.838 ;
      RECT MASK 1 56.005 97.41 56.065 108.838 ;
      RECT MASK 1 56.279 97.41 56.339 108.838 ;
      RECT MASK 1 56.553 97.41 56.613 108.838 ;
      RECT MASK 1 56.827 97.41 56.887 108.838 ;
      RECT MASK 1 57.101 97.41 57.161 108.838 ;
      RECT MASK 1 57.375 97.41 57.435 108.838 ;
      RECT MASK 1 57.649 97.41 57.709 108.838 ;
      RECT MASK 1 57.923 97.41 57.983 108.838 ;
      RECT MASK 1 58.197 97.41 58.257 108.838 ;
      RECT MASK 1 58.471 97.41 58.531 108.838 ;
      RECT MASK 1 58.745 97.41 58.805 108.838 ;
      RECT MASK 1 59.019 97.41 59.079 108.838 ;
      RECT MASK 1 59.293 97.41 59.353 108.838 ;
      RECT MASK 1 59.567 97.41 59.627 108.838 ;
      RECT MASK 1 59.841 97.41 59.901 108.838 ;
      RECT MASK 1 60.115 97.41 60.175 108.838 ;
      RECT MASK 1 60.389 97.41 60.449 108.838 ;
      RECT MASK 1 60.663 97.41 60.723 108.838 ;
      RECT MASK 1 60.937 97.41 60.997 108.838 ;
      RECT MASK 1 61.211 97.41 61.271 108.838 ;
      RECT MASK 1 61.485 97.41 61.545 108.838 ;
      RECT MASK 1 61.759 97.41 61.819 108.838 ;
      RECT MASK 1 62.033 97.41 62.093 108.838 ;
      RECT MASK 1 62.307 97.41 62.367 108.838 ;
      RECT MASK 1 62.581 97.41 62.641 108.838 ;
      RECT MASK 1 62.855 97.41 62.915 108.838 ;
      RECT MASK 1 63.129 97.41 63.189 108.838 ;
      RECT MASK 1 63.403 97.41 63.463 108.838 ;
      RECT MASK 1 63.677 97.41 63.737 108.838 ;
      RECT MASK 1 63.951 97.41 64.011 108.838 ;
      RECT MASK 1 64.225 97.41 64.285 108.838 ;
      RECT MASK 1 64.499 97.41 64.559 108.838 ;
      RECT MASK 1 64.773 97.41 64.833 108.838 ;
      RECT MASK 1 65.047 97.41 65.107 108.838 ;
      RECT MASK 1 65.321 97.41 65.381 108.838 ;
      RECT MASK 1 65.595 97.41 65.655 108.838 ;
      RECT MASK 1 65.869 97.41 65.929 108.838 ;
      RECT MASK 1 66.143 97.41 66.203 108.838 ;
      RECT MASK 1 66.417 97.41 66.477 108.838 ;
      RECT MASK 1 66.691 97.41 66.751 108.838 ;
      RECT MASK 1 66.965 97.41 67.025 108.838 ;
      RECT MASK 1 67.239 97.41 67.299 108.838 ;
      RECT MASK 1 67.513 97.41 67.573 108.838 ;
      RECT MASK 1 67.787 97.41 67.847 108.838 ;
      RECT MASK 1 68.061 97.41 68.121 108.838 ;
      RECT MASK 1 68.335 97.41 68.395 108.838 ;
      RECT MASK 1 68.609 97.41 68.669 108.838 ;
      RECT MASK 1 68.883 97.41 68.943 108.838 ;
      RECT MASK 1 69.157 97.41 69.217 108.838 ;
      RECT MASK 1 69.431 97.41 69.491 108.838 ;
      RECT MASK 1 69.705 97.41 69.765 108.838 ;
      RECT MASK 1 69.979 97.41 70.039 108.838 ;
      RECT MASK 1 70.253 97.41 70.313 108.838 ;
      RECT MASK 1 70.527 97.41 70.587 108.838 ;
      RECT MASK 1 70.801 97.41 70.861 108.838 ;
      RECT MASK 1 71.075 97.41 71.135 108.838 ;
      RECT MASK 1 71.349 97.41 71.409 108.838 ;
      RECT MASK 1 71.623 97.41 71.683 108.838 ;
      RECT MASK 1 71.897 97.41 71.957 108.838 ;
      RECT MASK 1 72.171 97.41 72.231 108.838 ;
      RECT MASK 1 72.445 97.41 72.505 108.838 ;
      RECT MASK 1 72.719 97.41 72.779 108.838 ;
      RECT MASK 1 72.993 97.41 73.053 108.838 ;
      RECT MASK 1 73.267 97.41 73.327 108.838 ;
      RECT MASK 1 73.541 97.41 73.601 108.838 ;
      RECT MASK 1 73.815 97.41 73.875 108.838 ;
      RECT MASK 1 74.089 97.41 74.149 108.838 ;
      RECT MASK 1 74.363 97.41 74.423 108.838 ;
      RECT MASK 1 74.637 97.41 74.697 108.838 ;
      RECT MASK 1 74.911 97.41 74.971 108.838 ;
      RECT MASK 1 75.185 97.41 75.245 108.838 ;
      RECT MASK 1 75.459 97.41 75.519 108.838 ;
      RECT MASK 1 75.733 97.41 75.793 108.838 ;
      RECT MASK 1 76.007 97.41 76.067 108.838 ;
      RECT MASK 1 76.281 97.41 76.341 108.838 ;
      RECT MASK 1 76.555 97.41 76.615 108.838 ;
      RECT MASK 1 76.829 97.41 76.889 108.838 ;
      RECT MASK 1 77.103 97.41 77.163 108.838 ;
      RECT MASK 1 77.377 97.41 77.437 108.838 ;
      RECT MASK 1 77.651 97.41 77.711 108.838 ;
      RECT MASK 1 77.925 97.41 77.985 108.838 ;
      RECT MASK 1 78.199 97.41 78.259 108.838 ;
      RECT MASK 1 78.473 97.41 78.533 108.838 ;
      RECT MASK 1 78.747 97.41 78.807 108.838 ;
      RECT MASK 1 79.021 97.41 79.081 108.838 ;
      RECT MASK 1 79.295 97.41 79.355 108.838 ;
      RECT MASK 1 79.569 97.41 79.629 108.838 ;
      RECT MASK 1 79.843 97.41 79.903 108.838 ;
      RECT MASK 1 80.117 97.41 80.177 108.838 ;
      RECT MASK 1 80.391 97.41 80.451 108.838 ;
      RECT MASK 1 80.665 97.41 80.725 108.838 ;
      RECT MASK 1 80.939 97.41 80.999 108.838 ;
      RECT MASK 1 81.213 97.41 81.273 108.838 ;
      RECT MASK 1 81.487 97.41 81.547 108.838 ;
      RECT MASK 1 81.761 97.41 81.821 108.838 ;
      RECT MASK 1 82.035 97.41 82.095 108.838 ;
      RECT MASK 1 82.309 97.41 82.369 108.838 ;
      RECT MASK 1 82.583 97.41 82.643 108.838 ;
      RECT MASK 1 82.857 97.41 82.917 108.838 ;
      RECT MASK 1 83.131 97.41 83.191 108.838 ;
      RECT MASK 1 83.405 97.41 83.465 108.838 ;
      RECT MASK 1 83.679 97.41 83.739 108.838 ;
      RECT MASK 1 83.953 97.41 84.013 108.838 ;
      RECT MASK 1 84.227 97.41 84.287 108.838 ;
      RECT MASK 1 84.501 97.41 84.561 108.838 ;
      RECT MASK 1 84.775 97.41 84.835 108.838 ;
      RECT MASK 1 85.049 97.41 85.109 108.838 ;
      RECT MASK 1 85.323 97.41 85.383 108.838 ;
      RECT MASK 1 85.597 97.41 85.657 108.838 ;
      RECT MASK 1 85.871 97.41 85.931 108.838 ;
      RECT MASK 1 86.145 97.41 86.205 108.838 ;
      RECT MASK 1 86.419 97.41 86.479 108.838 ;
      RECT MASK 1 86.693 97.41 86.753 108.838 ;
      RECT MASK 1 89.226 97.41 89.286 108.838 ;
      RECT MASK 1 89.5 97.41 89.56 108.838 ;
      RECT MASK 1 89.774 97.41 89.834 108.838 ;
      RECT MASK 1 90.048 97.41 90.108 108.838 ;
      RECT MASK 1 90.322 97.41 90.382 108.838 ;
      RECT MASK 1 90.596 97.41 90.656 108.838 ;
      RECT MASK 1 90.87 97.41 90.93 108.838 ;
      RECT MASK 1 91.144 97.41 91.204 108.838 ;
      RECT MASK 1 91.418 97.41 91.478 108.838 ;
      RECT MASK 1 91.692 97.41 91.752 108.838 ;
      RECT MASK 1 91.966 97.41 92.026 108.838 ;
      RECT MASK 1 92.24 97.41 92.3 108.838 ;
      RECT MASK 1 92.514 97.41 92.574 108.838 ;
      RECT MASK 1 92.788 97.41 92.848 108.838 ;
      RECT MASK 1 93.062 97.41 93.122 108.838 ;
      RECT MASK 1 93.336 97.41 93.396 108.838 ;
      RECT MASK 1 93.61 97.41 93.67 108.838 ;
      RECT MASK 1 93.884 97.41 93.944 108.838 ;
      RECT MASK 1 94.158 97.41 94.218 108.838 ;
      RECT MASK 1 94.432 97.41 94.492 108.838 ;
      RECT MASK 1 94.706 97.41 94.766 108.838 ;
      RECT MASK 1 94.98 97.41 95.04 108.838 ;
      RECT MASK 1 95.254 97.41 95.314 108.838 ;
      RECT MASK 1 95.528 97.41 95.588 108.838 ;
      RECT MASK 1 95.802 97.41 95.862 108.838 ;
      RECT MASK 1 96.076 97.41 96.136 108.838 ;
      RECT MASK 1 96.35 97.41 96.41 108.838 ;
      RECT MASK 1 96.624 97.41 96.684 108.838 ;
      RECT MASK 1 96.898 97.41 96.958 108.838 ;
      RECT MASK 1 97.172 97.41 97.232 108.838 ;
      RECT MASK 1 97.446 97.41 97.506 108.838 ;
      RECT MASK 1 97.72 97.41 97.78 108.838 ;
      RECT MASK 1 97.994 97.41 98.054 108.838 ;
      RECT MASK 1 98.268 97.41 98.328 108.838 ;
      RECT MASK 1 98.542 97.41 98.602 108.838 ;
      RECT MASK 1 98.816 97.41 98.876 108.838 ;
      RECT MASK 1 99.09 97.41 99.15 108.838 ;
      RECT MASK 1 99.364 97.41 99.424 108.838 ;
      RECT MASK 1 99.638 97.41 99.698 108.838 ;
      RECT MASK 1 99.912 97.41 99.972 108.838 ;
      RECT MASK 1 100.186 97.41 100.246 108.838 ;
      RECT MASK 1 100.46 97.41 100.52 108.838 ;
      RECT MASK 1 100.734 97.41 100.794 108.838 ;
      RECT MASK 1 101.008 97.41 101.068 108.838 ;
      RECT MASK 1 101.282 97.41 101.342 108.838 ;
      RECT MASK 1 101.556 97.41 101.616 108.838 ;
      RECT MASK 1 101.83 97.41 101.89 108.838 ;
      RECT MASK 1 102.104 97.41 102.164 108.838 ;
      RECT MASK 1 102.378 97.41 102.438 108.838 ;
      RECT MASK 1 102.652 97.41 102.712 108.838 ;
      RECT MASK 1 102.926 97.41 102.986 108.838 ;
      RECT MASK 1 103.2 97.41 103.26 108.838 ;
      RECT MASK 1 103.474 97.41 103.534 108.838 ;
      RECT MASK 1 103.748 97.41 103.808 108.838 ;
      RECT MASK 1 104.022 97.41 104.082 108.838 ;
      RECT MASK 1 104.296 97.41 104.356 108.838 ;
      RECT MASK 1 104.57 97.41 104.63 108.838 ;
      RECT MASK 1 104.844 97.41 104.904 108.838 ;
      RECT MASK 1 105.118 97.41 105.178 108.838 ;
      RECT MASK 1 105.392 97.41 105.452 108.838 ;
      RECT MASK 1 105.666 97.41 105.726 108.838 ;
      RECT MASK 1 105.94 97.41 106 108.838 ;
      RECT MASK 1 106.214 97.41 106.274 108.838 ;
      RECT MASK 1 106.488 97.41 106.548 108.838 ;
      RECT MASK 1 106.762 97.41 106.822 108.838 ;
      RECT MASK 1 107.036 97.41 107.096 108.838 ;
      RECT MASK 1 107.31 97.41 107.37 108.838 ;
      RECT MASK 1 107.584 97.41 107.644 108.838 ;
      RECT MASK 1 107.858 97.41 107.918 108.838 ;
      RECT MASK 1 108.132 97.41 108.192 108.838 ;
      RECT MASK 1 108.406 97.41 108.466 108.838 ;
      RECT MASK 1 108.68 97.41 108.74 108.838 ;
      RECT MASK 1 108.954 97.41 109.014 108.838 ;
      RECT MASK 1 109.228 97.41 109.288 108.838 ;
      RECT MASK 1 109.502 97.41 109.562 108.838 ;
      RECT MASK 1 109.776 97.41 109.836 108.838 ;
      RECT MASK 1 110.05 97.41 110.11 108.838 ;
      RECT MASK 1 110.324 97.41 110.384 108.838 ;
      RECT MASK 1 110.598 97.41 110.658 108.838 ;
      RECT MASK 1 110.872 97.41 110.932 108.838 ;
      RECT MASK 1 111.146 97.41 111.206 108.838 ;
      RECT MASK 1 111.42 97.41 111.48 108.838 ;
      RECT MASK 1 111.694 97.41 111.754 108.838 ;
      RECT MASK 1 111.968 97.41 112.028 108.838 ;
      RECT MASK 1 112.242 97.41 112.302 108.838 ;
      RECT MASK 1 112.516 97.41 112.576 108.838 ;
      RECT MASK 1 112.79 97.41 112.85 108.838 ;
      RECT MASK 1 113.064 97.41 113.124 108.838 ;
      RECT MASK 1 113.338 97.41 113.398 108.838 ;
      RECT MASK 1 113.612 97.41 113.672 108.838 ;
      RECT MASK 1 113.886 97.41 113.946 108.838 ;
      RECT MASK 1 114.16 97.41 114.22 108.838 ;
      RECT MASK 1 114.434 97.41 114.494 108.838 ;
      RECT MASK 1 114.708 97.41 114.768 108.838 ;
      RECT MASK 1 114.982 97.41 115.042 108.838 ;
      RECT MASK 1 115.256 97.41 115.316 108.838 ;
      RECT MASK 1 115.53 97.41 115.59 108.838 ;
      RECT MASK 1 115.804 97.41 115.864 108.838 ;
      RECT MASK 1 116.078 97.41 116.138 108.838 ;
      RECT MASK 1 116.352 97.41 116.412 108.838 ;
      RECT MASK 1 116.626 97.41 116.686 108.838 ;
      RECT MASK 1 116.9 97.41 116.96 108.838 ;
      RECT MASK 1 117.174 97.41 117.234 108.838 ;
      RECT MASK 1 117.448 97.41 117.508 108.838 ;
      RECT MASK 1 117.722 97.41 117.782 108.838 ;
      RECT MASK 1 117.996 97.41 118.056 108.838 ;
      RECT MASK 1 118.27 97.41 118.33 108.838 ;
      RECT MASK 1 118.544 97.41 118.604 108.838 ;
      RECT MASK 1 118.818 97.41 118.878 108.838 ;
      RECT MASK 1 119.092 97.41 119.152 108.838 ;
      RECT MASK 1 119.366 97.41 119.426 108.838 ;
      RECT MASK 1 119.64 97.41 119.7 108.838 ;
      RECT MASK 1 119.914 97.41 119.974 108.838 ;
      RECT MASK 1 120.188 97.41 120.248 108.838 ;
      RECT MASK 1 120.462 97.41 120.522 108.838 ;
      RECT MASK 1 120.736 97.41 120.796 108.838 ;
      RECT MASK 1 121.01 97.41 121.07 108.838 ;
      RECT MASK 1 121.284 97.41 121.344 108.838 ;
      RECT MASK 1 121.558 97.41 121.618 108.838 ;
      RECT MASK 1 121.832 97.41 121.892 108.838 ;
      RECT MASK 1 122.106 97.41 122.166 108.838 ;
      RECT MASK 1 122.38 97.41 122.44 108.838 ;
      RECT MASK 1 122.654 97.41 122.714 108.838 ;
      RECT MASK 1 122.928 97.41 122.988 108.838 ;
      RECT MASK 1 123.202 97.41 123.262 108.838 ;
      RECT MASK 1 123.476 97.41 123.536 108.838 ;
      RECT MASK 1 123.75 97.41 123.81 108.838 ;
      RECT MASK 1 124.024 97.41 124.084 108.838 ;
      RECT MASK 1 124.298 97.41 124.358 108.838 ;
      RECT MASK 1 124.572 97.41 124.632 108.838 ;
      RECT MASK 1 124.846 97.41 124.906 108.838 ;
      RECT MASK 1 125.12 97.41 125.18 108.838 ;
      RECT MASK 1 125.394 97.41 125.454 108.838 ;
      RECT MASK 1 125.668 97.41 125.728 108.838 ;
      RECT MASK 1 125.942 97.41 126.002 108.838 ;
      RECT MASK 1 126.216 97.41 126.276 108.838 ;
      RECT MASK 1 126.49 97.41 126.55 108.838 ;
      RECT MASK 1 126.764 97.41 126.824 108.838 ;
      RECT MASK 1 127.038 97.41 127.098 108.838 ;
      RECT MASK 1 127.312 97.41 127.372 108.838 ;
      RECT MASK 2 1.878 0.51 1.998 18.09 ;
      RECT MASK 2 2.256 0.51 2.376 18.09 ;
      RECT MASK 2 2.634 0.51 2.754 18.09 ;
      RECT MASK 2 3.012 0.51 3.132 18.09 ;
      RECT MASK 2 3.39 0.51 3.51 18.09 ;
      RECT MASK 2 3.768 0.51 3.888 18.09 ;
      RECT MASK 2 4.146 0.51 4.266 17.85 ;
      RECT MASK 2 4.524 0.51 4.644 10.77 ;
      RECT MASK 2 4.902 0.51 5.022 17.85 ;
      RECT MASK 2 5.28 0.51 5.4 10.77 ;
      RECT MASK 2 5.658 0.51 5.778 17.85 ;
      RECT MASK 2 6.036 0.51 6.156 10.77 ;
      RECT MASK 2 6.414 0.51 6.534 17.85 ;
      RECT MASK 2 6.82 0.51 6.94 17.85 ;
      RECT MASK 2 7.198 0.51 7.318 10.77 ;
      RECT MASK 2 7.576 0.51 7.696 17.85 ;
      RECT MASK 2 7.982 0.51 8.102 17.85 ;
      RECT MASK 2 8.36 0.51 8.48 10.77 ;
      RECT MASK 2 8.738 0.51 8.858 17.85 ;
      RECT MASK 2 9.144 0.51 9.264 17.85 ;
      RECT MASK 2 9.522 0.51 9.642 10.77 ;
      RECT MASK 2 9.9 0.51 10.02 17.85 ;
      RECT MASK 2 11.142 0.51 11.262 10.77 ;
      RECT MASK 2 11.52 0.51 11.64 17.85 ;
      RECT MASK 2 11.898 0.51 12.018 10.77 ;
      RECT MASK 2 12.276 0.51 12.396 17.85 ;
      RECT MASK 2 12.654 0.51 12.774 10.77 ;
      RECT MASK 2 13.032 0.51 13.152 17.85 ;
      RECT MASK 2 13.438 0.51 13.558 17.85 ;
      RECT MASK 2 14.194 0.51 14.314 17.85 ;
      RECT MASK 2 14.6 0.51 14.72 17.85 ;
      RECT MASK 2 15.356 0.51 15.476 14.322 ;
      RECT MASK 2 15.762 0.51 15.882 17.85 ;
      RECT MASK 2 16.518 0.51 16.638 17.85 ;
      RECT MASK 2 17.382 0.51 17.502 17.85 ;
      RECT MASK 2 18.138 0.51 18.258 14.4415 ;
      RECT MASK 2 18.894 0.51 19.014 17.85 ;
      RECT MASK 2 19.65 0.51 19.77 17.85 ;
      RECT MASK 2 20.056 0.51 20.176 17.85 ;
      RECT MASK 2 20.812 0.51 20.932 17.85 ;
      RECT MASK 2 21.218 0.51 21.338 17.85 ;
      RECT MASK 2 21.596 0.51 21.716 17.85 ;
      RECT MASK 2 22.38 0.51 22.5 17.82 ;
      RECT MASK 2 23.136 0.51 23.256 17.82 ;
      RECT MASK 2 23.622 0.51 23.742 11.1545 ;
      RECT MASK 2 24.378 0.51 24.498 11.1545 ;
      RECT MASK 2 24.756 0.51 24.876 17.85 ;
      RECT MASK 2 25.134 0.51 25.254 11.1545 ;
      RECT MASK 2 25.512 0.51 25.632 17.85 ;
      RECT MASK 2 26.268 0.51 26.388 17.85 ;
      RECT MASK 2 26.674 0.51 26.794 17.85 ;
      RECT MASK 2 27.052 0.51 27.172 11.1545 ;
      RECT MASK 2 27.43 0.51 27.55 17.85 ;
      RECT MASK 2 27.836 0.51 27.956 17.85 ;
      RECT MASK 2 28.214 0.51 28.334 11.1545 ;
      RECT MASK 2 28.592 0.51 28.712 14.322 ;
      RECT MASK 2 28.998 0.51 29.118 17.85 ;
      RECT MASK 2 29.376 0.51 29.496 11.1545 ;
      RECT MASK 2 29.754 0.51 29.874 17.85 ;
      RECT MASK 2 30.24 0.51 30.36 11.1545 ;
      RECT MASK 2 30.618 0.51 30.738 14.387 ;
      RECT MASK 2 30.996 0.51 31.116 9.1675 ;
      RECT MASK 2 31.374 0.51 31.494 9.1675 ;
      RECT MASK 2 31.752 0.51 31.872 9.1675 ;
      RECT MASK 2 32.13 0.51 32.25 17.85 ;
      RECT MASK 2 32.508 0.51 32.628 8.291 ;
      RECT MASK 2 32.886 0.51 33.006 17.85 ;
      RECT MASK 2 33.292 0.51 33.412 8.291 ;
      RECT MASK 2 33.67 0.51 33.79 10.77 ;
      RECT MASK 2 34.048 0.51 34.168 8.291 ;
      RECT MASK 2 34.454 0.51 34.574 17.85 ;
      RECT MASK 2 34.832 0.51 34.952 8.291 ;
      RECT MASK 2 35.21 0.51 35.33 17.85 ;
      RECT MASK 2 35.588 0.51 35.708 8.094 ;
      RECT MASK 2 35.994 0.51 36.114 10.77 ;
      RECT MASK 2 36.372 0.51 36.492 8.094 ;
      RECT MASK 2 36.858 0.51 36.978 8.291 ;
      RECT MASK 2 37.236 0.51 37.356 17.85 ;
      RECT MASK 2 37.614 0.51 37.734 8.291 ;
      RECT MASK 2 37.992 0.51 38.112 17.85 ;
      RECT MASK 2 38.37 0.51 38.49 8.291 ;
      RECT MASK 2 38.748 0.51 38.868 17.82 ;
      RECT MASK 2 39.126 0.51 39.246 8.291 ;
      RECT MASK 2 39.504 0.51 39.624 17.82 ;
      RECT MASK 2 39.91 0.51 40.03 17.85 ;
      RECT MASK 2 40.288 0.51 40.408 8.291 ;
      RECT MASK 2 40.666 0.51 40.786 17.85 ;
      RECT MASK 2 41.072 0.51 41.192 17.82 ;
      RECT MASK 2 41.45 0.51 41.57 8.291 ;
      RECT MASK 2 42.1535 0.51 42.2735 3.935 ;
      RECT MASK 2 42.612 0.51 42.732 8.291 ;
      RECT MASK 2 42.99 0.51 43.11 17.85 ;
      RECT MASK 2 43.854 0.51 43.974 14.322 ;
      RECT MASK 2 44.232 0.51 44.352 8.291 ;
      RECT MASK 2 44.61 0.51 44.73 17.85 ;
      RECT MASK 2 44.988 0.51 45.108 8.291 ;
      RECT MASK 2 45.366 0.51 45.486 17.85 ;
      RECT MASK 2 45.744 0.51 45.864 8.291 ;
      RECT MASK 2 46.122 0.51 46.242 17.85 ;
      RECT MASK 2 46.5 0.51 46.62 4.5 ;
      RECT MASK 2 46.878 0.51 46.998 10.77 ;
      RECT MASK 2 47.284 0.51 47.404 4.5 ;
      RECT MASK 2 47.662 0.51 47.782 10.77 ;
      RECT MASK 2 48.04 0.51 48.16 4.5 ;
      RECT MASK 2 48.446 0.51 48.566 17.82 ;
      RECT MASK 2 48.824 0.51 48.944 4.5 ;
      RECT MASK 2 49.986 0.51 50.106 1.5195 ;
      RECT MASK 2 50.472 0.51 50.592 17.85 ;
      RECT MASK 2 50.85 0.51 50.97 1.5195 ;
      RECT MASK 2 51.228 0.51 51.348 17.85 ;
      RECT MASK 2 51.606 0.51 51.726 1.5195 ;
      RECT MASK 2 51.984 0.51 52.104 17.82 ;
      RECT MASK 2 52.362 0.51 52.482 1.5195 ;
      RECT MASK 2 53.524 0.51 53.644 17.85 ;
      RECT MASK 2 53.874 0.51 53.994 10.77 ;
      RECT MASK 2 54.308 0.51 54.428 10.77 ;
      RECT MASK 2 54.686 0.51 54.806 10.77 ;
      RECT MASK 2 55.064 0.51 55.184 10.77 ;
      RECT MASK 2 55.47 0.51 55.59 17.85 ;
      RECT MASK 2 55.848 0.51 55.968 17.85 ;
      RECT MASK 2 56.226 0.51 56.346 17.85 ;
      RECT MASK 2 57.846 0.51 57.966 17.85 ;
      RECT MASK 2 58.224 0.51 58.344 22.36 ;
      RECT MASK 2 59.358 0.51 59.478 17.85 ;
      RECT MASK 2 60.52 0.51 60.64 17.85 ;
      RECT MASK 2 60.926 0.51 61.046 17.85 ;
      RECT MASK 2 61.304 0.51 61.424 10.4 ;
      RECT MASK 2 61.682 0.51 61.802 1.302 ;
      RECT MASK 2 62.088 0.51 62.208 10.4 ;
      RECT MASK 2 63.33 0.51 63.45 10.4 ;
      RECT MASK 2 64.086 0.51 64.206 1.3965 ;
      RECT MASK 2 64.464 0.51 64.584 10.4 ;
      RECT MASK 2 65.22 0.51 65.34 10.4 ;
      RECT MASK 2 65.598 0.51 65.718 10.56 ;
      RECT MASK 2 65.976 0.51 66.096 10.4 ;
      RECT MASK 2 67.544 0.51 67.664 10.4 ;
      RECT MASK 2 67.922 0.51 68.042 10.56 ;
      RECT MASK 2 68.3 0.51 68.42 10.4 ;
      RECT MASK 2 68.706 0.51 68.826 14.322 ;
      RECT MASK 2 69.084 0.51 69.204 10.4 ;
      RECT MASK 2 69.462 0.51 69.582 17.85 ;
      RECT MASK 2 69.948 0.51 70.068 10.4 ;
      RECT MASK 2 70.326 0.51 70.446 10.56 ;
      RECT MASK 2 70.704 0.51 70.824 10.4 ;
      RECT MASK 2 73.756 0.51 73.876 17.85 ;
      RECT MASK 2 74.162 0.51 74.282 17.85 ;
      RECT MASK 2 74.918 0.51 75.038 17.85 ;
      RECT MASK 2 75.324 0.51 75.444 17.85 ;
      RECT MASK 2 76.08 0.51 76.2 17.85 ;
      RECT MASK 2 76.944 0.51 77.064 17.85 ;
      RECT MASK 2 77.7 0.51 77.82 17.85 ;
      RECT MASK 2 78.456 0.51 78.576 17.85 ;
      RECT MASK 2 79.212 0.51 79.332 17.85 ;
      RECT MASK 2 79.618 0.51 79.738 17.85 ;
      RECT MASK 2 80.374 0.51 80.494 14.3385 ;
      RECT MASK 2 80.78 0.51 80.9 10.77 ;
      RECT MASK 2 81.158 0.51 81.278 10.77 ;
      RECT MASK 2 81.536 0.51 81.656 10.77 ;
      RECT MASK 2 81.942 0.51 82.062 14.379 ;
      RECT MASK 2 82.32 0.51 82.44 10.77 ;
      RECT MASK 2 82.698 0.51 82.818 17.85 ;
      RECT MASK 2 83.076 0.51 83.196 10.77 ;
      RECT MASK 2 83.562 0.51 83.682 17.85 ;
      RECT MASK 2 83.94 0.51 84.06 10.77 ;
      RECT MASK 2 84.318 0.51 84.438 17.85 ;
      RECT MASK 2 84.696 0.51 84.816 10.77 ;
      RECT MASK 2 85.074 0.51 85.194 17.85 ;
      RECT MASK 2 85.452 0.51 85.572 10.77 ;
      RECT MASK 2 85.83 0.51 85.95 17.85 ;
      RECT MASK 2 86.236 0.51 86.356 10.77 ;
      RECT MASK 2 86.614 0.51 86.734 10.77 ;
      RECT MASK 2 86.992 0.51 87.112 10.77 ;
      RECT MASK 2 87.398 0.51 87.518 17.85 ;
      RECT MASK 2 87.776 0.51 87.896 10.77 ;
      RECT MASK 2 88.154 0.51 88.274 17.85 ;
      RECT MASK 2 88.56 0.51 88.68 10.77 ;
      RECT MASK 2 88.938 0.51 89.058 10.77 ;
      RECT MASK 2 89.316 0.51 89.436 10.77 ;
      RECT MASK 2 89.802 0.51 89.922 10.77 ;
      RECT MASK 2 90.18 0.51 90.3 10.77 ;
      RECT MASK 2 90.558 0.51 90.678 10.77 ;
      RECT MASK 2 90.936 0.51 91.056 10.77 ;
      RECT MASK 2 91.314 0.51 91.434 10.77 ;
      RECT MASK 2 91.692 0.51 91.812 10.77 ;
      RECT MASK 2 92.07 0.51 92.19 10.77 ;
      RECT MASK 2 92.448 0.51 92.568 17.85 ;
      RECT MASK 2 92.854 0.51 92.974 17.85 ;
      RECT MASK 2 93.61 0.51 93.73 14.322 ;
      RECT MASK 2 94.016 0.51 94.136 17.85 ;
      RECT MASK 2 94.772 0.51 94.892 17.85 ;
      RECT MASK 2 95.178 0.51 95.298 17.85 ;
      RECT MASK 2 95.556 0.51 95.676 10.77 ;
      RECT MASK 2 95.934 0.51 96.054 17.85 ;
      RECT MASK 2 96.42 0.51 96.54 10.77 ;
      RECT MASK 2 96.798 0.51 96.918 17.85 ;
      RECT MASK 2 97.176 0.51 97.296 10.77 ;
      RECT MASK 2 97.554 0.51 97.674 14.322 ;
      RECT MASK 2 97.932 0.51 98.052 10.77 ;
      RECT MASK 2 98.31 0.51 98.43 17.85 ;
      RECT MASK 2 98.688 0.51 98.808 10.77 ;
      RECT MASK 2 99.066 0.51 99.186 17.85 ;
      RECT MASK 2 99.472 0.51 99.592 10.77 ;
      RECT MASK 2 99.85 0.51 99.97 10.77 ;
      RECT MASK 2 100.228 0.51 100.348 10.77 ;
      RECT MASK 2 100.634 0.51 100.754 17.85 ;
      RECT MASK 2 101.012 0.51 101.132 10.77 ;
      RECT MASK 2 101.39 0.51 101.51 17.85 ;
      RECT MASK 2 101.796 0.51 101.916 10.77 ;
      RECT MASK 2 102.174 0.51 102.294 10.77 ;
      RECT MASK 2 102.552 0.51 102.672 10.77 ;
      RECT MASK 2 103.038 0.51 103.158 10.77 ;
      RECT MASK 2 103.416 0.51 103.536 10.77 ;
      RECT MASK 2 103.794 0.51 103.914 10.77 ;
      RECT MASK 2 104.172 0.51 104.292 10.77 ;
      RECT MASK 2 104.55 0.51 104.67 10.77 ;
      RECT MASK 2 104.928 0.51 105.048 10.77 ;
      RECT MASK 2 105.306 0.51 105.426 10.77 ;
      RECT MASK 2 105.684 0.51 105.804 10.77 ;
      RECT MASK 2 106.09 0.51 106.21 10.77 ;
      RECT MASK 2 106.468 0.51 106.588 10.77 ;
      RECT MASK 2 106.846 0.51 106.966 14.322 ;
      RECT MASK 2 107.252 0.51 107.372 17.85 ;
      RECT MASK 2 108.008 0.51 108.128 10.77 ;
      RECT MASK 2 108.414 0.51 108.534 17.85 ;
      RECT MASK 2 109.17 0.51 109.29 17.85 ;
      RECT MASK 2 110.034 0.51 110.154 17.85 ;
      RECT MASK 2 110.79 0.51 110.91 17.85 ;
      RECT MASK 2 111.546 0.51 111.666 17.85 ;
      RECT MASK 2 111.924 0.51 112.044 17.85 ;
      RECT MASK 2 112.302 0.51 112.422 17.85 ;
      RECT MASK 2 112.68 0.51 112.8 17.85 ;
      RECT MASK 2 113.058 0.51 113.178 17.85 ;
      RECT MASK 2 113.436 0.51 113.556 17.85 ;
      RECT MASK 2 113.814 0.51 113.934 17.85 ;
      RECT MASK 2 24.0385 0.935 24.0985 4.825 ;
      RECT MASK 2 22.2 1.135 22.26 9.3965 ;
      RECT MASK 2 62.7385 1.299 62.8585 3.0225 ;
      RECT MASK 2 63.57 1.299 63.63 3.0225 ;
      RECT MASK 2 64.871 1.319 64.951 3.0225 ;
      RECT MASK 2 58.794 1.64 58.854 3.04 ;
      RECT MASK 2 61.566 1.64 61.626 3.28 ;
      RECT MASK 2 63.834 1.64 63.894 3.04 ;
      RECT MASK 2 116.291 1.6565 116.351 23.6505 ;
      RECT MASK 2 116.565 1.6565 116.625 23.6505 ;
      RECT MASK 2 116.839 1.6565 116.899 23.6505 ;
      RECT MASK 2 117.113 1.6565 117.173 23.6505 ;
      RECT MASK 2 117.387 1.6565 117.447 23.6505 ;
      RECT MASK 2 117.661 1.6565 117.721 23.6505 ;
      RECT MASK 2 117.935 1.6565 117.995 23.6505 ;
      RECT MASK 2 118.209 1.6565 118.269 23.6505 ;
      RECT MASK 2 118.483 1.6565 118.543 23.6505 ;
      RECT MASK 2 118.757 1.6565 118.817 23.6505 ;
      RECT MASK 2 119.031 1.6565 119.091 23.6505 ;
      RECT MASK 2 119.305 1.6565 119.365 23.6505 ;
      RECT MASK 2 119.579 1.6565 119.639 23.6505 ;
      RECT MASK 2 119.853 1.6565 119.913 23.6505 ;
      RECT MASK 2 120.127 1.6565 120.187 23.6505 ;
      RECT MASK 2 120.401 1.6565 120.461 23.6505 ;
      RECT MASK 2 120.675 1.6565 120.735 23.6505 ;
      RECT MASK 2 120.949 1.6565 121.009 23.6505 ;
      RECT MASK 2 121.223 1.6565 121.283 23.6505 ;
      RECT MASK 2 121.497 1.6565 121.557 23.6505 ;
      RECT MASK 2 121.771 1.6565 121.831 23.6505 ;
      RECT MASK 2 122.045 1.6565 122.105 23.6505 ;
      RECT MASK 2 122.319 1.6565 122.379 23.6505 ;
      RECT MASK 2 122.593 1.6565 122.653 23.6505 ;
      RECT MASK 2 122.867 1.6565 122.927 23.6505 ;
      RECT MASK 2 123.141 1.6565 123.201 23.6505 ;
      RECT MASK 2 123.415 1.6565 123.475 23.6505 ;
      RECT MASK 2 123.689 1.6565 123.749 23.6505 ;
      RECT MASK 2 123.963 1.6565 124.023 23.6505 ;
      RECT MASK 2 124.237 1.6565 124.297 23.6505 ;
      RECT MASK 2 124.511 1.6565 124.571 23.6505 ;
      RECT MASK 2 124.785 1.6565 124.845 23.6505 ;
      RECT MASK 2 125.059 1.6565 125.119 23.6505 ;
      RECT MASK 2 125.333 1.6565 125.393 23.6505 ;
      RECT MASK 2 125.607 1.6565 125.667 23.6505 ;
      RECT MASK 2 125.881 1.6565 125.941 23.6505 ;
      RECT MASK 2 126.155 1.6565 126.215 23.6505 ;
      RECT MASK 2 126.429 1.6565 126.489 23.6505 ;
      RECT MASK 2 126.703 1.6565 126.763 23.6505 ;
      RECT MASK 2 126.977 1.6565 127.037 23.6505 ;
      RECT MASK 2 127.251 1.6565 127.311 10.8495 ;
      RECT MASK 2 127.525 1.6565 127.585 10.8495 ;
      RECT MASK 2 127.799 1.6565 127.859 10.952 ;
      RECT MASK 2 22.956 2.861 23.016 6.57 ;
      RECT MASK 2 10.3885 3.03 10.5085 6.629 ;
      RECT MASK 2 56.712 3.1155 56.832 22.36 ;
      RECT MASK 2 57.09 3.1155 57.21 10.898 ;
      RECT MASK 2 57.468 3.1155 57.588 22.36 ;
      RECT MASK 2 58.98 3.12 59.1 84.25 ;
      RECT MASK 2 63.035 3.4905 63.155 4.5015 ;
      RECT MASK 2 58.602 3.51 58.722 4.6475 ;
      RECT MASK 2 42.1835 4.495 42.2435 8.384 ;
      RECT MASK 2 61.566 4.88 61.626 6.52 ;
      RECT MASK 2 46.5 4.95 46.62 10.77 ;
      RECT MASK 2 47.284 4.95 47.404 10.77 ;
      RECT MASK 2 48.04 4.95 48.16 10.77 ;
      RECT MASK 2 48.824 4.95 48.944 10.77 ;
      RECT MASK 2 58.794 5.12 58.854 6.52 ;
      RECT MASK 2 63.834 5.12 63.894 6.52 ;
      RECT MASK 2 24 5.1645 24.12 17.85 ;
      RECT MASK 2 64.867 5.213 64.947 10.575 ;
      RECT MASK 2 62.814 5.2165 62.894 10.575 ;
      RECT MASK 2 63.1095 5.2165 63.1895 10.575 ;
      RECT MASK 2 49.986 6.2695 50.106 10.77 ;
      RECT MASK 2 50.85 6.2695 50.97 10.77 ;
      RECT MASK 2 51.606 6.2695 51.726 17.85 ;
      RECT MASK 2 52.362 6.2695 52.482 17.82 ;
      RECT MASK 2 22.782 6.8415 22.862 10.9305 ;
      RECT MASK 2 42.0045 6.8675 42.0645 8.283 ;
      RECT MASK 2 58.794 7.88 58.854 9.28 ;
      RECT MASK 2 61.566 7.88 61.626 9.52 ;
      RECT MASK 2 63.834 7.88 63.894 9.28 ;
      RECT MASK 2 45.744 8.86 45.864 17.85 ;
      RECT MASK 2 36.858 8.9095 36.978 17.85 ;
      RECT MASK 2 37.614 8.9095 37.734 14.328 ;
      RECT MASK 2 38.37 8.9095 38.49 17.85 ;
      RECT MASK 2 39.126 8.9095 39.246 17.82 ;
      RECT MASK 2 40.288 8.9095 40.408 17.82 ;
      RECT MASK 2 44.232 8.9095 44.352 14.322 ;
      RECT MASK 2 44.988 8.9095 45.108 17.85 ;
      RECT MASK 2 32.508 8.91 32.628 17.85 ;
      RECT MASK 2 33.292 8.91 33.412 10.77 ;
      RECT MASK 2 34.048 8.91 34.168 10.77 ;
      RECT MASK 2 34.832 8.91 34.952 17.85 ;
      RECT MASK 2 35.616 8.91 35.736 10.77 ;
      RECT MASK 2 36.372 8.91 36.492 10.77 ;
      RECT MASK 2 53.009 9.325 53.069 10.845 ;
      RECT MASK 2 31.257 9.482 31.317 10.6735 ;
      RECT MASK 2 21.974 9.5605 22.094 17.85 ;
      RECT MASK 2 30.9355 9.684 30.9955 10.4715 ;
      RECT MASK 2 60.167 10.22 60.247 16.66 ;
      RECT MASK 2 31.7635 10.732 31.8235 11.0495 ;
      RECT MASK 2 127.358 11.063 127.478 76.891 ;
      RECT MASK 2 33.67 11.178 33.79 17.82 ;
      RECT MASK 2 35.994 11.178 36.114 17.82 ;
      RECT MASK 2 31.374 11.2745 31.494 17.85 ;
      RECT MASK 2 31.752 11.2745 31.872 17.85 ;
      RECT MASK 2 42.234 11.2745 42.354 17.85 ;
      RECT MASK 2 22.758 11.354 22.878 17.82 ;
      RECT MASK 2 25.89 11.354 26.01 17.82 ;
      RECT MASK 2 62.844 11.42 62.964 17.82 ;
      RECT MASK 2 63.708 11.42 63.828 17.85 ;
      RECT MASK 2 64.464 11.42 64.584 17.85 ;
      RECT MASK 2 65.22 11.42 65.34 18.137 ;
      RECT MASK 2 65.976 11.42 66.096 18.137 ;
      RECT MASK 2 66.382 11.42 66.502 18.137 ;
      RECT MASK 2 67.544 11.42 67.664 17.82 ;
      RECT MASK 2 68.3 11.42 68.42 17.82 ;
      RECT MASK 2 28.214 11.4705 28.334 17.82 ;
      RECT MASK 2 23.622 11.5145 23.742 17.85 ;
      RECT MASK 2 24.378 11.5145 24.498 17.85 ;
      RECT MASK 2 25.134 11.5145 25.254 17.85 ;
      RECT MASK 2 27.052 11.5145 27.172 17.82 ;
      RECT MASK 2 50.875 11.566 50.955 12.857 ;
      RECT MASK 2 53.062 11.566 53.142 13.814 ;
      RECT MASK 2 53.952 11.566 54.032 13.876 ;
      RECT MASK 2 4.524 11.67 4.644 17.85 ;
      RECT MASK 2 5.28 11.67 5.4 21.565 ;
      RECT MASK 2 6.036 11.67 6.156 26.01 ;
      RECT MASK 2 7.198 11.67 7.318 84.1645 ;
      RECT MASK 2 8.36 11.67 8.48 84.1645 ;
      RECT MASK 2 9.522 11.67 9.642 84.1645 ;
      RECT MASK 2 10.386 11.67 10.506 17.85 ;
      RECT MASK 2 10.764 11.67 10.884 17.85 ;
      RECT MASK 2 11.142 11.67 11.262 17.85 ;
      RECT MASK 2 11.898 11.67 12.018 17.85 ;
      RECT MASK 2 12.654 11.67 12.774 17.82 ;
      RECT MASK 2 13.816 11.67 13.936 17.82 ;
      RECT MASK 2 14.978 11.67 15.098 17.82 ;
      RECT MASK 2 16.14 11.67 16.26 17.82 ;
      RECT MASK 2 17.004 11.67 17.124 17.85 ;
      RECT MASK 2 17.76 11.67 17.88 17.85 ;
      RECT MASK 2 18.516 11.67 18.636 17.85 ;
      RECT MASK 2 19.272 11.67 19.392 17.82 ;
      RECT MASK 2 20.434 11.67 20.554 17.82 ;
      RECT MASK 2 29.376 11.67 29.496 17.82 ;
      RECT MASK 2 30.24 11.67 30.36 17.85 ;
      RECT MASK 2 30.996 11.67 31.116 17.85 ;
      RECT MASK 2 33.292 11.67 33.412 17.82 ;
      RECT MASK 2 34.048 11.67 34.168 17.82 ;
      RECT MASK 2 35.616 11.67 35.736 17.82 ;
      RECT MASK 2 36.372 11.67 36.492 17.82 ;
      RECT MASK 2 42.612 11.67 42.732 17.82 ;
      RECT MASK 2 43.476 11.67 43.596 17.85 ;
      RECT MASK 2 46.528 11.67 46.648 17.82 ;
      RECT MASK 2 46.906 11.67 47.026 17.82 ;
      RECT MASK 2 47.284 11.67 47.404 17.82 ;
      RECT MASK 2 47.69 11.67 47.81 17.85 ;
      RECT MASK 2 48.068 11.67 48.188 17.85 ;
      RECT MASK 2 48.852 11.67 48.972 17.82 ;
      RECT MASK 2 49.23 11.67 49.35 17.82 ;
      RECT MASK 2 49.608 11.67 49.728 17.82 ;
      RECT MASK 2 50.094 11.67 50.214 17.85 ;
      RECT MASK 2 54.308 11.67 54.428 17.82 ;
      RECT MASK 2 54.686 11.67 54.806 17.82 ;
      RECT MASK 2 55.064 11.67 55.184 14.322 ;
      RECT MASK 2 57.09 11.67 57.21 17.85 ;
      RECT MASK 2 58.602 11.67 58.722 17.82 ;
      RECT MASK 2 59.764 11.67 59.884 17.85 ;
      RECT MASK 2 61.304 11.67 61.424 84.25 ;
      RECT MASK 2 61.682 11.67 61.802 17.82 ;
      RECT MASK 2 62.088 11.67 62.208 17.82 ;
      RECT MASK 2 62.466 11.67 62.586 84.25 ;
      RECT MASK 2 63.33 11.67 63.45 17.85 ;
      RECT MASK 2 64.086 11.67 64.206 17.85 ;
      RECT MASK 2 64.842 11.67 64.962 17.85 ;
      RECT MASK 2 65.598 11.67 65.718 17.82 ;
      RECT MASK 2 66.76 11.67 66.88 17.82 ;
      RECT MASK 2 67.138 11.67 67.258 14.322 ;
      RECT MASK 2 67.922 11.67 68.042 17.82 ;
      RECT MASK 2 69.084 11.67 69.204 17.82 ;
      RECT MASK 2 69.948 11.67 70.068 17.85 ;
      RECT MASK 2 70.326 11.67 70.446 17.85 ;
      RECT MASK 2 70.704 11.67 70.824 17.85 ;
      RECT MASK 2 71.082 11.67 71.202 17.85 ;
      RECT MASK 2 71.46 11.67 71.58 17.85 ;
      RECT MASK 2 71.838 11.67 71.958 17.82 ;
      RECT MASK 2 72.216 11.67 72.336 17.82 ;
      RECT MASK 2 72.594 11.67 72.714 17.82 ;
      RECT MASK 2 73 11.67 73.12 17.82 ;
      RECT MASK 2 73.378 11.67 73.498 17.82 ;
      RECT MASK 2 74.54 11.67 74.66 17.82 ;
      RECT MASK 2 75.702 11.67 75.822 17.82 ;
      RECT MASK 2 76.566 11.67 76.686 17.85 ;
      RECT MASK 2 77.322 11.67 77.442 17.85 ;
      RECT MASK 2 78.078 11.67 78.198 17.85 ;
      RECT MASK 2 78.834 11.67 78.954 17.82 ;
      RECT MASK 2 79.996 11.67 80.116 17.82 ;
      RECT MASK 2 80.78 11.67 80.9 17.82 ;
      RECT MASK 2 81.536 11.67 81.656 17.82 ;
      RECT MASK 2 82.32 11.67 82.44 17.82 ;
      RECT MASK 2 83.94 11.67 84.06 14.441 ;
      RECT MASK 2 84.696 11.67 84.816 17.85 ;
      RECT MASK 2 85.452 11.67 85.572 17.82 ;
      RECT MASK 2 86.236 11.67 86.356 17.82 ;
      RECT MASK 2 86.614 11.67 86.734 17.82 ;
      RECT MASK 2 86.992 11.67 87.112 17.82 ;
      RECT MASK 2 87.776 11.67 87.896 17.82 ;
      RECT MASK 2 88.56 11.67 88.68 17.82 ;
      RECT MASK 2 88.938 11.67 89.058 17.82 ;
      RECT MASK 2 89.316 11.67 89.436 17.82 ;
      RECT MASK 2 89.802 11.67 89.922 17.85 ;
      RECT MASK 2 90.18 11.67 90.3 17.85 ;
      RECT MASK 2 90.558 11.67 90.678 17.85 ;
      RECT MASK 2 91.314 11.67 91.434 17.85 ;
      RECT MASK 2 91.692 11.67 91.812 17.82 ;
      RECT MASK 2 92.07 11.67 92.19 17.82 ;
      RECT MASK 2 93.232 11.67 93.352 17.82 ;
      RECT MASK 2 94.394 11.67 94.514 17.82 ;
      RECT MASK 2 95.556 11.67 95.676 17.82 ;
      RECT MASK 2 96.42 11.67 96.54 17.85 ;
      RECT MASK 2 97.176 11.67 97.296 14.322 ;
      RECT MASK 2 97.932 11.67 98.052 17.85 ;
      RECT MASK 2 98.688 11.67 98.808 17.82 ;
      RECT MASK 2 99.472 11.67 99.592 17.82 ;
      RECT MASK 2 99.85 11.67 99.97 17.82 ;
      RECT MASK 2 100.228 11.67 100.348 17.82 ;
      RECT MASK 2 101.012 11.67 101.132 17.82 ;
      RECT MASK 2 101.796 11.67 101.916 17.82 ;
      RECT MASK 2 102.174 11.67 102.294 17.82 ;
      RECT MASK 2 102.552 11.67 102.672 17.82 ;
      RECT MASK 2 103.038 11.67 103.158 17.85 ;
      RECT MASK 2 103.416 11.67 103.536 17.85 ;
      RECT MASK 2 103.794 11.67 103.914 17.85 ;
      RECT MASK 2 104.172 11.67 104.292 14.322 ;
      RECT MASK 2 104.55 11.67 104.67 17.85 ;
      RECT MASK 2 104.928 11.67 105.048 17.82 ;
      RECT MASK 2 105.306 11.67 105.426 17.82 ;
      RECT MASK 2 105.684 11.67 105.804 17.82 ;
      RECT MASK 2 106.09 11.67 106.21 17.82 ;
      RECT MASK 2 106.468 11.67 106.588 17.82 ;
      RECT MASK 2 107.63 11.67 107.75 17.82 ;
      RECT MASK 2 108.792 11.67 108.912 17.82 ;
      RECT MASK 2 109.656 11.67 109.776 17.85 ;
      RECT MASK 2 110.412 11.67 110.532 17.85 ;
      RECT MASK 2 111.168 11.67 111.288 17.85 ;
      RECT MASK 2 41.541 12.656 41.601 14.458 ;
      RECT MASK 2 52.775 13.13 52.835 16.672 ;
      RECT MASK 2 81.175 13.136 81.235 16.768 ;
      RECT MASK 2 15.391 14.672 15.451 16.768 ;
      RECT MASK 2 28.627 14.672 28.687 16.768 ;
      RECT MASK 2 41.863 14.672 41.923 16.768 ;
      RECT MASK 2 55.099 14.672 55.159 16.768 ;
      RECT MASK 2 68.741 14.672 68.801 16.768 ;
      RECT MASK 2 67.219 14.768 67.279 16.768 ;
      RECT MASK 2 93.691 14.768 93.751 16.768 ;
      RECT MASK 2 106.807 14.768 106.867 16.768 ;
      RECT MASK 2 53.097 14.864 53.157 16.768 ;
      RECT MASK 2 41.45 15.013 41.57 17.82 ;
      RECT MASK 2 44.191 15.05 44.251 17.434 ;
      RECT MASK 2 80.335 15.05 80.395 17.538 ;
      RECT MASK 2 97.613 15.05 97.673 17.434 ;
      RECT MASK 2 104.129 15.05 104.189 17.434 ;
      RECT MASK 2 67.169 17.23 67.249 18.1345 ;
      RECT MASK 2 60.142 17.52 60.262 84.25 ;
      RECT MASK 2 57.09 18.344 57.21 22.36 ;
      RECT MASK 2 57.846 18.38 57.966 22.36 ;
      RECT MASK 2 6.82 18.45 6.94 85.5325 ;
      RECT MASK 2 7.576 18.45 7.696 85.5325 ;
      RECT MASK 2 7.982 18.45 8.102 85.5325 ;
      RECT MASK 2 8.738 18.45 8.858 85.53 ;
      RECT MASK 2 9.144 18.45 9.264 85.5325 ;
      RECT MASK 2 9.9 18.45 10.02 85.5325 ;
      RECT MASK 2 12.276 18.45 12.396 85.5325 ;
      RECT MASK 2 13.032 18.45 13.152 85.5325 ;
      RECT MASK 2 13.438 18.45 13.558 85.5325 ;
      RECT MASK 2 14.194 18.45 14.314 85.5325 ;
      RECT MASK 2 14.6 18.45 14.72 85.5325 ;
      RECT MASK 2 15.356 18.45 15.476 85.5325 ;
      RECT MASK 2 15.762 18.45 15.882 85.5325 ;
      RECT MASK 2 16.518 18.45 16.638 85.5325 ;
      RECT MASK 2 18.894 18.45 19.014 85.5325 ;
      RECT MASK 2 19.65 18.45 19.77 85.5325 ;
      RECT MASK 2 20.056 18.45 20.176 85.5325 ;
      RECT MASK 2 20.812 18.45 20.932 85.5325 ;
      RECT MASK 2 21.218 18.45 21.338 85.5325 ;
      RECT MASK 2 21.974 18.45 22.094 85.5325 ;
      RECT MASK 2 22.38 18.45 22.5 85.5325 ;
      RECT MASK 2 23.136 18.45 23.256 85.5325 ;
      RECT MASK 2 25.512 18.45 25.632 85.5325 ;
      RECT MASK 2 26.268 18.45 26.388 85.5325 ;
      RECT MASK 2 26.674 18.45 26.794 85.5325 ;
      RECT MASK 2 27.43 18.45 27.55 85.5325 ;
      RECT MASK 2 27.836 18.45 27.956 85.5325 ;
      RECT MASK 2 28.592 18.45 28.712 85.5325 ;
      RECT MASK 2 28.998 18.45 29.118 85.5325 ;
      RECT MASK 2 29.754 18.45 29.874 85.5325 ;
      RECT MASK 2 32.13 18.45 32.25 85.5325 ;
      RECT MASK 2 32.886 18.45 33.006 85.5325 ;
      RECT MASK 2 33.292 18.45 33.412 85.5325 ;
      RECT MASK 2 34.048 18.45 34.168 85.5325 ;
      RECT MASK 2 34.454 18.45 34.574 85.5325 ;
      RECT MASK 2 35.21 18.45 35.33 85.5325 ;
      RECT MASK 2 35.616 18.45 35.736 85.5325 ;
      RECT MASK 2 36.372 18.45 36.492 85.5325 ;
      RECT MASK 2 38.748 18.45 38.868 85.5325 ;
      RECT MASK 2 39.504 18.45 39.624 85.5325 ;
      RECT MASK 2 39.91 18.45 40.03 85.5325 ;
      RECT MASK 2 40.666 18.45 40.786 85.5325 ;
      RECT MASK 2 41.072 18.45 41.192 85.5325 ;
      RECT MASK 2 41.828 18.45 41.948 85.5325 ;
      RECT MASK 2 42.234 18.45 42.354 85.5325 ;
      RECT MASK 2 42.99 18.45 43.11 85.5325 ;
      RECT MASK 2 45.366 18.45 45.486 85.5325 ;
      RECT MASK 2 46.122 18.45 46.242 85.5325 ;
      RECT MASK 2 46.528 18.45 46.648 85.5325 ;
      RECT MASK 2 47.284 18.45 47.404 85.5325 ;
      RECT MASK 2 47.69 18.45 47.81 85.5325 ;
      RECT MASK 2 48.446 18.45 48.566 85.5325 ;
      RECT MASK 2 48.852 18.45 48.972 85.5325 ;
      RECT MASK 2 49.608 18.45 49.728 85.5325 ;
      RECT MASK 2 51.984 18.45 52.104 85.5325 ;
      RECT MASK 2 52.74 18.45 52.86 85.5325 ;
      RECT MASK 2 53.146 18.45 53.266 85.5325 ;
      RECT MASK 2 53.902 18.45 54.022 85.5325 ;
      RECT MASK 2 54.308 18.45 54.428 85.5325 ;
      RECT MASK 2 55.064 18.45 55.184 85.5325 ;
      RECT MASK 2 55.47 18.45 55.59 85.5325 ;
      RECT MASK 2 56.226 18.45 56.346 85.5325 ;
      RECT MASK 2 58.602 18.45 58.722 85.5325 ;
      RECT MASK 2 59.358 18.45 59.478 85.5325 ;
      RECT MASK 2 59.764 18.45 59.884 85.5325 ;
      RECT MASK 2 60.52 18.45 60.64 85.5325 ;
      RECT MASK 2 60.926 18.45 61.046 85.5325 ;
      RECT MASK 2 61.682 18.45 61.802 85.5325 ;
      RECT MASK 2 62.088 18.45 62.208 85.5325 ;
      RECT MASK 2 62.844 18.45 62.964 85.5325 ;
      RECT MASK 2 65.22 18.45 65.34 85.5325 ;
      RECT MASK 2 65.976 18.45 66.096 85.5325 ;
      RECT MASK 2 66.382 18.45 66.502 85.5325 ;
      RECT MASK 2 67.138 18.45 67.258 85.5325 ;
      RECT MASK 2 67.544 18.45 67.664 85.5325 ;
      RECT MASK 2 68.3 18.45 68.42 85.5325 ;
      RECT MASK 2 68.706 18.45 68.826 85.5325 ;
      RECT MASK 2 69.462 18.45 69.582 85.5325 ;
      RECT MASK 2 71.838 18.45 71.958 85.5325 ;
      RECT MASK 2 72.594 18.45 72.714 85.5325 ;
      RECT MASK 2 73 18.45 73.12 85.5325 ;
      RECT MASK 2 73.756 18.45 73.876 85.5325 ;
      RECT MASK 2 74.162 18.45 74.282 85.5325 ;
      RECT MASK 2 74.918 18.45 75.038 85.5325 ;
      RECT MASK 2 75.324 18.45 75.444 85.5325 ;
      RECT MASK 2 76.08 18.45 76.2 85.5325 ;
      RECT MASK 2 78.456 18.45 78.576 85.5325 ;
      RECT MASK 2 79.212 18.45 79.332 85.5325 ;
      RECT MASK 2 79.618 18.45 79.738 85.5325 ;
      RECT MASK 2 80.374 18.45 80.494 85.5325 ;
      RECT MASK 2 80.78 18.45 80.9 85.5325 ;
      RECT MASK 2 81.536 18.45 81.656 85.5325 ;
      RECT MASK 2 81.942 18.45 82.062 85.5325 ;
      RECT MASK 2 82.698 18.45 82.818 85.5325 ;
      RECT MASK 2 85.074 18.45 85.194 85.5325 ;
      RECT MASK 2 85.83 18.45 85.95 85.5325 ;
      RECT MASK 2 86.236 18.45 86.356 85.5325 ;
      RECT MASK 2 86.992 18.45 87.112 85.5325 ;
      RECT MASK 2 87.398 18.45 87.518 85.5325 ;
      RECT MASK 2 88.154 18.45 88.274 85.5325 ;
      RECT MASK 2 88.56 18.45 88.68 85.5325 ;
      RECT MASK 2 89.316 18.45 89.436 85.5325 ;
      RECT MASK 2 91.692 18.45 91.812 85.5325 ;
      RECT MASK 2 92.448 18.45 92.568 85.5325 ;
      RECT MASK 2 92.854 18.45 92.974 85.5325 ;
      RECT MASK 2 93.61 18.45 93.73 85.5325 ;
      RECT MASK 2 94.016 18.45 94.136 85.5325 ;
      RECT MASK 2 94.772 18.45 94.892 85.5325 ;
      RECT MASK 2 95.178 18.45 95.298 85.5325 ;
      RECT MASK 2 95.934 18.45 96.054 85.5325 ;
      RECT MASK 2 98.31 18.45 98.43 85.5325 ;
      RECT MASK 2 99.066 18.45 99.186 85.5325 ;
      RECT MASK 2 99.472 18.45 99.592 85.5325 ;
      RECT MASK 2 100.228 18.45 100.348 85.5325 ;
      RECT MASK 2 100.634 18.45 100.754 85.5325 ;
      RECT MASK 2 101.39 18.45 101.51 85.5325 ;
      RECT MASK 2 101.796 18.45 101.916 85.5325 ;
      RECT MASK 2 102.552 18.45 102.672 85.5325 ;
      RECT MASK 2 104.928 18.45 105.048 85.5325 ;
      RECT MASK 2 105.684 18.45 105.804 85.5325 ;
      RECT MASK 2 106.09 18.45 106.21 85.5325 ;
      RECT MASK 2 106.846 18.45 106.966 85.5325 ;
      RECT MASK 2 107.252 18.45 107.372 85.5325 ;
      RECT MASK 2 108.008 18.45 108.128 85.5325 ;
      RECT MASK 2 108.414 18.45 108.534 85.5325 ;
      RECT MASK 2 109.17 18.45 109.29 85.5325 ;
      RECT MASK 2 12.654 19.535 12.774 84.1645 ;
      RECT MASK 2 13.816 19.535 13.936 84.1645 ;
      RECT MASK 2 14.978 19.535 15.098 84.1645 ;
      RECT MASK 2 16.14 19.535 16.26 84.1645 ;
      RECT MASK 2 19.272 19.535 19.392 84.1645 ;
      RECT MASK 2 20.434 19.535 20.554 84.1645 ;
      RECT MASK 2 21.596 19.535 21.716 84.1645 ;
      RECT MASK 2 22.758 19.535 22.878 84.1645 ;
      RECT MASK 2 25.89 19.535 26.01 84.1645 ;
      RECT MASK 2 27.052 19.535 27.172 84.1645 ;
      RECT MASK 2 28.214 19.535 28.334 84.1645 ;
      RECT MASK 2 29.376 19.535 29.496 84.1645 ;
      RECT MASK 2 32.508 19.535 32.628 84.1645 ;
      RECT MASK 2 33.67 19.535 33.79 84.1645 ;
      RECT MASK 2 34.832 19.535 34.952 84.1645 ;
      RECT MASK 2 35.994 19.535 36.114 84.1645 ;
      RECT MASK 2 39.126 19.535 39.246 84.1645 ;
      RECT MASK 2 40.288 19.535 40.408 84.1645 ;
      RECT MASK 2 41.45 19.535 41.57 84.1645 ;
      RECT MASK 2 42.612 19.535 42.732 84.1645 ;
      RECT MASK 2 45.744 19.535 45.864 84.1645 ;
      RECT MASK 2 46.906 19.535 47.026 84.1645 ;
      RECT MASK 2 48.068 19.535 48.188 84.1645 ;
      RECT MASK 2 49.23 19.535 49.35 84.1645 ;
      RECT MASK 2 52.362 19.535 52.482 84.1645 ;
      RECT MASK 2 53.524 19.535 53.644 84.1645 ;
      RECT MASK 2 54.686 19.535 54.806 84.1645 ;
      RECT MASK 2 55.848 19.535 55.968 84.1645 ;
      RECT MASK 2 65.598 19.535 65.718 84.1645 ;
      RECT MASK 2 66.76 19.535 66.88 84.1645 ;
      RECT MASK 2 67.922 19.535 68.042 84.1645 ;
      RECT MASK 2 69.084 19.535 69.204 84.1645 ;
      RECT MASK 2 72.216 19.535 72.336 84.1645 ;
      RECT MASK 2 73.378 19.535 73.498 84.1645 ;
      RECT MASK 2 74.54 19.535 74.66 84.1645 ;
      RECT MASK 2 75.702 19.535 75.822 84.1645 ;
      RECT MASK 2 78.834 19.535 78.954 84.1645 ;
      RECT MASK 2 79.996 19.535 80.116 84.1645 ;
      RECT MASK 2 81.158 19.535 81.278 84.1645 ;
      RECT MASK 2 82.32 19.535 82.44 84.1645 ;
      RECT MASK 2 85.452 19.535 85.572 84.1645 ;
      RECT MASK 2 86.614 19.535 86.734 84.1645 ;
      RECT MASK 2 87.776 19.535 87.896 84.1645 ;
      RECT MASK 2 88.938 19.535 89.058 84.1645 ;
      RECT MASK 2 92.07 19.535 92.19 84.1645 ;
      RECT MASK 2 93.232 19.535 93.352 84.1645 ;
      RECT MASK 2 94.394 19.535 94.514 84.1645 ;
      RECT MASK 2 95.556 19.535 95.676 84.1645 ;
      RECT MASK 2 98.688 19.535 98.808 84.1645 ;
      RECT MASK 2 99.85 19.535 99.97 84.1645 ;
      RECT MASK 2 101.012 19.535 101.132 84.1645 ;
      RECT MASK 2 102.174 19.535 102.294 84.1645 ;
      RECT MASK 2 105.306 19.535 105.426 84.1645 ;
      RECT MASK 2 106.468 19.535 106.588 84.1645 ;
      RECT MASK 2 107.63 19.535 107.75 84.1645 ;
      RECT MASK 2 108.792 19.535 108.912 84.1645 ;
      RECT MASK 2 2.362 19.63 2.422 24.53 ;
      RECT MASK 2 2.636 19.63 2.696 24.53 ;
      RECT MASK 2 2.91 19.63 2.97 24.53 ;
      RECT MASK 2 3.184 19.63 3.244 24.53 ;
      RECT MASK 2 3.458 19.63 3.518 24.53 ;
      RECT MASK 2 3.732 19.63 3.792 24.53 ;
      RECT MASK 2 5.658 21.27 5.778 26.01 ;
      RECT MASK 2 6.414 21.27 6.534 26.01 ;
      RECT MASK 2 112.592 22.51 112.712 81.47 ;
      RECT MASK 2 111.679 24.144 111.799 79.903 ;
      RECT MASK 2 110.47 26.1 110.59 77.719 ;
      RECT MASK 2 111.226 26.1 111.346 77.719 ;
      RECT MASK 2 113.116 26.1 113.236 77.719 ;
      RECT MASK 2 113.872 26.1 113.992 78.249 ;
      RECT MASK 2 116.701 26.94 116.841 29.48 ;
      RECT MASK 2 117.318 26.94 117.358 28.18 ;
      RECT MASK 2 117.696 26.94 117.736 28.18 ;
      RECT MASK 2 118.074 26.94 118.114 28.18 ;
      RECT MASK 2 118.452 26.94 118.492 28.18 ;
      RECT MASK 2 118.83 26.94 118.87 28.18 ;
      RECT MASK 2 119.208 26.94 119.248 28.18 ;
      RECT MASK 2 119.586 26.94 119.626 28.18 ;
      RECT MASK 2 119.964 26.94 120.004 28.18 ;
      RECT MASK 2 120.342 26.94 120.382 28.18 ;
      RECT MASK 2 120.72 26.94 120.76 28.18 ;
      RECT MASK 2 121.098 26.94 121.138 28.18 ;
      RECT MASK 2 121.476 26.94 121.516 28.18 ;
      RECT MASK 2 121.854 26.94 121.894 28.18 ;
      RECT MASK 2 122.232 26.94 122.272 28.18 ;
      RECT MASK 2 122.61 26.94 122.65 28.18 ;
      RECT MASK 2 122.988 26.94 123.028 28.18 ;
      RECT MASK 2 123.366 26.94 123.406 28.18 ;
      RECT MASK 2 123.744 26.94 123.784 28.18 ;
      RECT MASK 2 124.122 26.94 124.162 28.18 ;
      RECT MASK 2 124.5 26.94 124.54 28.18 ;
      RECT MASK 2 124.878 26.94 124.918 28.18 ;
      RECT MASK 2 125.256 26.94 125.296 28.18 ;
      RECT MASK 2 125.634 26.94 125.674 28.18 ;
      RECT MASK 2 115.006 27.027 115.126 72.532 ;
      RECT MASK 2 117.318 28.7615 117.358 51.3195 ;
      RECT MASK 2 117.696 28.7615 117.736 51.3195 ;
      RECT MASK 2 118.074 28.7615 118.114 51.3195 ;
      RECT MASK 2 118.452 28.7615 118.492 51.3195 ;
      RECT MASK 2 118.83 28.7615 118.87 51.3195 ;
      RECT MASK 2 119.208 28.7615 119.248 51.3195 ;
      RECT MASK 2 119.586 28.7615 119.626 51.3195 ;
      RECT MASK 2 119.964 28.7615 120.004 51.3195 ;
      RECT MASK 2 120.342 28.7615 120.382 51.3195 ;
      RECT MASK 2 120.72 28.7615 120.76 51.3195 ;
      RECT MASK 2 121.098 28.7615 121.138 51.3195 ;
      RECT MASK 2 121.476 28.7615 121.516 51.3195 ;
      RECT MASK 2 121.854 28.7615 121.894 51.3195 ;
      RECT MASK 2 122.232 28.7615 122.272 51.3195 ;
      RECT MASK 2 122.61 28.7615 122.65 51.3195 ;
      RECT MASK 2 122.988 28.7615 123.028 51.3195 ;
      RECT MASK 2 123.366 28.7615 123.406 51.3195 ;
      RECT MASK 2 123.744 28.7615 123.784 51.3195 ;
      RECT MASK 2 124.122 28.7615 124.162 51.3195 ;
      RECT MASK 2 124.5 28.7615 124.54 51.3195 ;
      RECT MASK 2 124.878 28.7615 124.918 51.3195 ;
      RECT MASK 2 125.256 28.7615 125.296 51.3195 ;
      RECT MASK 2 125.634 28.7615 125.674 51.3195 ;
      RECT MASK 2 126.5675 30.141 126.6875 72.484 ;
      RECT MASK 2 128.236 31.175 128.356 72.484 ;
      RECT MASK 2 117.467 51.78 117.587 69.9575 ;
      RECT MASK 2 118.223 51.78 118.343 69.9575 ;
      RECT MASK 2 118.979 51.78 119.099 69.9575 ;
      RECT MASK 2 119.735 51.78 119.855 69.9575 ;
      RECT MASK 2 120.491 51.78 120.611 69.9575 ;
      RECT MASK 2 121.247 51.78 121.367 69.9575 ;
      RECT MASK 2 122.003 51.78 122.123 69.9575 ;
      RECT MASK 2 122.759 51.78 122.879 69.9575 ;
      RECT MASK 2 123.515 51.78 123.635 69.9575 ;
      RECT MASK 2 124.271 51.78 124.391 69.9575 ;
      RECT MASK 2 125.027 51.78 125.147 69.9575 ;
      RECT MASK 2 125.783 51.78 125.903 69.9575 ;
      RECT MASK 2 117.079 52.687 117.219 76.57 ;
      RECT MASK 2 117.835 52.687 117.975 76.57 ;
      RECT MASK 2 118.591 52.687 118.731 76.57 ;
      RECT MASK 2 119.347 52.687 119.487 76.57 ;
      RECT MASK 2 120.103 52.687 120.243 76.57 ;
      RECT MASK 2 120.859 52.687 120.999 76.57 ;
      RECT MASK 2 121.615 52.687 121.755 76.57 ;
      RECT MASK 2 122.371 52.687 122.511 76.57 ;
      RECT MASK 2 123.127 52.687 123.267 76.57 ;
      RECT MASK 2 123.883 52.687 124.023 76.57 ;
      RECT MASK 2 124.639 52.687 124.779 76.57 ;
      RECT MASK 2 125.395 52.687 125.535 76.57 ;
      RECT MASK 2 116.701 70.8925 116.841 79.4 ;
      RECT MASK 2 117.457 70.8925 117.597 79.4 ;
      RECT MASK 2 118.213 70.8925 118.353 79.4 ;
      RECT MASK 2 118.969 70.8925 119.109 79.4 ;
      RECT MASK 2 119.725 70.8925 119.865 79.4 ;
      RECT MASK 2 120.481 70.8925 120.621 79.4 ;
      RECT MASK 2 121.237 70.8925 121.377 79.4 ;
      RECT MASK 2 121.993 70.8925 122.133 79.4 ;
      RECT MASK 2 122.749 70.8925 122.889 79.4 ;
      RECT MASK 2 123.505 70.8925 123.645 79.4 ;
      RECT MASK 2 124.261 70.8925 124.401 79.4 ;
      RECT MASK 2 125.017 70.8925 125.157 79.4 ;
      RECT MASK 2 125.773 70.8925 125.913 79.4 ;
      RECT MASK 2 117.079 77.12 117.219 80.393 ;
      RECT MASK 2 117.835 77.12 117.975 80.393 ;
      RECT MASK 2 118.591 77.12 118.731 80.393 ;
      RECT MASK 2 119.347 77.12 119.487 80.393 ;
      RECT MASK 2 120.103 77.12 120.243 80.393 ;
      RECT MASK 2 120.859 77.12 120.999 80.393 ;
      RECT MASK 2 121.615 77.12 121.755 80.393 ;
      RECT MASK 2 122.371 77.12 122.511 80.393 ;
      RECT MASK 2 123.127 77.12 123.267 80.393 ;
      RECT MASK 2 123.883 77.12 124.023 80.393 ;
      RECT MASK 2 124.639 77.12 124.779 80.393 ;
      RECT MASK 2 125.395 77.12 125.535 80.393 ;
      RECT MASK 2 112.095 77.613 112.215 85.549 ;
      RECT MASK 2 113.229 78.04 113.349 85.549 ;
      RECT MASK 2 2.204 79.12 2.264 95.78 ;
      RECT MASK 2 2.478 79.12 2.538 95.78 ;
      RECT MASK 2 2.752 79.12 2.812 95.78 ;
      RECT MASK 2 3.026 79.12 3.086 95.78 ;
      RECT MASK 2 3.3 79.12 3.36 95.78 ;
      RECT MASK 2 3.574 79.12 3.634 95.78 ;
      RECT MASK 2 3.848 79.12 3.908 95.78 ;
      RECT MASK 2 4.122 79.12 4.182 95.78 ;
      RECT MASK 2 4.396 79.12 4.456 95.78 ;
      RECT MASK 2 57.498 80.465 57.578 84.25 ;
      RECT MASK 2 57.876 80.465 57.956 84.25 ;
      RECT MASK 2 58.254 80.465 58.334 84.25 ;
      RECT MASK 2 63.106 80.465 63.186 84.25 ;
      RECT MASK 2 63.484 80.465 63.564 84.25 ;
      RECT MASK 2 63.862 80.465 63.942 84.25 ;
      RECT MASK 2 111.466 80.65 111.586 84.174 ;
      RECT MASK 2 116.599 81.814 116.659 96.653 ;
      RECT MASK 2 116.873 81.814 116.933 96.653 ;
      RECT MASK 2 117.147 81.814 117.207 96.653 ;
      RECT MASK 2 117.421 81.814 117.481 96.653 ;
      RECT MASK 2 117.695 81.814 117.755 96.653 ;
      RECT MASK 2 117.969 81.814 118.029 96.653 ;
      RECT MASK 2 118.243 81.814 118.303 96.653 ;
      RECT MASK 2 118.517 81.814 118.577 96.653 ;
      RECT MASK 2 118.791 81.814 118.851 96.653 ;
      RECT MASK 2 119.065 81.814 119.125 96.653 ;
      RECT MASK 2 119.339 81.814 119.399 96.653 ;
      RECT MASK 2 119.613 81.814 119.673 96.653 ;
      RECT MASK 2 119.887 81.814 119.947 96.653 ;
      RECT MASK 2 120.161 81.814 120.221 96.653 ;
      RECT MASK 2 120.435 81.814 120.495 96.653 ;
      RECT MASK 2 120.709 81.814 120.769 96.653 ;
      RECT MASK 2 120.983 81.814 121.043 96.653 ;
      RECT MASK 2 121.257 81.814 121.317 96.653 ;
      RECT MASK 2 121.531 81.814 121.591 96.653 ;
      RECT MASK 2 121.805 81.814 121.865 96.653 ;
      RECT MASK 2 122.079 81.814 122.139 96.653 ;
      RECT MASK 2 122.353 81.814 122.413 96.653 ;
      RECT MASK 2 122.627 81.814 122.687 96.653 ;
      RECT MASK 2 122.901 81.814 122.961 96.653 ;
      RECT MASK 2 123.175 81.814 123.235 96.653 ;
      RECT MASK 2 123.449 81.814 123.509 96.653 ;
      RECT MASK 2 123.723 81.814 123.783 96.653 ;
      RECT MASK 2 123.997 81.814 124.057 96.653 ;
      RECT MASK 2 124.271 81.814 124.331 96.653 ;
      RECT MASK 2 124.545 81.814 124.605 96.653 ;
      RECT MASK 2 124.819 81.814 124.879 96.653 ;
      RECT MASK 2 125.093 81.814 125.153 96.653 ;
      RECT MASK 2 125.367 81.814 125.427 96.653 ;
      RECT MASK 2 125.641 81.814 125.701 96.653 ;
      RECT MASK 2 125.915 81.814 125.975 96.653 ;
      RECT MASK 2 126.189 81.814 126.249 96.653 ;
      RECT MASK 2 126.463 81.814 126.523 96.653 ;
      RECT MASK 2 126.737 81.814 126.797 96.653 ;
      RECT MASK 2 127.011 81.814 127.071 96.653 ;
      RECT MASK 2 127.285 81.814 127.345 96.653 ;
      RECT MASK 2 127.559 81.814 127.619 96.653 ;
      RECT MASK 2 24.397 85.686 24.497 94.49 ;
      RECT MASK 2 18.2105 86.43 18.3105 93.48 ;
      RECT MASK 2 21.5305 86.43 21.6305 93.48 ;
      RECT MASK 2 36.328 86.996 36.778 94.67 ;
      RECT MASK 2 66.024 86.996 66.474 94.67 ;
      RECT MASK 2 72.718 86.996 73.168 94.67 ;
      RECT MASK 2 102.414 86.996 102.864 94.67 ;
      RECT MASK 2 37.048 87.021 65.754 87.081 ;
      RECT MASK 2 73.438 87.021 102.144 87.081 ;
      RECT MASK 2 14.7495 87.06 14.8295 89.2865 ;
      RECT MASK 2 15.0815 87.06 15.1615 89.2865 ;
      RECT MASK 2 15.4135 87.06 15.4935 89.2865 ;
      RECT MASK 2 25.68 87.101 25.74 88.982 ;
      RECT MASK 2 26.048 87.101 26.108 88.982 ;
      RECT MASK 2 26.36 87.101 26.42 88.982 ;
      RECT MASK 2 26.63 87.101 26.69 88.982 ;
      RECT MASK 2 26.9 87.101 26.96 88.982 ;
      RECT MASK 2 27.17 87.101 27.23 88.982 ;
      RECT MASK 2 27.44 87.101 27.5 88.982 ;
      RECT MASK 2 27.71 87.101 27.77 88.982 ;
      RECT MASK 2 27.98 87.101 28.04 88.982 ;
      RECT MASK 2 28.25 87.101 28.31 88.982 ;
      RECT MASK 2 28.52 87.101 28.58 88.982 ;
      RECT MASK 2 28.79 87.101 28.85 88.982 ;
      RECT MASK 2 29.06 87.101 29.12 88.982 ;
      RECT MASK 2 29.33 87.101 29.39 88.982 ;
      RECT MASK 2 29.6 87.101 29.66 88.982 ;
      RECT MASK 2 29.87 87.101 29.93 88.982 ;
      RECT MASK 2 30.182 87.101 30.242 88.982 ;
      RECT MASK 2 30.55 87.101 30.61 88.982 ;
      RECT MASK 2 6.309 87.244 6.409 94.316 ;
      RECT MASK 2 7.2325 87.244 7.3325 94.316 ;
      RECT MASK 2 37.048 87.273 65.754 87.333 ;
      RECT MASK 2 73.438 87.273 102.144 87.333 ;
      RECT MASK 2 22.758 87.285 22.878 96.81 ;
      RECT MASK 2 23.136 87.285 23.256 96.81 ;
      RECT MASK 2 67.5 87.416 71.692 87.516 ;
      RECT MASK 2 103.89 87.416 106.869 87.516 ;
      RECT MASK 2 32.279 87.431 35.302 87.531 ;
      RECT MASK 2 9.8675 87.52 9.9475 89.2865 ;
      RECT MASK 2 10.1995 87.52 10.2795 89.2865 ;
      RECT MASK 2 10.5315 87.52 10.6115 89.2865 ;
      RECT MASK 2 10.8635 87.52 10.9435 89.2865 ;
      RECT MASK 2 11.1955 87.52 11.2755 89.2865 ;
      RECT MASK 2 19.2995 87.52 19.3795 89.2865 ;
      RECT MASK 2 19.6315 87.52 19.7115 89.2865 ;
      RECT MASK 2 19.9635 87.52 20.0435 89.2865 ;
      RECT MASK 2 20.2955 87.52 20.3755 89.2865 ;
      RECT MASK 2 20.6275 87.52 20.7075 89.2865 ;
      RECT MASK 2 107.557 87.72 107.617 96.653 ;
      RECT MASK 2 107.831 87.72 107.891 96.653 ;
      RECT MASK 2 108.105 87.72 108.165 96.653 ;
      RECT MASK 2 108.379 87.72 108.439 96.653 ;
      RECT MASK 2 108.653 87.72 108.713 96.653 ;
      RECT MASK 2 108.927 87.72 108.987 96.653 ;
      RECT MASK 2 109.201 87.72 109.261 96.653 ;
      RECT MASK 2 109.475 87.72 109.535 96.653 ;
      RECT MASK 2 109.749 87.72 109.809 96.653 ;
      RECT MASK 2 110.023 87.72 110.083 96.653 ;
      RECT MASK 2 110.297 87.72 110.357 96.653 ;
      RECT MASK 2 110.571 87.72 110.631 96.653 ;
      RECT MASK 2 110.845 87.72 110.905 96.653 ;
      RECT MASK 2 111.119 87.72 111.179 96.653 ;
      RECT MASK 2 111.393 87.72 111.453 96.653 ;
      RECT MASK 2 111.667 87.72 111.727 96.653 ;
      RECT MASK 2 111.941 87.72 112.001 96.653 ;
      RECT MASK 2 112.215 87.72 112.275 96.653 ;
      RECT MASK 2 112.489 87.72 112.549 96.653 ;
      RECT MASK 2 112.763 87.72 112.823 96.653 ;
      RECT MASK 2 113.037 87.72 113.097 96.653 ;
      RECT MASK 2 113.311 87.72 113.371 96.653 ;
      RECT MASK 2 113.585 87.72 113.645 96.653 ;
      RECT MASK 2 113.859 87.72 113.919 96.653 ;
      RECT MASK 2 114.133 87.72 114.193 96.653 ;
      RECT MASK 2 114.407 87.72 114.467 96.653 ;
      RECT MASK 2 114.681 87.72 114.741 96.653 ;
      RECT MASK 2 114.955 87.72 115.015 96.653 ;
      RECT MASK 2 115.229 87.72 115.289 96.653 ;
      RECT MASK 2 115.503 87.72 115.563 96.653 ;
      RECT MASK 2 115.777 87.72 115.837 96.653 ;
      RECT MASK 2 116.051 87.72 116.111 96.653 ;
      RECT MASK 2 116.325 87.72 116.385 96.653 ;
      RECT MASK 2 67.5 87.768 71.692 87.868 ;
      RECT MASK 2 103.89 87.768 106.869 87.868 ;
      RECT MASK 2 32.279 87.783 35.302 87.883 ;
      RECT MASK 2 23.514 87.87 23.634 96.81 ;
      RECT MASK 2 23.892 87.87 24.012 96.81 ;
      RECT MASK 2 37.048 87.921 65.754 87.981 ;
      RECT MASK 2 73.438 87.921 102.144 87.981 ;
      RECT MASK 2 8.409 88.08 8.529 89.7135 ;
      RECT MASK 2 8.8115 88.08 8.9315 89.7135 ;
      RECT MASK 2 9.2115 88.08 9.3315 88.7365 ;
      RECT MASK 2 11.6115 88.08 11.7315 88.7365 ;
      RECT MASK 2 12.0635 88.08 12.1835 89.7135 ;
      RECT MASK 2 12.466 88.08 12.586 89.7135 ;
      RECT MASK 2 12.953 88.08 13.073 89.7135 ;
      RECT MASK 2 13.517 88.08 13.637 89.7135 ;
      RECT MASK 2 14.0115 88.08 14.1315 88.7365 ;
      RECT MASK 2 14.4115 88.08 14.5315 88.7365 ;
      RECT MASK 2 15.8115 88.08 15.9315 88.7365 ;
      RECT MASK 2 16.2115 88.08 16.3315 88.7365 ;
      RECT MASK 2 67.5 88.12 71.692 88.22 ;
      RECT MASK 2 103.89 88.12 106.869 88.22 ;
      RECT MASK 2 32.279 88.135 35.302 88.235 ;
      RECT MASK 2 37.048 88.173 65.754 88.233 ;
      RECT MASK 2 73.438 88.173 102.144 88.233 ;
      RECT MASK 2 9.5355 88.412 9.6155 89.8155 ;
      RECT MASK 2 18.9675 88.412 19.0475 89.8155 ;
      RECT MASK 2 67.5 88.472 71.692 88.572 ;
      RECT MASK 2 103.89 88.472 106.869 88.572 ;
      RECT MASK 2 32.279 88.487 35.302 88.587 ;
      RECT MASK 2 37.048 88.821 65.754 88.881 ;
      RECT MASK 2 73.438 88.821 102.144 88.881 ;
      RECT MASK 2 67.5 88.824 71.692 88.924 ;
      RECT MASK 2 103.89 88.824 106.869 88.924 ;
      RECT MASK 2 32.279 88.839 35.302 88.939 ;
      RECT MASK 2 9.2035 89.025 9.2835 92.535 ;
      RECT MASK 2 11.5275 89.025 11.6075 92.535 ;
      RECT MASK 2 11.8595 89.025 11.9395 92.535 ;
      RECT MASK 2 14.0855 89.025 14.1655 90.39 ;
      RECT MASK 2 14.4175 89.025 14.4975 90.39 ;
      RECT MASK 2 16.0775 89.025 16.1575 90.39 ;
      RECT MASK 2 18.6355 89.025 18.7155 92.535 ;
      RECT MASK 2 20.9595 89.025 21.0395 92.535 ;
      RECT MASK 2 21.2915 89.025 21.3715 92.535 ;
      RECT MASK 2 37.048 89.073 65.754 89.133 ;
      RECT MASK 2 73.438 89.073 102.144 89.133 ;
      RECT MASK 2 67.5 89.176 71.692 89.276 ;
      RECT MASK 2 103.89 89.176 106.869 89.276 ;
      RECT MASK 2 32.279 89.191 35.302 89.291 ;
      RECT MASK 2 25.68 89.441 25.74 91.322 ;
      RECT MASK 2 26.048 89.441 26.108 91.322 ;
      RECT MASK 2 26.36 89.441 26.42 91.322 ;
      RECT MASK 2 26.63 89.441 26.69 91.322 ;
      RECT MASK 2 26.9 89.441 26.96 91.322 ;
      RECT MASK 2 27.17 89.441 27.23 91.844 ;
      RECT MASK 2 27.44 89.441 27.5 91.844 ;
      RECT MASK 2 27.71 89.441 27.77 91.844 ;
      RECT MASK 2 27.98 89.441 28.04 91.844 ;
      RECT MASK 2 28.25 89.441 28.31 91.844 ;
      RECT MASK 2 28.52 89.441 28.58 91.844 ;
      RECT MASK 2 28.79 89.441 28.85 91.844 ;
      RECT MASK 2 29.06 89.441 29.12 91.844 ;
      RECT MASK 2 29.33 89.441 29.39 91.844 ;
      RECT MASK 2 29.6 89.441 29.66 91.844 ;
      RECT MASK 2 29.87 89.441 29.93 91.844 ;
      RECT MASK 2 30.182 89.441 30.242 91.322 ;
      RECT MASK 2 30.55 89.441 30.61 91.322 ;
      RECT MASK 2 67.5 89.528 71.692 89.628 ;
      RECT MASK 2 103.89 89.528 106.869 89.628 ;
      RECT MASK 2 32.279 89.543 35.302 89.643 ;
      RECT MASK 2 37.048 89.721 65.754 89.781 ;
      RECT MASK 2 73.438 89.721 102.144 89.781 ;
      RECT MASK 2 10.0325 89.8275 10.1125 91.7075 ;
      RECT MASK 2 10.3655 89.8275 10.4455 91.7075 ;
      RECT MASK 2 10.6995 89.8275 10.7795 91.7075 ;
      RECT MASK 2 11.0325 89.8275 11.1125 91.7075 ;
      RECT MASK 2 14.744 89.8275 14.824 91.913 ;
      RECT MASK 2 15.077 89.8275 15.157 91.913 ;
      RECT MASK 2 15.411 89.8275 15.491 91.913 ;
      RECT MASK 2 15.743 89.8275 15.823 91.913 ;
      RECT MASK 2 19.4665 89.8275 19.5465 91.665 ;
      RECT MASK 2 19.7995 89.8275 19.8795 91.665 ;
      RECT MASK 2 20.1335 89.8275 20.2135 91.665 ;
      RECT MASK 2 20.4665 89.8275 20.5465 91.665 ;
      RECT MASK 2 67.5 89.88 71.692 89.98 ;
      RECT MASK 2 103.89 89.88 106.869 89.98 ;
      RECT MASK 2 32.279 89.895 35.302 89.995 ;
      RECT MASK 2 37.048 89.973 65.754 90.033 ;
      RECT MASK 2 73.438 89.973 102.144 90.033 ;
      RECT MASK 2 13.6575 90.0145 13.7375 94.3995 ;
      RECT MASK 2 16.6715 90.03 16.7515 94.3995 ;
      RECT MASK 2 67.5 90.232 71.692 90.332 ;
      RECT MASK 2 103.89 90.232 106.869 90.332 ;
      RECT MASK 2 32.279 90.247 35.302 90.347 ;
      RECT MASK 2 67.5 90.584 71.692 90.684 ;
      RECT MASK 2 103.89 90.584 106.869 90.684 ;
      RECT MASK 2 32.279 90.599 35.302 90.699 ;
      RECT MASK 2 37.048 90.621 65.754 90.681 ;
      RECT MASK 2 73.438 90.621 102.144 90.681 ;
      RECT MASK 2 37.048 90.873 65.754 90.933 ;
      RECT MASK 2 73.438 90.873 102.144 90.933 ;
      RECT MASK 2 67.5 90.936 71.692 91.036 ;
      RECT MASK 2 103.89 90.936 106.869 91.036 ;
      RECT MASK 2 32.279 90.951 35.302 91.051 ;
      RECT MASK 2 14.0855 91.17 14.1655 92.535 ;
      RECT MASK 2 14.4175 91.17 14.4975 92.535 ;
      RECT MASK 2 16.0775 91.17 16.1575 92.535 ;
      RECT MASK 2 67.5 91.288 71.692 91.388 ;
      RECT MASK 2 103.89 91.288 106.869 91.388 ;
      RECT MASK 2 32.279 91.303 35.302 91.403 ;
      RECT MASK 2 26.36 91.4615 26.42 92.054 ;
      RECT MASK 2 26.63 91.4615 26.69 92.054 ;
      RECT MASK 2 26.9 91.4615 26.96 92.054 ;
      RECT MASK 2 37.048 91.521 65.754 91.581 ;
      RECT MASK 2 73.438 91.521 102.144 91.581 ;
      RECT MASK 2 67.5 91.64 71.692 91.74 ;
      RECT MASK 2 103.89 91.64 106.869 91.74 ;
      RECT MASK 2 32.279 91.655 35.302 91.755 ;
      RECT MASK 2 9.5355 91.7445 9.6155 93.148 ;
      RECT MASK 2 18.9675 91.7445 19.0475 93.148 ;
      RECT MASK 2 37.048 91.773 65.754 91.833 ;
      RECT MASK 2 73.438 91.773 102.144 91.833 ;
      RECT MASK 2 67.5 91.992 71.692 92.092 ;
      RECT MASK 2 103.89 91.992 106.869 92.092 ;
      RECT MASK 2 32.279 92.007 35.302 92.107 ;
      RECT MASK 2 9.8675 92.2735 9.9475 94.04 ;
      RECT MASK 2 10.1995 92.2735 10.2795 94.04 ;
      RECT MASK 2 10.5315 92.2735 10.6115 94.04 ;
      RECT MASK 2 10.8635 92.2735 10.9435 94.04 ;
      RECT MASK 2 14.7495 92.2735 14.8295 94.5 ;
      RECT MASK 2 15.0815 92.2735 15.1615 94.5 ;
      RECT MASK 2 15.4135 92.2735 15.4935 94.5 ;
      RECT MASK 2 19.2995 92.2735 19.3795 94.04 ;
      RECT MASK 2 19.6315 92.2735 19.7115 94.04 ;
      RECT MASK 2 19.9635 92.2735 20.0435 94.04 ;
      RECT MASK 2 20.2955 92.2735 20.3755 94.04 ;
      RECT MASK 2 20.6275 92.2735 20.7075 94.04 ;
      RECT MASK 2 67.5 92.344 71.692 92.444 ;
      RECT MASK 2 103.89 92.344 106.869 92.444 ;
      RECT MASK 2 32.279 92.359 35.302 92.459 ;
      RECT MASK 2 37.048 92.421 65.754 92.481 ;
      RECT MASK 2 73.438 92.421 102.144 92.481 ;
      RECT MASK 2 37.048 92.673 65.754 92.733 ;
      RECT MASK 2 73.438 92.673 102.144 92.733 ;
      RECT MASK 2 67.5 92.696 71.692 92.796 ;
      RECT MASK 2 103.89 92.696 106.869 92.796 ;
      RECT MASK 2 32.279 92.711 35.302 92.811 ;
      RECT MASK 2 8.8675 92.736 8.9675 93.196 ;
      RECT MASK 2 14.0845 92.7795 14.1645 94.3995 ;
      RECT MASK 2 14.4175 92.7795 14.4975 94.3995 ;
      RECT MASK 2 15.7455 92.7795 15.8255 94.3995 ;
      RECT MASK 2 16.0785 92.7795 16.1585 94.3995 ;
      RECT MASK 2 67.5 93.048 71.692 93.148 ;
      RECT MASK 2 103.89 93.048 106.869 93.148 ;
      RECT MASK 2 32.279 93.063 35.302 93.163 ;
      RECT MASK 2 37.048 93.321 65.754 93.381 ;
      RECT MASK 2 73.438 93.321 102.144 93.381 ;
      RECT MASK 2 67.5 93.4 71.692 93.5 ;
      RECT MASK 2 103.89 93.4 106.869 93.5 ;
      RECT MASK 2 32.279 93.415 35.302 93.515 ;
      RECT MASK 2 37.048 93.573 65.754 93.633 ;
      RECT MASK 2 73.438 93.573 102.144 93.633 ;
      RECT MASK 2 25.237 93.748 31.053 94.134 ;
      RECT MASK 2 67.5 93.752 71.692 93.852 ;
      RECT MASK 2 103.89 93.752 106.869 93.852 ;
      RECT MASK 2 32.279 93.767 35.302 93.867 ;
      RECT MASK 2 67.5 94.104 71.692 94.204 ;
      RECT MASK 2 103.89 94.104 106.869 94.204 ;
      RECT MASK 2 32.279 94.119 35.302 94.219 ;
      RECT MASK 2 37.048 94.221 65.754 94.281 ;
      RECT MASK 2 73.438 94.221 102.144 94.281 ;
      RECT MASK 2 37.048 94.473 65.754 94.533 ;
      RECT MASK 2 73.438 94.473 102.144 94.533 ;
      RECT MASK 2 25.026 94.59 25.146 96.81 ;
      RECT MASK 2 25.404 94.59 25.524 96.81 ;
      RECT MASK 2 25.782 94.59 25.902 96.81 ;
      RECT MASK 2 26.16 94.59 26.28 96.81 ;
      RECT MASK 2 26.538 94.59 26.658 96.81 ;
      RECT MASK 2 26.916 94.59 27.036 96.81 ;
      RECT MASK 2 27.294 94.59 27.414 96.81 ;
      RECT MASK 2 27.672 94.59 27.792 96.81 ;
      RECT MASK 2 28.05 94.59 28.17 96.81 ;
      RECT MASK 2 28.428 94.59 28.548 96.81 ;
      RECT MASK 2 28.806 94.59 28.926 96.81 ;
      RECT MASK 2 29.184 94.59 29.304 96.81 ;
      RECT MASK 2 29.562 94.59 29.682 96.81 ;
      RECT MASK 2 29.94 94.59 30.06 96.81 ;
      RECT MASK 2 30.318 94.59 30.438 96.81 ;
      RECT MASK 2 30.696 94.59 30.816 96.81 ;
      RECT MASK 2 31.074 94.59 31.194 96.81 ;
      RECT MASK 2 24.27 95.01 24.39 96.81 ;
      RECT MASK 2 24.648 95.01 24.768 96.81 ;
      RECT MASK 2 31.452 95.85 31.572 96.81 ;
      RECT MASK 2 31.83 95.85 31.95 96.81 ;
      RECT MASK 2 32.208 95.85 32.328 96.81 ;
      RECT MASK 2 32.586 95.85 32.706 96.81 ;
      RECT MASK 2 32.964 95.85 33.084 96.81 ;
      RECT MASK 2 33.342 95.85 33.462 96.81 ;
      RECT MASK 2 33.72 95.85 33.84 96.81 ;
      RECT MASK 2 34.098 95.85 34.218 96.81 ;
      RECT MASK 2 34.476 95.85 34.596 96.81 ;
      RECT MASK 2 34.854 95.85 34.974 96.81 ;
      RECT MASK 2 35.232 95.85 35.352 96.81 ;
      RECT MASK 2 35.61 95.85 35.73 96.81 ;
      RECT MASK 2 35.988 95.85 36.108 96.81 ;
      RECT MASK 2 36.366 95.85 36.486 96.81 ;
      RECT MASK 2 2.338 97.41 2.398 108.838 ;
      RECT MASK 2 2.612 97.41 2.672 108.838 ;
      RECT MASK 2 2.886 97.41 2.946 108.838 ;
      RECT MASK 2 3.16 97.41 3.22 108.838 ;
      RECT MASK 2 3.434 97.41 3.494 108.838 ;
      RECT MASK 2 3.708 97.41 3.768 108.838 ;
      RECT MASK 2 3.982 97.41 4.042 108.838 ;
      RECT MASK 2 4.256 97.41 4.316 108.838 ;
      RECT MASK 2 4.53 97.41 4.59 108.838 ;
      RECT MASK 2 4.804 97.41 4.864 108.838 ;
      RECT MASK 2 5.078 97.41 5.138 108.838 ;
      RECT MASK 2 5.352 97.41 5.412 108.838 ;
      RECT MASK 2 5.626 97.41 5.686 108.838 ;
      RECT MASK 2 5.9 97.41 5.96 108.838 ;
      RECT MASK 2 6.174 97.41 6.234 108.838 ;
      RECT MASK 2 6.448 97.41 6.508 108.838 ;
      RECT MASK 2 6.722 97.41 6.782 108.838 ;
      RECT MASK 2 6.996 97.41 7.056 108.838 ;
      RECT MASK 2 7.27 97.41 7.33 108.838 ;
      RECT MASK 2 7.544 97.41 7.604 108.838 ;
      RECT MASK 2 7.818 97.41 7.878 108.838 ;
      RECT MASK 2 8.092 97.41 8.152 108.838 ;
      RECT MASK 2 8.366 97.41 8.426 108.838 ;
      RECT MASK 2 8.64 97.41 8.7 108.838 ;
      RECT MASK 2 8.914 97.41 8.974 108.838 ;
      RECT MASK 2 9.188 97.41 9.248 108.838 ;
      RECT MASK 2 9.462 97.41 9.522 108.838 ;
      RECT MASK 2 9.736 97.41 9.796 108.838 ;
      RECT MASK 2 10.01 97.41 10.07 108.838 ;
      RECT MASK 2 10.284 97.41 10.344 108.838 ;
      RECT MASK 2 10.558 97.41 10.618 108.838 ;
      RECT MASK 2 10.832 97.41 10.892 108.838 ;
      RECT MASK 2 11.106 97.41 11.166 108.838 ;
      RECT MASK 2 11.38 97.41 11.44 108.838 ;
      RECT MASK 2 11.654 97.41 11.714 108.838 ;
      RECT MASK 2 11.928 97.41 11.988 108.838 ;
      RECT MASK 2 12.202 97.41 12.262 108.838 ;
      RECT MASK 2 12.476 97.41 12.536 108.838 ;
      RECT MASK 2 12.75 97.41 12.81 108.838 ;
      RECT MASK 2 13.024 97.41 13.084 108.838 ;
      RECT MASK 2 13.298 97.41 13.358 108.838 ;
      RECT MASK 2 13.572 97.41 13.632 108.838 ;
      RECT MASK 2 13.846 97.41 13.906 108.838 ;
      RECT MASK 2 14.12 97.41 14.18 108.838 ;
      RECT MASK 2 14.394 97.41 14.454 108.838 ;
      RECT MASK 2 14.668 97.41 14.728 108.838 ;
      RECT MASK 2 14.942 97.41 15.002 108.838 ;
      RECT MASK 2 15.216 97.41 15.276 108.838 ;
      RECT MASK 2 15.49 97.41 15.55 108.838 ;
      RECT MASK 2 15.764 97.41 15.824 108.838 ;
      RECT MASK 2 16.038 97.41 16.098 108.838 ;
      RECT MASK 2 16.312 97.41 16.372 108.838 ;
      RECT MASK 2 16.586 97.41 16.646 108.838 ;
      RECT MASK 2 16.86 97.41 16.92 108.838 ;
      RECT MASK 2 17.134 97.41 17.194 108.838 ;
      RECT MASK 2 17.408 97.41 17.468 108.838 ;
      RECT MASK 2 17.682 97.41 17.742 108.838 ;
      RECT MASK 2 17.956 97.41 18.016 108.838 ;
      RECT MASK 2 18.23 97.41 18.29 108.838 ;
      RECT MASK 2 18.504 97.41 18.564 108.838 ;
      RECT MASK 2 18.778 97.41 18.838 108.838 ;
      RECT MASK 2 19.052 97.41 19.112 108.838 ;
      RECT MASK 2 19.326 97.41 19.386 108.838 ;
      RECT MASK 2 19.6 97.41 19.66 108.838 ;
      RECT MASK 2 19.874 97.41 19.934 108.838 ;
      RECT MASK 2 20.148 97.41 20.208 108.838 ;
      RECT MASK 2 20.422 97.41 20.482 108.838 ;
      RECT MASK 2 20.696 97.41 20.756 108.838 ;
      RECT MASK 2 20.97 97.41 21.03 108.838 ;
      RECT MASK 2 21.244 97.41 21.304 108.838 ;
      RECT MASK 2 21.518 97.41 21.578 108.838 ;
      RECT MASK 2 21.792 97.41 21.852 108.838 ;
      RECT MASK 2 22.066 97.41 22.126 108.838 ;
      RECT MASK 2 22.34 97.41 22.4 108.838 ;
      RECT MASK 2 22.614 97.41 22.674 108.838 ;
      RECT MASK 2 22.888 97.41 22.948 108.838 ;
      RECT MASK 2 23.162 97.41 23.222 108.838 ;
      RECT MASK 2 23.436 97.41 23.496 108.838 ;
      RECT MASK 2 23.71 97.41 23.77 108.838 ;
      RECT MASK 2 23.984 97.41 24.044 108.838 ;
      RECT MASK 2 24.258 97.41 24.318 108.838 ;
      RECT MASK 2 24.532 97.41 24.592 108.838 ;
      RECT MASK 2 24.806 97.41 24.866 108.838 ;
      RECT MASK 2 25.08 97.41 25.14 108.838 ;
      RECT MASK 2 25.354 97.41 25.414 108.838 ;
      RECT MASK 2 25.628 97.41 25.688 108.838 ;
      RECT MASK 2 25.902 97.41 25.962 108.838 ;
      RECT MASK 2 26.176 97.41 26.236 108.838 ;
      RECT MASK 2 26.45 97.41 26.51 108.838 ;
      RECT MASK 2 26.724 97.41 26.784 108.838 ;
      RECT MASK 2 26.998 97.41 27.058 108.838 ;
      RECT MASK 2 27.272 97.41 27.332 108.838 ;
      RECT MASK 2 27.546 97.41 27.606 108.838 ;
      RECT MASK 2 27.82 97.41 27.88 108.838 ;
      RECT MASK 2 28.094 97.41 28.154 108.838 ;
      RECT MASK 2 28.368 97.41 28.428 108.838 ;
      RECT MASK 2 28.642 97.41 28.702 108.838 ;
      RECT MASK 2 28.916 97.41 28.976 108.838 ;
      RECT MASK 2 29.19 97.41 29.25 108.838 ;
      RECT MASK 2 29.464 97.41 29.524 108.838 ;
      RECT MASK 2 29.738 97.41 29.798 108.838 ;
      RECT MASK 2 30.012 97.41 30.072 108.838 ;
      RECT MASK 2 30.286 97.41 30.346 108.838 ;
      RECT MASK 2 30.56 97.41 30.62 108.838 ;
      RECT MASK 2 30.834 97.41 30.894 108.838 ;
      RECT MASK 2 31.108 97.41 31.168 108.838 ;
      RECT MASK 2 31.382 97.41 31.442 108.838 ;
      RECT MASK 2 31.656 97.41 31.716 108.838 ;
      RECT MASK 2 31.93 97.41 31.99 108.838 ;
      RECT MASK 2 32.204 97.41 32.264 108.838 ;
      RECT MASK 2 32.478 97.41 32.538 108.838 ;
      RECT MASK 2 32.752 97.41 32.812 108.838 ;
      RECT MASK 2 33.026 97.41 33.086 108.838 ;
      RECT MASK 2 33.3 97.41 33.36 108.838 ;
      RECT MASK 2 33.574 97.41 33.634 108.838 ;
      RECT MASK 2 33.848 97.41 33.908 108.838 ;
      RECT MASK 2 34.122 97.41 34.182 108.838 ;
      RECT MASK 2 34.396 97.41 34.456 108.838 ;
      RECT MASK 2 34.67 97.41 34.73 108.838 ;
      RECT MASK 2 34.944 97.41 35.004 108.838 ;
      RECT MASK 2 35.218 97.41 35.278 108.838 ;
      RECT MASK 2 35.492 97.41 35.552 108.838 ;
      RECT MASK 2 35.766 97.41 35.826 108.838 ;
      RECT MASK 2 36.04 97.41 36.1 108.838 ;
      RECT MASK 2 36.314 97.41 36.374 108.838 ;
      RECT MASK 2 36.588 97.41 36.648 108.838 ;
      RECT MASK 2 36.862 97.41 36.922 108.838 ;
      RECT MASK 2 37.136 97.41 37.196 108.838 ;
      RECT MASK 2 37.41 97.41 37.47 108.838 ;
      RECT MASK 2 37.684 97.41 37.744 108.838 ;
      RECT MASK 2 37.958 97.41 38.018 108.838 ;
      RECT MASK 2 38.232 97.41 38.292 108.838 ;
      RECT MASK 2 38.506 97.41 38.566 108.838 ;
      RECT MASK 2 38.78 97.41 38.84 108.838 ;
      RECT MASK 2 39.054 97.41 39.114 108.838 ;
      RECT MASK 2 39.328 97.41 39.388 108.838 ;
      RECT MASK 2 39.602 97.41 39.662 108.838 ;
      RECT MASK 2 39.876 97.41 39.936 108.838 ;
      RECT MASK 2 40.15 97.41 40.21 108.838 ;
      RECT MASK 2 40.424 97.41 40.484 108.838 ;
      RECT MASK 2 40.698 97.41 40.758 108.838 ;
      RECT MASK 2 40.972 97.41 41.032 108.838 ;
      RECT MASK 2 41.246 97.41 41.306 108.838 ;
      RECT MASK 2 41.52 97.41 41.58 108.838 ;
      RECT MASK 2 41.794 97.41 41.854 108.838 ;
      RECT MASK 2 42.068 97.41 42.128 108.838 ;
      RECT MASK 2 42.342 97.41 42.402 108.838 ;
      RECT MASK 2 42.616 97.41 42.676 108.838 ;
      RECT MASK 2 42.89 97.41 42.95 108.838 ;
      RECT MASK 2 43.164 97.41 43.224 108.838 ;
      RECT MASK 2 43.438 97.41 43.498 108.838 ;
      RECT MASK 2 45.73 97.41 45.79 108.838 ;
      RECT MASK 2 46.004 97.41 46.064 108.838 ;
      RECT MASK 2 46.278 97.41 46.338 108.838 ;
      RECT MASK 2 46.552 97.41 46.612 108.838 ;
      RECT MASK 2 46.826 97.41 46.886 108.838 ;
      RECT MASK 2 47.1 97.41 47.16 108.838 ;
      RECT MASK 2 47.374 97.41 47.434 108.838 ;
      RECT MASK 2 47.648 97.41 47.708 108.838 ;
      RECT MASK 2 47.922 97.41 47.982 108.838 ;
      RECT MASK 2 48.196 97.41 48.256 108.838 ;
      RECT MASK 2 48.47 97.41 48.53 108.838 ;
      RECT MASK 2 48.744 97.41 48.804 108.838 ;
      RECT MASK 2 49.018 97.41 49.078 108.838 ;
      RECT MASK 2 49.292 97.41 49.352 108.838 ;
      RECT MASK 2 49.566 97.41 49.626 108.838 ;
      RECT MASK 2 49.84 97.41 49.9 108.838 ;
      RECT MASK 2 50.114 97.41 50.174 108.838 ;
      RECT MASK 2 50.388 97.41 50.448 108.838 ;
      RECT MASK 2 50.662 97.41 50.722 108.838 ;
      RECT MASK 2 50.936 97.41 50.996 108.838 ;
      RECT MASK 2 51.21 97.41 51.27 108.838 ;
      RECT MASK 2 51.484 97.41 51.544 108.838 ;
      RECT MASK 2 51.758 97.41 51.818 108.838 ;
      RECT MASK 2 52.032 97.41 52.092 108.838 ;
      RECT MASK 2 52.306 97.41 52.366 108.838 ;
      RECT MASK 2 52.58 97.41 52.64 108.838 ;
      RECT MASK 2 52.854 97.41 52.914 108.838 ;
      RECT MASK 2 53.128 97.41 53.188 108.838 ;
      RECT MASK 2 53.402 97.41 53.462 108.838 ;
      RECT MASK 2 53.676 97.41 53.736 108.838 ;
      RECT MASK 2 53.95 97.41 54.01 108.838 ;
      RECT MASK 2 54.224 97.41 54.284 108.838 ;
      RECT MASK 2 54.498 97.41 54.558 108.838 ;
      RECT MASK 2 54.772 97.41 54.832 108.838 ;
      RECT MASK 2 55.046 97.41 55.106 108.838 ;
      RECT MASK 2 55.32 97.41 55.38 108.838 ;
      RECT MASK 2 55.594 97.41 55.654 108.838 ;
      RECT MASK 2 55.868 97.41 55.928 108.838 ;
      RECT MASK 2 56.142 97.41 56.202 108.838 ;
      RECT MASK 2 56.416 97.41 56.476 108.838 ;
      RECT MASK 2 56.69 97.41 56.75 108.838 ;
      RECT MASK 2 56.964 97.41 57.024 108.838 ;
      RECT MASK 2 57.238 97.41 57.298 108.838 ;
      RECT MASK 2 57.512 97.41 57.572 108.838 ;
      RECT MASK 2 57.786 97.41 57.846 108.838 ;
      RECT MASK 2 58.06 97.41 58.12 108.838 ;
      RECT MASK 2 58.334 97.41 58.394 108.838 ;
      RECT MASK 2 58.608 97.41 58.668 108.838 ;
      RECT MASK 2 58.882 97.41 58.942 108.838 ;
      RECT MASK 2 59.156 97.41 59.216 108.838 ;
      RECT MASK 2 59.43 97.41 59.49 108.838 ;
      RECT MASK 2 59.704 97.41 59.764 108.838 ;
      RECT MASK 2 59.978 97.41 60.038 108.838 ;
      RECT MASK 2 60.252 97.41 60.312 108.838 ;
      RECT MASK 2 60.526 97.41 60.586 108.838 ;
      RECT MASK 2 60.8 97.41 60.86 108.838 ;
      RECT MASK 2 61.074 97.41 61.134 108.838 ;
      RECT MASK 2 61.348 97.41 61.408 108.838 ;
      RECT MASK 2 61.622 97.41 61.682 108.838 ;
      RECT MASK 2 61.896 97.41 61.956 108.838 ;
      RECT MASK 2 62.17 97.41 62.23 108.838 ;
      RECT MASK 2 62.444 97.41 62.504 108.838 ;
      RECT MASK 2 62.718 97.41 62.778 108.838 ;
      RECT MASK 2 62.992 97.41 63.052 108.838 ;
      RECT MASK 2 63.266 97.41 63.326 108.838 ;
      RECT MASK 2 63.54 97.41 63.6 108.838 ;
      RECT MASK 2 63.814 97.41 63.874 108.838 ;
      RECT MASK 2 64.088 97.41 64.148 108.838 ;
      RECT MASK 2 64.362 97.41 64.422 108.838 ;
      RECT MASK 2 64.636 97.41 64.696 108.838 ;
      RECT MASK 2 64.91 97.41 64.97 108.838 ;
      RECT MASK 2 65.184 97.41 65.244 108.838 ;
      RECT MASK 2 65.458 97.41 65.518 108.838 ;
      RECT MASK 2 65.732 97.41 65.792 108.838 ;
      RECT MASK 2 66.006 97.41 66.066 108.838 ;
      RECT MASK 2 66.28 97.41 66.34 108.838 ;
      RECT MASK 2 66.554 97.41 66.614 108.838 ;
      RECT MASK 2 66.828 97.41 66.888 108.838 ;
      RECT MASK 2 67.102 97.41 67.162 108.838 ;
      RECT MASK 2 67.376 97.41 67.436 108.838 ;
      RECT MASK 2 67.65 97.41 67.71 108.838 ;
      RECT MASK 2 67.924 97.41 67.984 108.838 ;
      RECT MASK 2 68.198 97.41 68.258 108.838 ;
      RECT MASK 2 68.472 97.41 68.532 108.838 ;
      RECT MASK 2 68.746 97.41 68.806 108.838 ;
      RECT MASK 2 69.02 97.41 69.08 108.838 ;
      RECT MASK 2 69.294 97.41 69.354 108.838 ;
      RECT MASK 2 69.568 97.41 69.628 108.838 ;
      RECT MASK 2 69.842 97.41 69.902 108.838 ;
      RECT MASK 2 70.116 97.41 70.176 108.838 ;
      RECT MASK 2 70.39 97.41 70.45 108.838 ;
      RECT MASK 2 70.664 97.41 70.724 108.838 ;
      RECT MASK 2 70.938 97.41 70.998 108.838 ;
      RECT MASK 2 71.212 97.41 71.272 108.838 ;
      RECT MASK 2 71.486 97.41 71.546 108.838 ;
      RECT MASK 2 71.76 97.41 71.82 108.838 ;
      RECT MASK 2 72.034 97.41 72.094 108.838 ;
      RECT MASK 2 72.308 97.41 72.368 108.838 ;
      RECT MASK 2 72.582 97.41 72.642 108.838 ;
      RECT MASK 2 72.856 97.41 72.916 108.838 ;
      RECT MASK 2 73.13 97.41 73.19 108.838 ;
      RECT MASK 2 73.404 97.41 73.464 108.838 ;
      RECT MASK 2 73.678 97.41 73.738 108.838 ;
      RECT MASK 2 73.952 97.41 74.012 108.838 ;
      RECT MASK 2 74.226 97.41 74.286 108.838 ;
      RECT MASK 2 74.5 97.41 74.56 108.838 ;
      RECT MASK 2 74.774 97.41 74.834 108.838 ;
      RECT MASK 2 75.048 97.41 75.108 108.838 ;
      RECT MASK 2 75.322 97.41 75.382 108.838 ;
      RECT MASK 2 75.596 97.41 75.656 108.838 ;
      RECT MASK 2 75.87 97.41 75.93 108.838 ;
      RECT MASK 2 76.144 97.41 76.204 108.838 ;
      RECT MASK 2 76.418 97.41 76.478 108.838 ;
      RECT MASK 2 76.692 97.41 76.752 108.838 ;
      RECT MASK 2 76.966 97.41 77.026 108.838 ;
      RECT MASK 2 77.24 97.41 77.3 108.838 ;
      RECT MASK 2 77.514 97.41 77.574 108.838 ;
      RECT MASK 2 77.788 97.41 77.848 108.838 ;
      RECT MASK 2 78.062 97.41 78.122 108.838 ;
      RECT MASK 2 78.336 97.41 78.396 108.838 ;
      RECT MASK 2 78.61 97.41 78.67 108.838 ;
      RECT MASK 2 78.884 97.41 78.944 108.838 ;
      RECT MASK 2 79.158 97.41 79.218 108.838 ;
      RECT MASK 2 79.432 97.41 79.492 108.838 ;
      RECT MASK 2 79.706 97.41 79.766 108.838 ;
      RECT MASK 2 79.98 97.41 80.04 108.838 ;
      RECT MASK 2 80.254 97.41 80.314 108.838 ;
      RECT MASK 2 80.528 97.41 80.588 108.838 ;
      RECT MASK 2 80.802 97.41 80.862 108.838 ;
      RECT MASK 2 81.076 97.41 81.136 108.838 ;
      RECT MASK 2 81.35 97.41 81.41 108.838 ;
      RECT MASK 2 81.624 97.41 81.684 108.838 ;
      RECT MASK 2 81.898 97.41 81.958 108.838 ;
      RECT MASK 2 82.172 97.41 82.232 108.838 ;
      RECT MASK 2 82.446 97.41 82.506 108.838 ;
      RECT MASK 2 82.72 97.41 82.78 108.838 ;
      RECT MASK 2 82.994 97.41 83.054 108.838 ;
      RECT MASK 2 83.268 97.41 83.328 108.838 ;
      RECT MASK 2 83.542 97.41 83.602 108.838 ;
      RECT MASK 2 83.816 97.41 83.876 108.838 ;
      RECT MASK 2 84.09 97.41 84.15 108.838 ;
      RECT MASK 2 84.364 97.41 84.424 108.838 ;
      RECT MASK 2 84.638 97.41 84.698 108.838 ;
      RECT MASK 2 84.912 97.41 84.972 108.838 ;
      RECT MASK 2 85.186 97.41 85.246 108.838 ;
      RECT MASK 2 85.46 97.41 85.52 108.838 ;
      RECT MASK 2 85.734 97.41 85.794 108.838 ;
      RECT MASK 2 86.008 97.41 86.068 108.838 ;
      RECT MASK 2 86.282 97.41 86.342 108.838 ;
      RECT MASK 2 86.556 97.41 86.616 108.838 ;
      RECT MASK 2 86.83 97.41 86.89 108.838 ;
      RECT MASK 2 89.089 97.41 89.149 108.838 ;
      RECT MASK 2 89.363 97.41 89.423 108.838 ;
      RECT MASK 2 89.637 97.41 89.697 108.838 ;
      RECT MASK 2 89.911 97.41 89.971 108.838 ;
      RECT MASK 2 90.185 97.41 90.245 108.838 ;
      RECT MASK 2 90.459 97.41 90.519 108.838 ;
      RECT MASK 2 90.733 97.41 90.793 108.838 ;
      RECT MASK 2 91.007 97.41 91.067 108.838 ;
      RECT MASK 2 91.281 97.41 91.341 108.838 ;
      RECT MASK 2 91.555 97.41 91.615 108.838 ;
      RECT MASK 2 91.829 97.41 91.889 108.838 ;
      RECT MASK 2 92.103 97.41 92.163 108.838 ;
      RECT MASK 2 92.377 97.41 92.437 108.838 ;
      RECT MASK 2 92.651 97.41 92.711 108.838 ;
      RECT MASK 2 92.925 97.41 92.985 108.838 ;
      RECT MASK 2 93.199 97.41 93.259 108.838 ;
      RECT MASK 2 93.473 97.41 93.533 108.838 ;
      RECT MASK 2 93.747 97.41 93.807 108.838 ;
      RECT MASK 2 94.021 97.41 94.081 108.838 ;
      RECT MASK 2 94.295 97.41 94.355 108.838 ;
      RECT MASK 2 94.569 97.41 94.629 108.838 ;
      RECT MASK 2 94.843 97.41 94.903 108.838 ;
      RECT MASK 2 95.117 97.41 95.177 108.838 ;
      RECT MASK 2 95.391 97.41 95.451 108.838 ;
      RECT MASK 2 95.665 97.41 95.725 108.838 ;
      RECT MASK 2 95.939 97.41 95.999 108.838 ;
      RECT MASK 2 96.213 97.41 96.273 108.838 ;
      RECT MASK 2 96.487 97.41 96.547 108.838 ;
      RECT MASK 2 96.761 97.41 96.821 108.838 ;
      RECT MASK 2 97.035 97.41 97.095 108.838 ;
      RECT MASK 2 97.309 97.41 97.369 108.838 ;
      RECT MASK 2 97.583 97.41 97.643 108.838 ;
      RECT MASK 2 97.857 97.41 97.917 108.838 ;
      RECT MASK 2 98.131 97.41 98.191 108.838 ;
      RECT MASK 2 98.405 97.41 98.465 108.838 ;
      RECT MASK 2 98.679 97.41 98.739 108.838 ;
      RECT MASK 2 98.953 97.41 99.013 108.838 ;
      RECT MASK 2 99.227 97.41 99.287 108.838 ;
      RECT MASK 2 99.501 97.41 99.561 108.838 ;
      RECT MASK 2 99.775 97.41 99.835 108.838 ;
      RECT MASK 2 100.049 97.41 100.109 108.838 ;
      RECT MASK 2 100.323 97.41 100.383 108.838 ;
      RECT MASK 2 100.597 97.41 100.657 108.838 ;
      RECT MASK 2 100.871 97.41 100.931 108.838 ;
      RECT MASK 2 101.145 97.41 101.205 108.838 ;
      RECT MASK 2 101.419 97.41 101.479 108.838 ;
      RECT MASK 2 101.693 97.41 101.753 108.838 ;
      RECT MASK 2 101.967 97.41 102.027 108.838 ;
      RECT MASK 2 102.241 97.41 102.301 108.838 ;
      RECT MASK 2 102.515 97.41 102.575 108.838 ;
      RECT MASK 2 102.789 97.41 102.849 108.838 ;
      RECT MASK 2 103.063 97.41 103.123 108.838 ;
      RECT MASK 2 103.337 97.41 103.397 108.838 ;
      RECT MASK 2 103.611 97.41 103.671 108.838 ;
      RECT MASK 2 103.885 97.41 103.945 108.838 ;
      RECT MASK 2 104.159 97.41 104.219 108.838 ;
      RECT MASK 2 104.433 97.41 104.493 108.838 ;
      RECT MASK 2 104.707 97.41 104.767 108.838 ;
      RECT MASK 2 104.981 97.41 105.041 108.838 ;
      RECT MASK 2 105.255 97.41 105.315 108.838 ;
      RECT MASK 2 105.529 97.41 105.589 108.838 ;
      RECT MASK 2 105.803 97.41 105.863 108.838 ;
      RECT MASK 2 106.077 97.41 106.137 108.838 ;
      RECT MASK 2 106.351 97.41 106.411 108.838 ;
      RECT MASK 2 106.625 97.41 106.685 108.838 ;
      RECT MASK 2 106.899 97.41 106.959 108.838 ;
      RECT MASK 2 107.173 97.41 107.233 108.838 ;
      RECT MASK 2 107.447 97.41 107.507 108.838 ;
      RECT MASK 2 107.721 97.41 107.781 108.838 ;
      RECT MASK 2 107.995 97.41 108.055 108.838 ;
      RECT MASK 2 108.269 97.41 108.329 108.838 ;
      RECT MASK 2 108.543 97.41 108.603 108.838 ;
      RECT MASK 2 108.817 97.41 108.877 108.838 ;
      RECT MASK 2 109.091 97.41 109.151 108.838 ;
      RECT MASK 2 109.365 97.41 109.425 108.838 ;
      RECT MASK 2 109.639 97.41 109.699 108.838 ;
      RECT MASK 2 109.913 97.41 109.973 108.838 ;
      RECT MASK 2 110.187 97.41 110.247 108.838 ;
      RECT MASK 2 110.461 97.41 110.521 108.838 ;
      RECT MASK 2 110.735 97.41 110.795 108.838 ;
      RECT MASK 2 111.009 97.41 111.069 108.838 ;
      RECT MASK 2 111.283 97.41 111.343 108.838 ;
      RECT MASK 2 111.557 97.41 111.617 108.838 ;
      RECT MASK 2 111.831 97.41 111.891 108.838 ;
      RECT MASK 2 112.105 97.41 112.165 108.838 ;
      RECT MASK 2 112.379 97.41 112.439 108.838 ;
      RECT MASK 2 112.653 97.41 112.713 108.838 ;
      RECT MASK 2 112.927 97.41 112.987 108.838 ;
      RECT MASK 2 113.201 97.41 113.261 108.838 ;
      RECT MASK 2 113.475 97.41 113.535 108.838 ;
      RECT MASK 2 113.749 97.41 113.809 108.838 ;
      RECT MASK 2 114.023 97.41 114.083 108.838 ;
      RECT MASK 2 114.297 97.41 114.357 108.838 ;
      RECT MASK 2 114.571 97.41 114.631 108.838 ;
      RECT MASK 2 114.845 97.41 114.905 108.838 ;
      RECT MASK 2 115.119 97.41 115.179 108.838 ;
      RECT MASK 2 115.393 97.41 115.453 108.838 ;
      RECT MASK 2 115.667 97.41 115.727 108.838 ;
      RECT MASK 2 115.941 97.41 116.001 108.838 ;
      RECT MASK 2 116.215 97.41 116.275 108.838 ;
      RECT MASK 2 116.489 97.41 116.549 108.838 ;
      RECT MASK 2 116.763 97.41 116.823 108.838 ;
      RECT MASK 2 117.037 97.41 117.097 108.838 ;
      RECT MASK 2 117.311 97.41 117.371 108.838 ;
      RECT MASK 2 117.585 97.41 117.645 108.838 ;
      RECT MASK 2 117.859 97.41 117.919 108.838 ;
      RECT MASK 2 118.133 97.41 118.193 108.838 ;
      RECT MASK 2 118.407 97.41 118.467 108.838 ;
      RECT MASK 2 118.681 97.41 118.741 108.838 ;
      RECT MASK 2 118.955 97.41 119.015 108.838 ;
      RECT MASK 2 119.229 97.41 119.289 108.838 ;
      RECT MASK 2 119.503 97.41 119.563 108.838 ;
      RECT MASK 2 119.777 97.41 119.837 108.838 ;
      RECT MASK 2 120.051 97.41 120.111 108.838 ;
      RECT MASK 2 120.325 97.41 120.385 108.838 ;
      RECT MASK 2 120.599 97.41 120.659 108.838 ;
      RECT MASK 2 120.873 97.41 120.933 108.838 ;
      RECT MASK 2 121.147 97.41 121.207 108.838 ;
      RECT MASK 2 121.421 97.41 121.481 108.838 ;
      RECT MASK 2 121.695 97.41 121.755 108.838 ;
      RECT MASK 2 121.969 97.41 122.029 108.838 ;
      RECT MASK 2 122.243 97.41 122.303 108.838 ;
      RECT MASK 2 122.517 97.41 122.577 108.838 ;
      RECT MASK 2 122.791 97.41 122.851 108.838 ;
      RECT MASK 2 123.065 97.41 123.125 108.838 ;
      RECT MASK 2 123.339 97.41 123.399 108.838 ;
      RECT MASK 2 123.613 97.41 123.673 108.838 ;
      RECT MASK 2 123.887 97.41 123.947 108.838 ;
      RECT MASK 2 124.161 97.41 124.221 108.838 ;
      RECT MASK 2 124.435 97.41 124.495 108.838 ;
      RECT MASK 2 124.709 97.41 124.769 108.838 ;
      RECT MASK 2 124.983 97.41 125.043 108.838 ;
      RECT MASK 2 125.257 97.41 125.317 108.838 ;
      RECT MASK 2 125.531 97.41 125.591 108.838 ;
      RECT MASK 2 125.805 97.41 125.865 108.838 ;
      RECT MASK 2 126.079 97.41 126.139 108.838 ;
      RECT MASK 2 126.353 97.41 126.413 108.838 ;
      RECT MASK 2 126.627 97.41 126.687 108.838 ;
      RECT MASK 2 126.901 97.41 126.961 108.838 ;
      RECT MASK 2 127.175 97.41 127.235 108.838 ;
      RECT MASK 2 127.449 97.41 127.509 108.838 ;
    LAYER M4 SPACING 0 ;
      RECT 0 0 130.416 109.44 ;
      RECT MASK 1 54.1255 11.218 127.698 11.298 ;
      RECT MASK 1 32.335 86.35 32.735 95.33 ;
      RECT MASK 1 35.562 86.35 67.24 86.71 ;
      RECT MASK 1 71.952 86.35 103.63 86.71 ;
      RECT MASK 1 25.387 87.081 31.9635 87.543 ;
      RECT MASK 1 37.021 87.89 65.781 88.39 ;
      RECT MASK 1 73.412 87.89 102.17 88.39 ;
      RECT MASK 1 25.6065 88.05 31.963 88.13 ;
      RECT MASK 1 25.387 89.458 31.963 89.92 ;
      RECT MASK 1 37.021 89.69 65.781 90.19 ;
      RECT MASK 1 73.412 89.69 102.17 90.19 ;
      RECT MASK 1 37.021 91.49 65.781 91.99 ;
      RECT MASK 1 73.412 91.49 102.17 91.99 ;
      RECT MASK 1 25.237 91.919 31.963 92.31 ;
      RECT MASK 1 37.021 93.29 65.781 93.79 ;
      RECT MASK 1 73.412 93.29 102.17 93.79 ;
      RECT MASK 1 25.237 93.748 31.961 94.134 ;
      RECT MASK 1 35.562 94.97 67.24 95.33 ;
      RECT MASK 1 71.952 94.97 103.63 95.33 ;
      RECT MASK 1 25.6665 95.25 31.9625 95.33 ;
      RECT MASK 1 4.371 95.28 4.481 95.3 ;
      RECT MASK 1 31.6175 95.64 107.542 95.82 ;
      RECT MASK 2 18.1755 86.43 31.963 86.821 ;
      RECT MASK 2 36.328 86.99 66.474 87.49 ;
      RECT MASK 2 72.718 86.99 102.864 87.49 ;
      RECT MASK 2 25.387 88.52 31.9635 88.982 ;
      RECT MASK 2 36.328 88.79 66.474 89.29 ;
      RECT MASK 2 72.718 88.79 102.864 89.29 ;
      RECT MASK 2 36.328 90.59 66.474 91.09 ;
      RECT MASK 2 72.718 90.59 102.864 91.09 ;
      RECT MASK 2 25.387 90.897 31.963 91.359 ;
      RECT MASK 2 36.328 92.39 66.474 92.89 ;
      RECT MASK 2 72.718 92.39 102.864 92.89 ;
      RECT MASK 2 36.328 94.19 66.474 94.69 ;
      RECT MASK 2 72.718 94.19 102.864 94.69 ;
    LAYER M5 SPACING 0 ;
      POLYGON 130.416 0 130.416 109.44 5.5175 109.44 5.5175 109.36 5.4375 109.36 5.4375 109.44 4.7765 109.44 4.7765 109.36 4.6965 109.36 4.6965 109.44 4.1955 109.44 4.1955 109.36 4.1155 109.36 4.1155 109.44 4.0355 109.44 4.0355 109.36 3.9555 109.36 3.9555 109.44 3.4545 109.44 3.4545 109.36 3.3745 109.36 3.3745 109.44 3.2945 109.44 3.2945 109.36 3.2145 109.36 3.2145 109.44 2.7135 109.44 2.7135 109.36 2.6335 109.36 2.6335 109.44 2.5535 109.44 2.5535 109.36 2.4735 109.36 2.4735 109.44 1.9725 109.44 1.9725 109.36 1.8925 109.36 1.8925 109.44 1.8125 109.44 1.8125 109.36 1.7325 109.36 1.7325 109.44 1.2315 109.44 1.2315 109.36 1.1515 109.36 1.1515 109.44 1.0715 109.44 1.0715 109.36 0.9915 109.36 0.9915 109.44 0 109.44 0 0 ;
      RECT MASK 1 32.335 86.35 32.735 95.53 ;
      RECT MASK 1 33.135 86.35 33.535 95.53 ;
      RECT MASK 1 33.935 86.35 34.335 95.53 ;
      RECT MASK 1 34.735 86.35 35.135 95.53 ;
      RECT MASK 1 24.353 86.365 24.553 96.987 ;
    LAYER M6 SPACING 0 ;
      RECT 0 0 130.416 109.44 ;
      RECT MASK 1 24.017 86.35 69.396 86.71 ;
      RECT MASK 1 24.017 86.99 69.396 87.49 ;
      RECT MASK 1 24.017 88.79 69.396 89.29 ;
      RECT MASK 1 24.017 90.59 69.396 91.09 ;
      RECT MASK 1 24.017 92.39 69.396 92.89 ;
      RECT MASK 1 24.017 94.19 69.396 94.69 ;
      RECT MASK 1 24.017 94.97 69.396 95.33 ;
      RECT MASK 1 0.2 95.55 130.199 95.91 ;
    LAYER M7 SPACING 0 ;
      POLYGON 130.416 0 130.416 109.44 15.853 109.44 15.853 108.99 15.403 108.99 15.403 109.44 0 109.44 0 0 ;
    LAYER M8 SPACING 0 ;
      POLYGON 0 0 0 109.44 130.416 109.44 130.416 109.28 0.2 109.28 0.2 108.83 130.216 108.83 130.216 109.28 130.416 109.28 130.416 108.48 0.2 108.48 0.2 108.03 130.216 108.03 130.216 108.48 130.416 108.48 130.416 107.68 0.2 107.68 0.2 107.23 130.216 107.23 130.216 107.68 130.416 107.68 130.416 106.88 0.2 106.88 0.2 106.43 130.216 106.43 130.216 106.88 130.416 106.88 130.416 106.08 0.2 106.08 0.2 105.63 130.216 105.63 130.216 106.08 130.416 106.08 130.416 105.28 0.2 105.28 0.2 104.83 130.216 104.83 130.216 105.28 130.416 105.28 130.416 104.48 0.2 104.48 0.2 104.03 130.216 104.03 130.216 104.48 130.416 104.48 130.416 103.68 0.2 103.68 0.2 103.23 130.216 103.23 130.216 103.68 130.416 103.68 130.416 102.88 0.2 102.88 0.2 102.43 130.216 102.43 130.216 102.88 130.416 102.88 130.416 102.08 0.2 102.08 0.2 101.63 130.216 101.63 130.216 102.08 130.416 102.08 130.416 101.28 0.2 101.28 0.2 100.83 130.216 100.83 130.216 101.28 130.416 101.28 130.416 100.48 0.2 100.48 0.2 100.03 130.216 100.03 130.216 100.48 130.416 100.48 130.416 99.68 0.2 99.68 0.2 99.23 130.216 99.23 130.216 99.68 130.416 99.68 130.416 98.88 0.2 98.88 0.2 98.43 130.216 98.43 130.216 98.88 130.416 98.88 130.416 98.08 0.2 98.08 0.2 97.63 130.216 97.63 130.216 98.08 130.416 98.08 130.416 97.28 0.2 97.28 0.2 96.83 130.199 96.83 130.199 97.28 130.416 97.28 130.416 96.48 0.2 96.48 0.2 96.03 130.216 96.03 130.216 96.48 130.416 96.48 130.416 95.705 0.2 95.705 0.2 95.255 23.817 95.255 23.817 95.705 107.51 95.705 107.51 95.255 130.199 95.255 130.199 95.705 130.416 95.705 130.416 94.905 0.2 94.905 0.2 94.455 23.817 94.455 23.817 94.905 107.51 94.905 107.51 94.69 24.017 94.69 24.017 94.19 69.396 94.19 69.396 94.69 69.796 94.69 69.796 94.19 107.057 94.19 107.057 94.69 107.51 94.69 107.51 94.455 130.199 94.455 130.199 94.905 130.416 94.905 130.416 94.105 0.2 94.105 0.2 93.655 23.817 93.655 23.817 94.105 107.51 94.105 107.51 93.79 24.017 93.79 24.017 93.35 0.2 93.35 0.2 92.9 23.817 92.9 23.817 93.35 24.017 93.35 24.017 93.29 102.87 93.29 102.87 93.79 103.27 93.79 103.27 93.29 107.057 93.29 107.057 93.79 107.51 93.79 107.51 93.655 130.199 93.655 130.199 94.105 130.416 94.105 130.416 93.35 107.51 93.35 107.51 92.9 130.199 92.9 130.199 93.35 130.416 93.35 130.416 92.89 24.017 92.89 24.017 92.55 0.2 92.55 0.2 92.1 23.817 92.1 23.817 92.55 24.017 92.55 24.017 92.39 69.396 92.39 69.396 92.89 69.796 92.89 69.796 92.39 107.057 92.39 107.057 92.89 130.416 92.89 130.416 92.55 107.51 92.55 107.51 92.1 130.199 92.1 130.199 92.55 130.416 92.55 130.416 91.99 24.017 91.99 24.017 91.795 0.2 91.795 0.2 91.345 23.817 91.345 23.817 91.795 24.017 91.795 24.017 91.49 102.87 91.49 102.87 91.99 103.27 91.99 103.27 91.49 107.057 91.49 107.057 91.99 130.416 91.99 130.416 91.795 107.51 91.795 107.51 91.345 130.199 91.345 130.199 91.795 130.416 91.795 130.416 91.09 24.017 91.09 24.017 90.995 0.2 90.995 0.2 90.545 23.817 90.545 23.817 90.995 24.017 90.995 24.017 90.59 69.396 90.59 69.396 91.09 69.796 91.09 69.796 90.59 107.057 90.59 107.057 91.09 130.416 91.09 130.416 90.995 107.51 90.995 107.51 90.545 130.199 90.545 130.199 90.995 130.416 90.995 130.416 90.24 0.2 90.24 0.2 89.79 23.817 89.79 23.817 90.24 107.51 90.24 107.51 90.19 24.017 90.19 24.017 89.69 102.87 89.69 102.87 90.19 103.27 90.19 103.27 89.69 107.057 89.69 107.057 90.19 107.51 90.19 107.51 89.79 130.199 89.79 130.199 90.24 130.416 90.24 130.416 89.57 9.355 89.57 9.355 89.52 0.2 89.52 0.2 89.07 8.997 89.07 8.997 89.52 9.355 89.52 9.355 89.07 23.817 89.07 23.817 89.57 130.416 89.57 130.416 89.52 107.51 89.52 107.51 89.29 24.017 89.29 24.017 88.79 69.396 88.79 69.396 89.29 69.796 89.29 69.796 88.79 107.057 88.79 107.057 89.29 107.51 89.29 107.51 89.07 130.199 89.07 130.199 89.52 130.416 89.52 130.416 88.71 0.2 88.71 0.2 88.26 8.997 88.26 8.997 88.71 9.355 88.71 9.355 88.21 23.817 88.21 23.817 88.71 107.51 88.71 107.51 88.39 24.017 88.39 24.017 87.99 0.2 87.99 0.2 87.54 23.817 87.54 23.817 87.99 24.017 87.99 24.017 87.89 102.87 87.89 102.87 88.39 103.27 88.39 103.27 87.89 107.057 87.89 107.057 88.39 107.51 88.39 107.51 88.26 130.199 88.26 130.199 88.71 130.416 88.71 130.416 87.99 107.51 87.99 107.51 87.54 130.199 87.54 130.199 87.99 130.416 87.99 130.416 87.49 24.017 87.49 24.017 87.24 0.2 87.24 0.2 86.79 23.817 86.79 23.817 87.24 24.017 87.24 24.017 86.99 69.396 86.99 69.396 87.49 69.796 87.49 69.796 86.99 107.057 86.99 107.057 87.49 130.416 87.49 130.416 87.24 107.51 87.24 107.51 86.79 130.199 86.79 130.199 87.24 130.416 87.24 130.416 86.55 9.355 86.55 9.355 86.525 0.2 86.525 0.2 86.075 8.997 86.075 8.997 86.525 9.355 86.525 9.355 86.05 23.817 86.05 23.817 86.55 130.416 86.55 130.416 86.525 107.51 86.525 107.51 86.075 130.199 86.075 130.199 86.525 130.416 86.525 130.416 85.65 0.2 85.65 0.2 85.2 130.199 85.2 130.199 85.65 130.416 85.65 130.416 84.85 0.2 84.85 0.2 84.4 130.199 84.4 130.199 84.85 130.416 84.85 130.416 84.05 0.2 84.05 0.2 83.6 130.199 83.6 130.199 84.05 130.416 84.05 130.416 83.25 0.2 83.25 0.2 82.8 130.199 82.8 130.199 83.25 130.416 83.25 130.416 82.45 0.2 82.45 0.2 82 130.199 82 130.199 82.45 130.416 82.45 130.416 81.65 0.2 81.65 0.2 81.2 130.199 81.2 130.199 81.65 130.416 81.65 130.416 80.85 0.2 80.85 0.2 80.4 130.199 80.4 130.199 80.85 130.416 80.85 130.416 80.05 0.2 80.05 0.2 79.6 130.199 79.6 130.199 80.05 130.416 80.05 130.416 79.25 0.2 79.25 0.2 78.8 130.199 78.8 130.199 79.25 130.416 79.25 130.416 78.45 0.2 78.45 0.2 78 130.199 78 130.199 78.45 130.416 78.45 130.416 77.65 0.2 77.65 0.2 77.2 130.199 77.2 130.199 77.65 130.416 77.65 130.416 76.85 0.2 76.85 0.2 76.4 130.199 76.4 130.199 76.85 130.416 76.85 130.416 76.05 0.2 76.05 0.2 75.6 130.199 75.6 130.199 76.05 130.416 76.05 130.416 75.25 0.2 75.25 0.2 74.8 130.199 74.8 130.199 75.25 130.416 75.25 130.416 74.45 0.2 74.45 0.2 74 130.199 74 130.199 74.45 130.416 74.45 130.416 73.65 0.2 73.65 0.2 73.2 130.199 73.2 130.199 73.65 130.416 73.65 130.416 72.85 0.2 72.85 0.2 72.4 130.199 72.4 130.199 72.85 130.416 72.85 130.416 72.05 0.2 72.05 0.2 71.6 130.199 71.6 130.199 72.05 130.416 72.05 130.416 71.25 0.2 71.25 0.2 70.8 130.199 70.8 130.199 71.25 130.416 71.25 130.416 70.45 0.2 70.45 0.2 70 130.199 70 130.199 70.45 130.416 70.45 130.416 69.65 0.2 69.65 0.2 69.2 130.199 69.2 130.199 69.65 130.416 69.65 130.416 68.85 0.2 68.85 0.2 68.4 130.199 68.4 130.199 68.85 130.416 68.85 130.416 68.05 0.2 68.05 0.2 67.6 130.199 67.6 130.199 68.05 130.416 68.05 130.416 67.25 0.2 67.25 0.2 66.8 130.199 66.8 130.199 67.25 130.416 67.25 130.416 66.45 0.2 66.45 0.2 66 130.199 66 130.199 66.45 130.416 66.45 130.416 65.65 0.2 65.65 0.2 65.2 130.199 65.2 130.199 65.65 130.416 65.65 130.416 64.85 0.2 64.85 0.2 64.4 130.199 64.4 130.199 64.85 130.416 64.85 130.416 64.05 0.2 64.05 0.2 63.6 130.199 63.6 130.199 64.05 130.416 64.05 130.416 63.25 0.2 63.25 0.2 62.8 130.199 62.8 130.199 63.25 130.416 63.25 130.416 62.45 0.2 62.45 0.2 62 130.199 62 130.199 62.45 130.416 62.45 130.416 61.65 0.2 61.65 0.2 61.2 130.199 61.2 130.199 61.65 130.416 61.65 130.416 60.85 0.2 60.85 0.2 60.4 130.199 60.4 130.199 60.85 130.416 60.85 130.416 60.05 0.2 60.05 0.2 59.6 130.199 59.6 130.199 60.05 130.416 60.05 130.416 59.25 0.2 59.25 0.2 58.8 130.199 58.8 130.199 59.25 130.416 59.25 130.416 58.45 0.2 58.45 0.2 58 130.199 58 130.199 58.45 130.416 58.45 130.416 57.65 0.2 57.65 0.2 57.2 130.199 57.2 130.199 57.65 130.416 57.65 130.416 56.85 0.2 56.85 0.2 56.4 130.199 56.4 130.199 56.85 130.416 56.85 130.416 56.05 0.2 56.05 0.2 55.6 130.199 55.6 130.199 56.05 130.416 56.05 130.416 55.25 0.2 55.25 0.2 54.8 130.199 54.8 130.199 55.25 130.416 55.25 130.416 54.45 0.2 54.45 0.2 54 130.199 54 130.199 54.45 130.416 54.45 130.416 53.65 0.2 53.65 0.2 53.2 130.199 53.2 130.199 53.65 130.416 53.65 130.416 52.85 0.2 52.85 0.2 52.4 130.199 52.4 130.199 52.85 130.416 52.85 130.416 52.05 0.2 52.05 0.2 51.6 130.199 51.6 130.199 52.05 130.416 52.05 130.416 51.25 0.2 51.25 0.2 50.8 130.199 50.8 130.199 51.25 130.416 51.25 130.416 50.45 0.2 50.45 0.2 50 130.199 50 130.199 50.45 130.416 50.45 130.416 49.65 0.2 49.65 0.2 49.2 130.199 49.2 130.199 49.65 130.416 49.65 130.416 48.85 0.2 48.85 0.2 48.4 130.199 48.4 130.199 48.85 130.416 48.85 130.416 48.05 0.2 48.05 0.2 47.6 130.199 47.6 130.199 48.05 130.416 48.05 130.416 47.25 0.2 47.25 0.2 46.8 130.199 46.8 130.199 47.25 130.416 47.25 130.416 46.45 0.2 46.45 0.2 46 130.199 46 130.199 46.45 130.416 46.45 130.416 45.65 0.2 45.65 0.2 45.2 130.199 45.2 130.199 45.65 130.416 45.65 130.416 44.85 0.2 44.85 0.2 44.4 130.199 44.4 130.199 44.85 130.416 44.85 130.416 44.05 0.2 44.05 0.2 43.6 130.199 43.6 130.199 44.05 130.416 44.05 130.416 43.25 0.2 43.25 0.2 42.8 130.199 42.8 130.199 43.25 130.416 43.25 130.416 42.45 0.2 42.45 0.2 42 130.199 42 130.199 42.45 130.416 42.45 130.416 41.65 0.2 41.65 0.2 41.2 130.199 41.2 130.199 41.65 130.416 41.65 130.416 40.85 0.2 40.85 0.2 40.4 130.199 40.4 130.199 40.85 130.416 40.85 130.416 40.05 0.2 40.05 0.2 39.6 130.199 39.6 130.199 40.05 130.416 40.05 130.416 39.25 0.2 39.25 0.2 38.8 130.199 38.8 130.199 39.25 130.416 39.25 130.416 38.45 0.2 38.45 0.2 38 130.199 38 130.199 38.45 130.416 38.45 130.416 37.65 0.2 37.65 0.2 37.2 130.199 37.2 130.199 37.65 130.416 37.65 130.416 36.85 0.2 36.85 0.2 36.4 130.199 36.4 130.199 36.85 130.416 36.85 130.416 36.05 0.2 36.05 0.2 35.6 130.199 35.6 130.199 36.05 130.416 36.05 130.416 35.25 0.2 35.25 0.2 34.8 130.199 34.8 130.199 35.25 130.416 35.25 130.416 34.45 0.2 34.45 0.2 34 130.199 34 130.199 34.45 130.416 34.45 130.416 33.65 0.2 33.65 0.2 33.2 130.199 33.2 130.199 33.65 130.416 33.65 130.416 32.85 0.2 32.85 0.2 32.4 130.199 32.4 130.199 32.85 130.416 32.85 130.416 32.05 0.2 32.05 0.2 31.6 130.199 31.6 130.199 32.05 130.416 32.05 130.416 31.25 0.2 31.25 0.2 30.8 130.199 30.8 130.199 31.25 130.416 31.25 130.416 30.45 0.2 30.45 0.2 30 130.199 30 130.199 30.45 130.416 30.45 130.416 29.65 0.2 29.65 0.2 29.2 130.199 29.2 130.199 29.65 130.416 29.65 130.416 28.85 0.2 28.85 0.2 28.4 130.199 28.4 130.199 28.85 130.416 28.85 130.416 28.05 0.2 28.05 0.2 27.6 130.199 27.6 130.199 28.05 130.416 28.05 130.416 27.25 0.2 27.25 0.2 26.8 130.199 26.8 130.199 27.25 130.416 27.25 130.416 26.45 0.2 26.45 0.2 26 130.199 26 130.199 26.45 130.416 26.45 130.416 25.65 0.2 25.65 0.2 25.2 130.199 25.2 130.199 25.65 130.416 25.65 130.416 24.85 0.2 24.85 0.2 24.4 130.199 24.4 130.199 24.85 130.416 24.85 130.416 24.05 0.2 24.05 0.2 23.6 130.199 23.6 130.199 24.05 130.416 24.05 130.416 23.25 0.2 23.25 0.2 22.8 130.199 22.8 130.199 23.25 130.416 23.25 130.416 22.45 0.2 22.45 0.2 22 130.199 22 130.199 22.45 130.416 22.45 130.416 21.65 0.2 21.65 0.2 21.2 130.199 21.2 130.199 21.65 130.416 21.65 130.416 20.85 0.2 20.85 0.2 20.4 130.199 20.4 130.199 20.85 130.416 20.85 130.416 20.05 0.2 20.05 0.2 19.6 130.199 19.6 130.199 20.05 130.416 20.05 130.416 19.25 0.2 19.25 0.2 18.8 130.199 18.8 130.199 19.25 130.416 19.25 130.416 18.45 0.2 18.45 0.2 18 130.199 18 130.199 18.45 130.416 18.45 130.416 17.65 0.2 17.65 0.2 17.2 130.199 17.2 130.199 17.65 130.416 17.65 130.416 16.85 0.2 16.85 0.2 16.4 130.199 16.4 130.199 16.85 130.416 16.85 130.416 16.05 0.2 16.05 0.2 15.6 130.199 15.6 130.199 16.05 130.416 16.05 130.416 15.25 0.2 15.25 0.2 14.8 130.199 14.8 130.199 15.25 130.416 15.25 130.416 14.45 0.2 14.45 0.2 14 130.199 14 130.199 14.45 130.416 14.45 130.416 13.65 0.2 13.65 0.2 13.2 130.199 13.2 130.199 13.65 130.416 13.65 130.416 12.85 0.2 12.85 0.2 12.4 130.199 12.4 130.199 12.85 130.416 12.85 130.416 12.05 0.2 12.05 0.2 11.6 130.199 11.6 130.199 12.05 130.416 12.05 130.416 11.25 0.2 11.25 0.2 10.8 130.199 10.8 130.199 11.25 130.416 11.25 130.416 10.45 0.2 10.45 0.2 10 130.199 10 130.199 10.45 130.416 10.45 130.416 9.65 0.2 9.65 0.2 9.2 130.199 9.2 130.199 9.65 130.416 9.65 130.416 8.85 0.2 8.85 0.2 8.4 130.199 8.4 130.199 8.85 130.416 8.85 130.416 8.05 0.2 8.05 0.2 7.6 130.199 7.6 130.199 8.05 130.416 8.05 130.416 7.25 0.2 7.25 0.2 6.8 130.199 6.8 130.199 7.25 130.416 7.25 130.416 6.45 0.2 6.45 0.2 6 130.199 6 130.199 6.45 130.416 6.45 130.416 5.65 0.2 5.65 0.2 5.2 130.199 5.2 130.199 5.65 130.416 5.65 130.416 4.85 0.2 4.85 0.2 4.4 130.199 4.4 130.199 4.85 130.416 4.85 130.416 4.05 0.2 4.05 0.2 3.6 130.199 3.6 130.199 4.05 130.416 4.05 130.416 3.25 0.2 3.25 0.2 2.8 130.199 2.8 130.199 3.25 130.416 3.25 130.416 2.45 0.2 2.45 0.2 2 130.199 2 130.199 2.45 130.416 2.45 130.416 1.65 0.2 1.65 0.2 1.2 130.199 1.2 130.199 1.65 130.416 1.65 130.416 0.85 0.2 0.85 0.2 0.4 130.199 0.4 130.199 0.85 130.416 0.85 130.416 0 ;
    LAYER M0 SPACING 0 ;
      RECT 0 0 130.416 109.44 ;
      RECT MASK 1 57.7415 0.7 65.984 0.74 ;
      RECT MASK 1 65.0585 1.05 65.949 1.078 ;
      RECT MASK 1 49.9395 1.12 52.6895 1.16 ;
      RECT MASK 1 58.765 1.198 58.825 1.378 ;
      RECT MASK 1 59.223 1.198 59.283 1.378 ;
      RECT MASK 1 59.681 1.198 59.741 1.378 ;
      RECT MASK 1 60.826 1.198 60.886 1.378 ;
      RECT MASK 1 61.284 1.198 61.344 1.378 ;
      RECT MASK 1 61.742 1.198 61.802 1.378 ;
      RECT MASK 1 62.2 1.198 62.26 1.378 ;
      RECT MASK 1 62.658 1.198 62.718 1.378 ;
      RECT MASK 1 63.116 1.198 63.176 1.378 ;
      RECT MASK 1 63.803 1.198 63.863 1.378 ;
      RECT MASK 1 64.261 1.198 64.321 1.378 ;
      RECT MASK 1 64.719 1.198 64.779 1.378 ;
      RECT MASK 1 115.425 1.435 129.001 1.475 ;
      RECT MASK 1 57.789 1.4575 57.969 1.4975 ;
      RECT MASK 1 60.1675 1.4575 60.3475 1.4975 ;
      RECT MASK 1 65.575 1.4575 65.984 1.4975 ;
      RECT MASK 1 50.0575 1.46 50.5795 1.5 ;
      RECT MASK 1 50.7215 1.46 51.2435 1.5 ;
      RECT MASK 1 51.3855 1.46 51.9075 1.5 ;
      RECT MASK 1 52.0495 1.46 52.5715 1.5 ;
      RECT MASK 1 61.259 1.518 62.6185 1.558 ;
      RECT MASK 1 50.0985 1.62 50.529 1.66 ;
      RECT MASK 1 50.7625 1.62 51.193 1.66 ;
      RECT MASK 1 51.4265 1.62 51.857 1.66 ;
      RECT MASK 1 52.0905 1.62 52.521 1.66 ;
      RECT MASK 1 1.6805 1.63 10.7245 1.67 ;
      RECT MASK 1 11.1705 1.63 12.9295 1.67 ;
      RECT MASK 1 13.4005 1.63 21.7575 1.67 ;
      RECT MASK 1 25.1795 1.63 33.5365 1.67 ;
      RECT MASK 1 34.0075 1.63 35.7665 1.67 ;
      RECT MASK 1 36.2125 1.63 45.2565 1.67 ;
      RECT MASK 1 58.74 1.72 64.804 1.76 ;
      RECT MASK 1 115.45 1.7435 115.53 23.5765 ;
      RECT MASK 1 128.896 1.7435 128.976 23.5765 ;
      RECT MASK 1 50.0575 1.78 50.476 1.82 ;
      RECT MASK 1 50.7215 1.78 51.14 1.82 ;
      RECT MASK 1 51.3855 1.78 51.804 1.82 ;
      RECT MASK 1 52.0495 1.78 52.468 1.82 ;
      RECT MASK 1 22.2235 1.878 23.3235 1.902 ;
      RECT MASK 1 23.6135 1.878 24.7135 1.902 ;
      RECT MASK 1 116.154 1.89 116.214 2.94 ;
      RECT MASK 1 116.428 1.89 116.488 2.94 ;
      RECT MASK 1 116.702 1.89 116.762 2.94 ;
      RECT MASK 1 116.976 1.89 117.036 2.94 ;
      RECT MASK 1 117.25 1.89 117.31 2.94 ;
      RECT MASK 1 117.524 1.89 117.584 2.94 ;
      RECT MASK 1 117.798 1.89 117.858 2.94 ;
      RECT MASK 1 118.072 1.89 118.132 2.94 ;
      RECT MASK 1 118.346 1.89 118.406 2.94 ;
      RECT MASK 1 118.62 1.89 118.68 2.94 ;
      RECT MASK 1 118.894 1.89 118.954 2.94 ;
      RECT MASK 1 119.168 1.89 119.228 2.94 ;
      RECT MASK 1 119.442 1.89 119.502 2.94 ;
      RECT MASK 1 119.716 1.89 119.776 2.94 ;
      RECT MASK 1 119.99 1.89 120.05 2.94 ;
      RECT MASK 1 120.264 1.89 120.324 2.94 ;
      RECT MASK 1 120.538 1.89 120.598 2.94 ;
      RECT MASK 1 120.812 1.89 120.872 2.94 ;
      RECT MASK 1 121.086 1.89 121.146 2.94 ;
      RECT MASK 1 121.36 1.89 121.42 2.94 ;
      RECT MASK 1 121.634 1.89 121.694 2.94 ;
      RECT MASK 1 121.908 1.89 121.968 2.94 ;
      RECT MASK 1 122.182 1.89 122.242 2.94 ;
      RECT MASK 1 122.456 1.89 122.516 2.94 ;
      RECT MASK 1 122.73 1.89 122.79 2.94 ;
      RECT MASK 1 123.004 1.89 123.064 2.94 ;
      RECT MASK 1 123.278 1.89 123.338 2.94 ;
      RECT MASK 1 123.552 1.89 123.612 2.94 ;
      RECT MASK 1 123.826 1.89 123.886 2.94 ;
      RECT MASK 1 124.1 1.89 124.16 2.94 ;
      RECT MASK 1 124.374 1.89 124.434 2.94 ;
      RECT MASK 1 124.648 1.89 124.708 2.94 ;
      RECT MASK 1 124.922 1.89 124.982 2.94 ;
      RECT MASK 1 125.196 1.89 125.256 2.94 ;
      RECT MASK 1 125.47 1.89 125.53 2.94 ;
      RECT MASK 1 125.744 1.89 125.804 2.94 ;
      RECT MASK 1 126.018 1.89 126.078 2.94 ;
      RECT MASK 1 126.292 1.89 126.352 2.94 ;
      RECT MASK 1 126.566 1.89 126.626 2.94 ;
      RECT MASK 1 126.84 1.89 126.9 2.94 ;
      RECT MASK 1 127.114 1.89 127.174 2.94 ;
      RECT MASK 1 127.388 1.89 127.448 2.94 ;
      RECT MASK 1 127.662 1.89 127.722 2.94 ;
      RECT MASK 1 127.936 1.89 127.996 2.94 ;
      RECT MASK 1 128.21 1.89 128.27 2.94 ;
      RECT MASK 1 61.3835 1.922 62.743 1.962 ;
      RECT MASK 1 57.789 1.9825 57.969 2.0225 ;
      RECT MASK 1 50.0985 2.055 50.529 2.095 ;
      RECT MASK 1 50.7625 2.055 51.193 2.095 ;
      RECT MASK 1 51.4265 2.055 51.857 2.095 ;
      RECT MASK 1 52.0905 2.055 52.521 2.095 ;
      RECT MASK 1 58.765 2.102 58.825 2.282 ;
      RECT MASK 1 59.223 2.102 59.283 2.282 ;
      RECT MASK 1 59.681 2.102 59.741 2.282 ;
      RECT MASK 1 60.826 2.102 60.886 2.282 ;
      RECT MASK 1 61.284 2.102 61.344 2.282 ;
      RECT MASK 1 61.742 2.102 61.802 2.282 ;
      RECT MASK 1 62.2 2.102 62.26 2.282 ;
      RECT MASK 1 62.658 2.102 62.718 2.282 ;
      RECT MASK 1 63.116 2.102 63.176 2.282 ;
      RECT MASK 1 63.803 2.102 63.863 2.282 ;
      RECT MASK 1 64.261 2.102 64.321 2.282 ;
      RECT MASK 1 64.719 2.102 64.779 2.282 ;
      RECT MASK 1 60.1675 2.1025 60.3475 2.1425 ;
      RECT MASK 1 65.575 2.1025 65.984 2.1425 ;
      RECT MASK 1 46.6605 2.12 49.2605 2.14 ;
      RECT MASK 1 2.4035 2.128 2.4635 2.308 ;
      RECT MASK 1 2.8615 2.128 2.9215 2.309 ;
      RECT MASK 1 3.3195 2.128 3.3795 2.308 ;
      RECT MASK 1 3.5485 2.128 3.6085 2.308 ;
      RECT MASK 1 3.7775 2.128 3.8375 2.308 ;
      RECT MASK 1 4.0065 2.128 4.0665 2.308 ;
      RECT MASK 1 4.2355 2.128 4.2955 2.308 ;
      RECT MASK 1 4.4645 2.128 4.5245 2.308 ;
      RECT MASK 1 4.6935 2.128 4.7535 2.308 ;
      RECT MASK 1 4.9225 2.128 4.9825 2.308 ;
      RECT MASK 1 5.1515 2.128 5.2115 2.309 ;
      RECT MASK 1 5.6095 2.128 5.6695 2.308 ;
      RECT MASK 1 6.0675 2.128 6.1275 2.308 ;
      RECT MASK 1 6.5255 2.128 6.5855 2.308 ;
      RECT MASK 1 6.9835 2.128 7.0435 2.308 ;
      RECT MASK 1 7.4415 2.128 7.5015 2.308 ;
      RECT MASK 1 7.8995 2.128 7.9595 2.308 ;
      RECT MASK 1 8.3575 2.128 8.4175 2.308 ;
      RECT MASK 1 8.8155 2.128 8.8755 2.308 ;
      RECT MASK 1 9.0445 2.128 9.1045 2.308 ;
      RECT MASK 1 9.2735 2.128 9.3335 2.308 ;
      RECT MASK 1 9.5025 2.128 9.5625 2.308 ;
      RECT MASK 1 9.7315 2.128 9.7915 2.308 ;
      RECT MASK 1 11.3455 2.128 11.4055 2.308 ;
      RECT MASK 1 11.8035 2.128 11.8635 2.308 ;
      RECT MASK 1 12.2615 2.128 12.3215 2.308 ;
      RECT MASK 1 12.7195 2.128 12.7795 2.308 ;
      RECT MASK 1 14.5735 2.128 14.6335 2.308 ;
      RECT MASK 1 15.0315 2.128 15.0915 2.308 ;
      RECT MASK 1 15.4895 2.128 15.5495 2.308 ;
      RECT MASK 1 15.9475 2.128 16.0075 2.308 ;
      RECT MASK 1 16.4055 2.128 16.4655 2.308 ;
      RECT MASK 1 16.8635 2.128 16.9235 2.308 ;
      RECT MASK 1 17.3215 2.128 17.3815 2.308 ;
      RECT MASK 1 17.7795 2.128 17.8395 2.308 ;
      RECT MASK 1 18.2375 2.128 18.2975 2.308 ;
      RECT MASK 1 18.6955 2.128 18.7555 2.308 ;
      RECT MASK 1 19.1535 2.128 19.2135 2.308 ;
      RECT MASK 1 19.6115 2.128 19.6715 2.308 ;
      RECT MASK 1 20.0695 2.128 20.1295 2.308 ;
      RECT MASK 1 20.5275 2.128 20.5875 2.308 ;
      RECT MASK 1 20.9855 2.128 21.0455 2.308 ;
      RECT MASK 1 21.4435 2.128 21.5035 2.308 ;
      RECT MASK 1 25.4335 2.128 25.4935 2.308 ;
      RECT MASK 1 25.8915 2.128 25.9515 2.308 ;
      RECT MASK 1 26.3495 2.128 26.4095 2.308 ;
      RECT MASK 1 26.8075 2.128 26.8675 2.308 ;
      RECT MASK 1 27.2655 2.128 27.3255 2.308 ;
      RECT MASK 1 27.7235 2.128 27.7835 2.308 ;
      RECT MASK 1 28.1815 2.128 28.2415 2.308 ;
      RECT MASK 1 28.6395 2.128 28.6995 2.308 ;
      RECT MASK 1 29.0975 2.128 29.1575 2.308 ;
      RECT MASK 1 29.5555 2.128 29.6155 2.308 ;
      RECT MASK 1 30.0135 2.128 30.0735 2.308 ;
      RECT MASK 1 30.4715 2.128 30.5315 2.308 ;
      RECT MASK 1 30.9295 2.128 30.9895 2.308 ;
      RECT MASK 1 31.3875 2.128 31.4475 2.308 ;
      RECT MASK 1 31.8455 2.128 31.9055 2.308 ;
      RECT MASK 1 32.3035 2.128 32.3635 2.308 ;
      RECT MASK 1 34.1575 2.128 34.2175 2.308 ;
      RECT MASK 1 34.6155 2.128 34.6755 2.308 ;
      RECT MASK 1 35.0735 2.128 35.1335 2.308 ;
      RECT MASK 1 35.5315 2.128 35.5915 2.308 ;
      RECT MASK 1 37.1455 2.128 37.2055 2.308 ;
      RECT MASK 1 37.3745 2.128 37.4345 2.308 ;
      RECT MASK 1 37.6035 2.128 37.6635 2.308 ;
      RECT MASK 1 37.8325 2.128 37.8925 2.308 ;
      RECT MASK 1 38.0615 2.128 38.1215 2.308 ;
      RECT MASK 1 38.5195 2.128 38.5795 2.308 ;
      RECT MASK 1 38.9775 2.128 39.0375 2.308 ;
      RECT MASK 1 39.4355 2.128 39.4955 2.308 ;
      RECT MASK 1 39.8935 2.128 39.9535 2.308 ;
      RECT MASK 1 40.3515 2.128 40.4115 2.308 ;
      RECT MASK 1 40.8095 2.128 40.8695 2.308 ;
      RECT MASK 1 41.2675 2.128 41.3275 2.308 ;
      RECT MASK 1 41.7255 2.128 41.7855 2.309 ;
      RECT MASK 1 41.9545 2.128 42.0145 2.308 ;
      RECT MASK 1 42.1835 2.128 42.2435 2.308 ;
      RECT MASK 1 42.4125 2.128 42.4725 2.308 ;
      RECT MASK 1 42.6415 2.128 42.7015 2.308 ;
      RECT MASK 1 42.8705 2.128 42.9305 2.308 ;
      RECT MASK 1 43.0995 2.128 43.1595 2.308 ;
      RECT MASK 1 43.3285 2.128 43.3885 2.308 ;
      RECT MASK 1 43.5575 2.128 43.6175 2.308 ;
      RECT MASK 1 44.0155 2.128 44.0755 2.309 ;
      RECT MASK 1 44.4735 2.128 44.5335 2.308 ;
      RECT MASK 1 46.6605 2.2 49.2605 2.22 ;
      RECT MASK 1 50.055 2.215 50.586 2.255 ;
      RECT MASK 1 50.719 2.215 51.25 2.255 ;
      RECT MASK 1 51.383 2.215 51.914 2.255 ;
      RECT MASK 1 52.047 2.215 52.578 2.255 ;
      RECT MASK 1 22.4135 2.238 22.7135 2.262 ;
      RECT MASK 1 22.8235 2.238 23.1235 2.262 ;
      RECT MASK 1 23.8135 2.238 24.1135 2.262 ;
      RECT MASK 1 24.2235 2.238 24.5235 2.262 ;
      RECT MASK 1 46.6605 2.28 49.2605 2.3 ;
      RECT MASK 1 22.4135 2.328 22.7135 2.352 ;
      RECT MASK 1 22.8235 2.328 23.1235 2.352 ;
      RECT MASK 1 23.8135 2.328 24.1135 2.352 ;
      RECT MASK 1 24.2235 2.328 24.5235 2.352 ;
      RECT MASK 1 46.6605 2.36 49.2605 2.38 ;
      RECT MASK 1 10.3585 2.3875 10.5385 2.4275 ;
      RECT MASK 1 13.5865 2.3875 13.7665 2.4275 ;
      RECT MASK 1 33.1705 2.3875 33.3505 2.4275 ;
      RECT MASK 1 36.3985 2.3875 36.5785 2.4275 ;
      RECT MASK 1 65.0475 2.402 65.949 2.43 ;
      RECT MASK 1 22.4135 2.418 22.7135 2.442 ;
      RECT MASK 1 22.8235 2.418 23.1235 2.442 ;
      RECT MASK 1 23.8135 2.418 24.1135 2.442 ;
      RECT MASK 1 24.2235 2.418 24.5235 2.442 ;
      RECT MASK 1 46.6605 2.44 49.2605 2.46 ;
      RECT MASK 1 1.6135 2.4475 1.8575 2.4875 ;
      RECT MASK 1 45.0795 2.4475 45.3235 2.4875 ;
      RECT MASK 1 22.2135 2.508 23.3235 2.532 ;
      RECT MASK 1 23.6135 2.508 24.7235 2.532 ;
      RECT MASK 1 46.6605 2.52 49.2605 2.54 ;
      RECT MASK 1 2.5025 2.549 2.7175 2.589 ;
      RECT MASK 1 2.8365 2.549 4.196 2.589 ;
      RECT MASK 1 5.7055 2.549 8.57 2.589 ;
      RECT MASK 1 9.373 2.549 10.0665 2.589 ;
      RECT MASK 1 11.0705 2.549 11.764 2.589 ;
      RECT MASK 1 12.361 2.549 13.0765 2.589 ;
      RECT MASK 1 14.663 2.549 21.414 2.589 ;
      RECT MASK 1 25.523 2.549 32.274 2.589 ;
      RECT MASK 1 33.8605 2.549 34.576 2.589 ;
      RECT MASK 1 35.173 2.549 35.8665 2.589 ;
      RECT MASK 1 36.8705 2.549 37.564 2.589 ;
      RECT MASK 1 38.367 2.549 41.2315 2.589 ;
      RECT MASK 1 42.741 2.549 44.1005 2.589 ;
      RECT MASK 1 44.2195 2.549 44.4345 2.589 ;
      RECT MASK 1 49.9395 2.59 52.6895 2.63 ;
      RECT MASK 1 22.7735 2.598 23.299 2.622 ;
      RECT MASK 1 23.684 2.598 24.1635 2.622 ;
      RECT MASK 1 46.6605 2.6 49.2605 2.62 ;
      RECT MASK 1 62.5395 2.61 62.743 2.638 ;
      RECT MASK 1 65.839 2.61 66.042 2.638 ;
      RECT MASK 1 2.5025 2.751 2.7175 2.791 ;
      RECT MASK 1 3.5235 2.751 9.692 2.791 ;
      RECT MASK 1 10.9455 2.751 11.764 2.791 ;
      RECT MASK 1 14.663 2.751 21.414 2.791 ;
      RECT MASK 1 25.523 2.751 32.274 2.791 ;
      RECT MASK 1 35.173 2.751 35.9915 2.791 ;
      RECT MASK 1 37.245 2.751 43.4135 2.791 ;
      RECT MASK 1 44.2195 2.751 44.4345 2.791 ;
      RECT MASK 1 58.536 2.758 58.596 2.938 ;
      RECT MASK 1 58.994 2.758 59.054 2.938 ;
      RECT MASK 1 59.452 2.758 59.512 2.938 ;
      RECT MASK 1 59.91 2.758 59.97 2.938 ;
      RECT MASK 1 60.368 2.758 60.428 2.938 ;
      RECT MASK 1 62.887 2.758 62.947 2.938 ;
      RECT MASK 1 63.345 2.758 63.405 2.938 ;
      RECT MASK 1 63.803 2.758 63.863 2.938 ;
      RECT MASK 1 64.261 2.758 64.321 2.938 ;
      RECT MASK 1 64.719 2.758 64.779 2.938 ;
      RECT MASK 1 65.177 2.758 65.237 2.938 ;
      RECT MASK 1 65.635 2.758 65.695 2.938 ;
      RECT MASK 1 46.6605 2.84 49.2605 2.86 ;
      RECT MASK 1 1.6135 2.8525 1.8575 2.8925 ;
      RECT MASK 1 45.0795 2.8525 45.3235 2.8925 ;
      RECT MASK 1 60.995 2.8975 61.404 2.9375 ;
      RECT MASK 1 61.911 2.8975 62.091 2.9375 ;
      RECT MASK 1 10.107 2.9125 10.7505 2.9525 ;
      RECT MASK 1 13.5865 2.9125 13.7665 2.9525 ;
      RECT MASK 1 33.1705 2.9125 33.3505 2.9525 ;
      RECT MASK 1 36.3985 2.9125 36.5785 2.9525 ;
      RECT MASK 1 46.6605 2.92 49.2605 2.94 ;
      RECT MASK 1 22.2135 2.958 23.3235 2.982 ;
      RECT MASK 1 23.6135 2.958 24.7235 2.982 ;
      RECT MASK 1 46.6605 3 49.2605 3.02 ;
      RECT MASK 1 49.9395 3.01 52.6895 3.05 ;
      RECT MASK 1 57.789 3.0175 57.969 3.0575 ;
      RECT MASK 1 2.4035 3.032 2.4635 3.212 ;
      RECT MASK 1 2.8615 3.032 2.9215 3.212 ;
      RECT MASK 1 3.3195 3.032 3.3795 3.212 ;
      RECT MASK 1 3.5485 3.032 3.6085 3.212 ;
      RECT MASK 1 3.7775 3.032 3.8375 3.212 ;
      RECT MASK 1 4.0065 3.032 4.0665 3.212 ;
      RECT MASK 1 4.2355 3.032 4.2955 3.212 ;
      RECT MASK 1 4.4645 3.032 4.5245 3.212 ;
      RECT MASK 1 4.6935 3.032 4.7535 3.212 ;
      RECT MASK 1 4.9225 3.032 4.9825 3.212 ;
      RECT MASK 1 5.1515 3.032 5.2115 3.212 ;
      RECT MASK 1 5.6095 3.032 5.6695 3.212 ;
      RECT MASK 1 6.0675 3.032 6.1275 3.212 ;
      RECT MASK 1 6.5255 3.032 6.5855 3.212 ;
      RECT MASK 1 6.9835 3.032 7.0435 3.212 ;
      RECT MASK 1 7.4415 3.032 7.5015 3.212 ;
      RECT MASK 1 7.8995 3.032 7.9595 3.212 ;
      RECT MASK 1 8.3575 3.032 8.4175 3.212 ;
      RECT MASK 1 8.8155 3.032 8.8755 3.212 ;
      RECT MASK 1 9.0445 3.032 9.1045 3.212 ;
      RECT MASK 1 9.2735 3.032 9.3335 3.212 ;
      RECT MASK 1 9.5025 3.032 9.5625 3.212 ;
      RECT MASK 1 9.7315 3.032 9.7915 3.212 ;
      RECT MASK 1 11.3455 3.032 11.4055 3.212 ;
      RECT MASK 1 11.8035 3.032 11.8635 3.212 ;
      RECT MASK 1 12.2615 3.032 12.3215 3.212 ;
      RECT MASK 1 12.7195 3.032 12.7795 3.212 ;
      RECT MASK 1 14.5735 3.032 14.6335 3.212 ;
      RECT MASK 1 15.0315 3.032 15.0915 3.212 ;
      RECT MASK 1 15.4895 3.032 15.5495 3.212 ;
      RECT MASK 1 15.9475 3.032 16.0075 3.212 ;
      RECT MASK 1 16.4055 3.032 16.4655 3.212 ;
      RECT MASK 1 16.8635 3.032 16.9235 3.212 ;
      RECT MASK 1 17.3215 3.032 17.3815 3.212 ;
      RECT MASK 1 17.7795 3.032 17.8395 3.212 ;
      RECT MASK 1 18.2375 3.032 18.2975 3.212 ;
      RECT MASK 1 18.6955 3.032 18.7555 3.212 ;
      RECT MASK 1 19.1535 3.032 19.2135 3.212 ;
      RECT MASK 1 19.6115 3.032 19.6715 3.212 ;
      RECT MASK 1 20.0695 3.032 20.1295 3.212 ;
      RECT MASK 1 20.5275 3.032 20.5875 3.212 ;
      RECT MASK 1 20.9855 3.032 21.0455 3.212 ;
      RECT MASK 1 21.4435 3.032 21.5035 3.212 ;
      RECT MASK 1 25.4335 3.032 25.4935 3.212 ;
      RECT MASK 1 25.8915 3.032 25.9515 3.212 ;
      RECT MASK 1 26.3495 3.032 26.4095 3.212 ;
      RECT MASK 1 26.8075 3.032 26.8675 3.212 ;
      RECT MASK 1 27.2655 3.032 27.3255 3.212 ;
      RECT MASK 1 27.7235 3.032 27.7835 3.212 ;
      RECT MASK 1 28.1815 3.032 28.2415 3.212 ;
      RECT MASK 1 28.6395 3.032 28.6995 3.212 ;
      RECT MASK 1 29.0975 3.032 29.1575 3.212 ;
      RECT MASK 1 29.5555 3.032 29.6155 3.212 ;
      RECT MASK 1 30.0135 3.032 30.0735 3.212 ;
      RECT MASK 1 30.4715 3.032 30.5315 3.212 ;
      RECT MASK 1 30.9295 3.032 30.9895 3.212 ;
      RECT MASK 1 31.3875 3.032 31.4475 3.212 ;
      RECT MASK 1 31.8455 3.032 31.9055 3.212 ;
      RECT MASK 1 32.3035 3.032 32.3635 3.212 ;
      RECT MASK 1 34.1575 3.032 34.2175 3.212 ;
      RECT MASK 1 34.6155 3.032 34.6755 3.212 ;
      RECT MASK 1 35.0735 3.032 35.1335 3.212 ;
      RECT MASK 1 35.5315 3.032 35.5915 3.212 ;
      RECT MASK 1 37.1455 3.032 37.2055 3.212 ;
      RECT MASK 1 37.3745 3.032 37.4345 3.212 ;
      RECT MASK 1 37.6035 3.032 37.6635 3.212 ;
      RECT MASK 1 37.8325 3.032 37.8925 3.212 ;
      RECT MASK 1 38.0615 3.032 38.1215 3.212 ;
      RECT MASK 1 38.5195 3.032 38.5795 3.212 ;
      RECT MASK 1 38.9775 3.032 39.0375 3.212 ;
      RECT MASK 1 39.4355 3.032 39.4955 3.212 ;
      RECT MASK 1 39.8935 3.032 39.9535 3.212 ;
      RECT MASK 1 40.3515 3.032 40.4115 3.212 ;
      RECT MASK 1 40.8095 3.032 40.8695 3.212 ;
      RECT MASK 1 41.2675 3.032 41.3275 3.212 ;
      RECT MASK 1 41.7255 3.032 41.7855 3.212 ;
      RECT MASK 1 41.9545 3.032 42.0145 3.212 ;
      RECT MASK 1 42.1835 3.032 42.2435 3.212 ;
      RECT MASK 1 42.4125 3.032 42.4725 3.212 ;
      RECT MASK 1 42.6415 3.032 42.7015 3.212 ;
      RECT MASK 1 42.8705 3.032 42.9305 3.212 ;
      RECT MASK 1 43.0995 3.032 43.1595 3.212 ;
      RECT MASK 1 43.3285 3.032 43.3885 3.212 ;
      RECT MASK 1 43.5575 3.032 43.6175 3.212 ;
      RECT MASK 1 44.0155 3.032 44.0755 3.212 ;
      RECT MASK 1 44.4735 3.032 44.5335 3.212 ;
      RECT MASK 1 22.2135 3.048 23.3235 3.072 ;
      RECT MASK 1 23.6135 3.048 24.7235 3.072 ;
      RECT MASK 1 62.633 3.078 63.0765 3.118 ;
      RECT MASK 1 63.6735 3.078 65.3665 3.118 ;
      RECT MASK 1 65.5055 3.078 65.949 3.118 ;
      RECT MASK 1 46.6605 3.08 49.2605 3.1 ;
      RECT MASK 1 22.2135 3.138 23.3235 3.162 ;
      RECT MASK 1 23.6135 3.138 24.7235 3.162 ;
      RECT MASK 1 46.6605 3.16 49.2605 3.18 ;
      RECT MASK 1 46.6605 3.24 49.2605 3.26 ;
      RECT MASK 1 46.6605 3.32 49.2605 3.34 ;
      RECT MASK 1 62.633 3.482 63.0765 3.522 ;
      RECT MASK 1 63.549 3.482 64.2215 3.522 ;
      RECT MASK 1 64.465 3.482 65.8245 3.522 ;
      RECT MASK 1 57.789 3.5425 57.969 3.5825 ;
      RECT MASK 1 60.995 3.5425 61.404 3.5825 ;
      RECT MASK 1 61.911 3.5425 62.091 3.5825 ;
      RECT MASK 1 46.6605 3.56 49.2605 3.58 ;
      RECT MASK 1 50.0675 3.57 50.2475 3.63 ;
      RECT MASK 1 50.3895 3.57 50.5695 3.63 ;
      RECT MASK 1 50.7315 3.57 50.9115 3.63 ;
      RECT MASK 1 51.0535 3.57 51.2335 3.63 ;
      RECT MASK 1 51.3955 3.57 51.5755 3.63 ;
      RECT MASK 1 51.7175 3.57 51.8975 3.63 ;
      RECT MASK 1 52.0595 3.57 52.2395 3.63 ;
      RECT MASK 1 52.3815 3.57 52.5615 3.63 ;
      RECT MASK 1 116.154 3.6 116.214 4.65 ;
      RECT MASK 1 116.428 3.6 116.488 4.65 ;
      RECT MASK 1 116.702 3.6 116.762 4.65 ;
      RECT MASK 1 116.976 3.6 117.036 4.65 ;
      RECT MASK 1 117.25 3.6 117.31 4.65 ;
      RECT MASK 1 117.524 3.6 117.584 4.65 ;
      RECT MASK 1 117.798 3.6 117.858 4.65 ;
      RECT MASK 1 118.072 3.6 118.132 4.65 ;
      RECT MASK 1 118.346 3.6 118.406 4.65 ;
      RECT MASK 1 118.62 3.6 118.68 4.65 ;
      RECT MASK 1 118.894 3.6 118.954 4.65 ;
      RECT MASK 1 119.168 3.6 119.228 4.65 ;
      RECT MASK 1 119.442 3.6 119.502 4.65 ;
      RECT MASK 1 119.716 3.6 119.776 4.65 ;
      RECT MASK 1 119.99 3.6 120.05 4.65 ;
      RECT MASK 1 120.264 3.6 120.324 4.65 ;
      RECT MASK 1 120.538 3.6 120.598 4.65 ;
      RECT MASK 1 120.812 3.6 120.872 4.65 ;
      RECT MASK 1 121.086 3.6 121.146 4.65 ;
      RECT MASK 1 121.36 3.6 121.42 4.65 ;
      RECT MASK 1 121.634 3.6 121.694 4.65 ;
      RECT MASK 1 121.908 3.6 121.968 4.65 ;
      RECT MASK 1 122.182 3.6 122.242 4.65 ;
      RECT MASK 1 122.456 3.6 122.516 4.65 ;
      RECT MASK 1 122.73 3.6 122.79 4.65 ;
      RECT MASK 1 123.004 3.6 123.064 4.65 ;
      RECT MASK 1 123.278 3.6 123.338 4.65 ;
      RECT MASK 1 123.552 3.6 123.612 4.65 ;
      RECT MASK 1 123.826 3.6 123.886 4.65 ;
      RECT MASK 1 124.1 3.6 124.16 4.65 ;
      RECT MASK 1 124.374 3.6 124.434 4.65 ;
      RECT MASK 1 124.648 3.6 124.708 4.65 ;
      RECT MASK 1 124.922 3.6 124.982 4.65 ;
      RECT MASK 1 125.196 3.6 125.256 4.65 ;
      RECT MASK 1 125.47 3.6 125.53 4.65 ;
      RECT MASK 1 125.744 3.6 125.804 4.65 ;
      RECT MASK 1 126.018 3.6 126.078 4.65 ;
      RECT MASK 1 126.292 3.6 126.352 4.65 ;
      RECT MASK 1 126.566 3.6 126.626 4.65 ;
      RECT MASK 1 126.84 3.6 126.9 4.65 ;
      RECT MASK 1 127.114 3.6 127.174 4.65 ;
      RECT MASK 1 127.388 3.6 127.448 4.65 ;
      RECT MASK 1 127.662 3.6 127.722 4.65 ;
      RECT MASK 1 127.936 3.6 127.996 4.65 ;
      RECT MASK 1 128.21 3.6 128.27 4.65 ;
      RECT MASK 1 46.6605 3.64 49.2605 3.66 ;
      RECT MASK 1 72.7245 3.64 76.9845 3.68 ;
      RECT MASK 1 77.4385 3.64 82.3625 3.68 ;
      RECT MASK 1 104.3425 3.64 109.2665 3.68 ;
      RECT MASK 1 109.7205 3.64 113.9805 3.68 ;
      RECT MASK 1 58.536 3.662 58.596 3.842 ;
      RECT MASK 1 58.994 3.662 59.054 3.842 ;
      RECT MASK 1 59.452 3.662 59.512 3.842 ;
      RECT MASK 1 59.91 3.662 59.97 3.842 ;
      RECT MASK 1 60.368 3.662 60.428 3.842 ;
      RECT MASK 1 62.887 3.662 62.947 3.842 ;
      RECT MASK 1 63.345 3.662 63.405 3.842 ;
      RECT MASK 1 63.803 3.662 63.863 3.842 ;
      RECT MASK 1 64.261 3.662 64.321 3.842 ;
      RECT MASK 1 64.719 3.662 64.779 3.842 ;
      RECT MASK 1 65.177 3.662 65.237 3.842 ;
      RECT MASK 1 65.635 3.662 65.695 3.842 ;
      RECT MASK 1 1.6805 3.67 13.9525 3.71 ;
      RECT MASK 1 14.3195 3.67 21.7575 3.71 ;
      RECT MASK 1 25.1795 3.67 32.6175 3.71 ;
      RECT MASK 1 32.9845 3.67 45.2565 3.71 ;
      RECT MASK 1 46.6605 3.72 49.2605 3.74 ;
      RECT MASK 1 46.6605 3.8 49.2605 3.82 ;
      RECT MASK 1 50.0675 3.81 50.2475 3.87 ;
      RECT MASK 1 50.3895 3.81 50.5695 3.87 ;
      RECT MASK 1 50.7315 3.81 50.9115 3.87 ;
      RECT MASK 1 51.0535 3.81 51.2335 3.87 ;
      RECT MASK 1 51.3955 3.81 51.5755 3.87 ;
      RECT MASK 1 51.7175 3.81 51.8975 3.87 ;
      RECT MASK 1 52.0595 3.81 52.2395 3.87 ;
      RECT MASK 1 52.3815 3.81 52.5615 3.87 ;
      RECT MASK 1 46.6605 3.88 49.2605 3.9 ;
      RECT MASK 1 83.7885 3.88 93.0585 3.92 ;
      RECT MASK 1 93.6465 3.88 102.9165 3.92 ;
      RECT MASK 1 72.7395 3.9335 72.8195 8.4265 ;
      RECT MASK 1 76.8895 3.9335 76.9695 8.4265 ;
      RECT MASK 1 77.4535 3.9335 77.5335 10.1365 ;
      RECT MASK 1 82.2675 3.9335 82.3475 10.1365 ;
      RECT MASK 1 104.3575 3.9335 104.4375 10.1365 ;
      RECT MASK 1 109.1715 3.9335 109.2515 10.1365 ;
      RECT MASK 1 109.7355 3.9335 109.8155 8.4265 ;
      RECT MASK 1 113.8855 3.9335 113.9655 8.4265 ;
      RECT MASK 1 62.5395 3.9595 62.743 3.9875 ;
      RECT MASK 1 65.839 3.9595 66.042 3.9875 ;
      RECT MASK 1 46.6605 3.96 49.2605 3.98 ;
      RECT MASK 1 46.6605 4.04 49.2605 4.06 ;
      RECT MASK 1 49.8465 4.08 50.0265 4.14 ;
      RECT MASK 1 50.3565 4.08 50.6125 4.14 ;
      RECT MASK 1 51.0205 4.08 51.2765 4.14 ;
      RECT MASK 1 51.6845 4.08 51.9405 4.14 ;
      RECT MASK 1 52.3485 4.08 52.6045 4.14 ;
      RECT MASK 1 83.8035 4.11 83.8835 6.21 ;
      RECT MASK 1 92.9635 4.11 93.0435 6.21 ;
      RECT MASK 1 93.6615 4.11 93.7415 6.21 ;
      RECT MASK 1 102.8215 4.11 102.9015 6.21 ;
      RECT MASK 1 2.4035 4.168 2.4635 4.348 ;
      RECT MASK 1 2.8615 4.168 2.9215 4.348 ;
      RECT MASK 1 3.3195 4.168 3.3795 4.348 ;
      RECT MASK 1 3.5485 4.168 3.6085 4.348 ;
      RECT MASK 1 3.7775 4.168 3.8375 4.348 ;
      RECT MASK 1 4.0065 4.168 4.0665 4.348 ;
      RECT MASK 1 4.2355 4.168 4.2955 4.348 ;
      RECT MASK 1 4.4645 4.168 4.5245 4.348 ;
      RECT MASK 1 4.6935 4.168 4.7535 4.348 ;
      RECT MASK 1 4.9225 4.168 4.9825 4.348 ;
      RECT MASK 1 5.1515 4.168 5.2115 4.348 ;
      RECT MASK 1 5.6095 4.168 5.6695 4.348 ;
      RECT MASK 1 6.0675 4.168 6.1275 4.348 ;
      RECT MASK 1 6.5255 4.168 6.5855 4.348 ;
      RECT MASK 1 6.9835 4.168 7.0435 4.348 ;
      RECT MASK 1 7.4415 4.168 7.5015 4.348 ;
      RECT MASK 1 7.8995 4.168 7.9595 4.348 ;
      RECT MASK 1 8.3575 4.168 8.4175 4.348 ;
      RECT MASK 1 8.8155 4.168 8.8755 4.348 ;
      RECT MASK 1 9.0445 4.168 9.1045 4.348 ;
      RECT MASK 1 9.2735 4.168 9.3335 4.348 ;
      RECT MASK 1 9.5025 4.168 9.5625 4.348 ;
      RECT MASK 1 9.7315 4.168 9.7915 4.348 ;
      RECT MASK 1 11.3455 4.168 11.4055 4.348 ;
      RECT MASK 1 11.8035 4.168 11.8635 4.348 ;
      RECT MASK 1 12.2615 4.168 12.3215 4.348 ;
      RECT MASK 1 12.7195 4.168 12.7795 4.348 ;
      RECT MASK 1 14.5735 4.168 14.6335 4.348 ;
      RECT MASK 1 15.0315 4.168 15.0915 4.348 ;
      RECT MASK 1 15.4895 4.168 15.5495 4.348 ;
      RECT MASK 1 15.9475 4.168 16.0075 4.348 ;
      RECT MASK 1 16.4055 4.168 16.4655 4.348 ;
      RECT MASK 1 16.8635 4.168 16.9235 4.348 ;
      RECT MASK 1 17.3215 4.168 17.3815 4.348 ;
      RECT MASK 1 17.7795 4.168 17.8395 4.348 ;
      RECT MASK 1 18.2375 4.168 18.2975 4.348 ;
      RECT MASK 1 18.6955 4.168 18.7555 4.348 ;
      RECT MASK 1 19.1535 4.168 19.2135 4.348 ;
      RECT MASK 1 19.6115 4.168 19.6715 4.348 ;
      RECT MASK 1 20.0695 4.168 20.1295 4.348 ;
      RECT MASK 1 20.5275 4.168 20.5875 4.348 ;
      RECT MASK 1 20.9855 4.168 21.0455 4.348 ;
      RECT MASK 1 21.4435 4.168 21.5035 4.348 ;
      RECT MASK 1 25.4335 4.168 25.4935 4.348 ;
      RECT MASK 1 25.8915 4.168 25.9515 4.348 ;
      RECT MASK 1 26.3495 4.168 26.4095 4.348 ;
      RECT MASK 1 26.8075 4.168 26.8675 4.348 ;
      RECT MASK 1 27.2655 4.168 27.3255 4.348 ;
      RECT MASK 1 27.7235 4.168 27.7835 4.348 ;
      RECT MASK 1 28.1815 4.168 28.2415 4.348 ;
      RECT MASK 1 28.6395 4.168 28.6995 4.348 ;
      RECT MASK 1 29.0975 4.168 29.1575 4.348 ;
      RECT MASK 1 29.5555 4.168 29.6155 4.348 ;
      RECT MASK 1 30.0135 4.168 30.0735 4.348 ;
      RECT MASK 1 30.4715 4.168 30.5315 4.348 ;
      RECT MASK 1 30.9295 4.168 30.9895 4.348 ;
      RECT MASK 1 31.3875 4.168 31.4475 4.348 ;
      RECT MASK 1 31.8455 4.168 31.9055 4.348 ;
      RECT MASK 1 32.3035 4.168 32.3635 4.348 ;
      RECT MASK 1 34.1575 4.168 34.2175 4.348 ;
      RECT MASK 1 34.6155 4.168 34.6755 4.348 ;
      RECT MASK 1 35.0735 4.168 35.1335 4.348 ;
      RECT MASK 1 35.5315 4.168 35.5915 4.348 ;
      RECT MASK 1 37.1455 4.168 37.2055 4.348 ;
      RECT MASK 1 37.3745 4.168 37.4345 4.348 ;
      RECT MASK 1 37.6035 4.168 37.6635 4.348 ;
      RECT MASK 1 37.8325 4.168 37.8925 4.348 ;
      RECT MASK 1 38.0615 4.168 38.1215 4.348 ;
      RECT MASK 1 38.5195 4.168 38.5795 4.348 ;
      RECT MASK 1 38.9775 4.168 39.0375 4.348 ;
      RECT MASK 1 39.4355 4.168 39.4955 4.348 ;
      RECT MASK 1 39.8935 4.168 39.9535 4.348 ;
      RECT MASK 1 40.3515 4.168 40.4115 4.348 ;
      RECT MASK 1 40.8095 4.168 40.8695 4.348 ;
      RECT MASK 1 41.2675 4.168 41.3275 4.348 ;
      RECT MASK 1 41.7255 4.168 41.7855 4.348 ;
      RECT MASK 1 41.9545 4.168 42.0145 4.348 ;
      RECT MASK 1 42.1835 4.168 42.2435 4.348 ;
      RECT MASK 1 42.4125 4.168 42.4725 4.348 ;
      RECT MASK 1 42.6415 4.168 42.7015 4.348 ;
      RECT MASK 1 42.8705 4.168 42.9305 4.348 ;
      RECT MASK 1 43.0995 4.168 43.1595 4.348 ;
      RECT MASK 1 43.3285 4.168 43.3885 4.348 ;
      RECT MASK 1 43.5575 4.168 43.6175 4.348 ;
      RECT MASK 1 44.0155 4.168 44.0755 4.348 ;
      RECT MASK 1 44.4735 4.168 44.5335 4.348 ;
      RECT MASK 1 62.5395 4.1725 62.743 4.2005 ;
      RECT MASK 1 65.839 4.1725 66.042 4.2005 ;
      RECT MASK 1 22.2135 4.218 23.3235 4.242 ;
      RECT MASK 1 23.6135 4.218 24.7235 4.242 ;
      RECT MASK 1 22.2135 4.308 23.3235 4.332 ;
      RECT MASK 1 23.6135 4.308 24.7235 4.332 ;
      RECT MASK 1 58.536 4.318 58.596 4.498 ;
      RECT MASK 1 58.994 4.318 59.054 4.498 ;
      RECT MASK 1 59.452 4.318 59.512 4.498 ;
      RECT MASK 1 59.91 4.318 59.97 4.498 ;
      RECT MASK 1 60.368 4.318 60.428 4.498 ;
      RECT MASK 1 62.887 4.318 62.947 4.498 ;
      RECT MASK 1 63.345 4.318 63.405 4.498 ;
      RECT MASK 1 63.803 4.318 63.863 4.498 ;
      RECT MASK 1 64.261 4.318 64.321 4.498 ;
      RECT MASK 1 64.719 4.318 64.779 4.498 ;
      RECT MASK 1 65.177 4.318 65.237 4.498 ;
      RECT MASK 1 65.635 4.318 65.695 4.498 ;
      RECT MASK 1 22.2135 4.398 23.3235 4.422 ;
      RECT MASK 1 23.6135 4.398 24.7235 4.422 ;
      RECT MASK 1 10.107 4.4275 10.7505 4.4675 ;
      RECT MASK 1 13.5865 4.4275 13.7665 4.4675 ;
      RECT MASK 1 33.1705 4.4275 33.3505 4.4675 ;
      RECT MASK 1 36.3985 4.4275 36.5785 4.4675 ;
      RECT MASK 1 1.6135 4.4875 1.8575 4.5275 ;
      RECT MASK 1 45.0795 4.4875 45.3235 4.5275 ;
      RECT MASK 1 49.8465 4.5 50.0265 4.56 ;
      RECT MASK 1 50.3565 4.5 50.6125 4.56 ;
      RECT MASK 1 51.0205 4.5 51.2765 4.56 ;
      RECT MASK 1 51.6845 4.5 51.9405 4.56 ;
      RECT MASK 1 52.3485 4.5 52.6045 4.56 ;
      RECT MASK 1 57.789 4.5775 57.969 4.6175 ;
      RECT MASK 1 60.995 4.5775 61.404 4.6175 ;
      RECT MASK 1 61.911 4.5775 62.091 4.6175 ;
      RECT MASK 1 2.5025 4.589 2.7175 4.629 ;
      RECT MASK 1 3.5235 4.589 9.692 4.629 ;
      RECT MASK 1 10.9455 4.589 11.764 4.629 ;
      RECT MASK 1 14.663 4.589 21.414 4.629 ;
      RECT MASK 1 25.523 4.589 32.274 4.629 ;
      RECT MASK 1 35.173 4.589 35.9915 4.629 ;
      RECT MASK 1 37.245 4.589 43.4135 4.629 ;
      RECT MASK 1 44.2195 4.589 44.4345 4.629 ;
      RECT MASK 1 84.7145 4.619 86.3915 4.679 ;
      RECT MASK 1 86.5465 4.619 90.3005 4.679 ;
      RECT MASK 1 90.6685 4.619 92.1325 4.679 ;
      RECT MASK 1 94.5725 4.619 96.0365 4.679 ;
      RECT MASK 1 96.4045 4.619 100.1585 4.679 ;
      RECT MASK 1 100.3135 4.619 101.9905 4.679 ;
      RECT MASK 1 62.633 4.638 63.0765 4.678 ;
      RECT MASK 1 63.549 4.638 64.2215 4.678 ;
      RECT MASK 1 64.465 4.638 65.8245 4.678 ;
      RECT MASK 1 22.7735 4.758 23.1635 4.782 ;
      RECT MASK 1 23.7135 4.758 24.1635 4.782 ;
      RECT MASK 1 50.0675 4.77 50.2475 4.83 ;
      RECT MASK 1 50.3895 4.77 50.5695 4.83 ;
      RECT MASK 1 50.7315 4.77 50.9115 4.83 ;
      RECT MASK 1 51.0535 4.77 51.2335 4.83 ;
      RECT MASK 1 51.3955 4.77 51.5755 4.83 ;
      RECT MASK 1 51.7175 4.77 51.8975 4.83 ;
      RECT MASK 1 52.0595 4.77 52.2395 4.83 ;
      RECT MASK 1 52.3815 4.77 52.5615 4.83 ;
      RECT MASK 1 2.5025 4.791 2.7175 4.831 ;
      RECT MASK 1 2.8365 4.791 4.196 4.831 ;
      RECT MASK 1 5.7055 4.791 8.57 4.831 ;
      RECT MASK 1 9.373 4.791 10.0665 4.831 ;
      RECT MASK 1 11.0705 4.791 11.764 4.831 ;
      RECT MASK 1 12.361 4.791 13.0765 4.831 ;
      RECT MASK 1 14.663 4.791 21.414 4.831 ;
      RECT MASK 1 25.523 4.791 32.274 4.831 ;
      RECT MASK 1 33.8605 4.791 34.576 4.831 ;
      RECT MASK 1 35.173 4.791 35.8665 4.831 ;
      RECT MASK 1 36.8705 4.791 37.564 4.831 ;
      RECT MASK 1 38.367 4.791 41.2315 4.831 ;
      RECT MASK 1 42.741 4.791 44.1005 4.831 ;
      RECT MASK 1 44.2195 4.791 44.4345 4.831 ;
      RECT MASK 1 22.2135 4.848 23.3235 4.872 ;
      RECT MASK 1 23.6135 4.848 24.7235 4.872 ;
      RECT MASK 1 1.6135 4.8925 1.8575 4.9325 ;
      RECT MASK 1 45.0795 4.8925 45.3235 4.9325 ;
      RECT MASK 1 22.4135 4.938 22.7135 4.962 ;
      RECT MASK 1 22.8235 4.938 23.1235 4.962 ;
      RECT MASK 1 23.8135 4.938 24.1135 4.962 ;
      RECT MASK 1 24.2235 4.938 24.5235 4.962 ;
      RECT MASK 1 10.3585 4.9525 10.5385 4.9925 ;
      RECT MASK 1 13.5865 4.9525 13.7665 4.9925 ;
      RECT MASK 1 33.1705 4.9525 33.3505 4.9925 ;
      RECT MASK 1 36.3985 4.9525 36.5785 4.9925 ;
      RECT MASK 1 50.0675 5.01 50.2475 5.07 ;
      RECT MASK 1 50.3895 5.01 50.5695 5.07 ;
      RECT MASK 1 50.7315 5.01 50.9115 5.07 ;
      RECT MASK 1 51.0535 5.01 51.2335 5.07 ;
      RECT MASK 1 51.3955 5.01 51.5755 5.07 ;
      RECT MASK 1 51.7175 5.01 51.8975 5.07 ;
      RECT MASK 1 52.0595 5.01 52.2395 5.07 ;
      RECT MASK 1 52.3815 5.01 52.5615 5.07 ;
      RECT MASK 1 22.4135 5.028 22.7135 5.052 ;
      RECT MASK 1 22.8235 5.028 23.1235 5.052 ;
      RECT MASK 1 23.8135 5.028 24.1135 5.052 ;
      RECT MASK 1 24.2235 5.028 24.5235 5.052 ;
      RECT MASK 1 62.633 5.042 63.0765 5.082 ;
      RECT MASK 1 63.6735 5.042 65.3665 5.082 ;
      RECT MASK 1 65.5055 5.042 65.949 5.082 ;
      RECT MASK 1 2.8615 5.071 2.9215 5.252 ;
      RECT MASK 1 5.1515 5.071 5.2115 5.252 ;
      RECT MASK 1 41.7255 5.071 41.7855 5.252 ;
      RECT MASK 1 44.0155 5.071 44.0755 5.252 ;
      RECT MASK 1 2.4035 5.072 2.4635 5.252 ;
      RECT MASK 1 3.3195 5.072 3.3795 5.252 ;
      RECT MASK 1 3.5485 5.072 3.6085 5.252 ;
      RECT MASK 1 3.7775 5.072 3.8375 5.252 ;
      RECT MASK 1 4.0065 5.072 4.0665 5.252 ;
      RECT MASK 1 4.2355 5.072 4.2955 5.252 ;
      RECT MASK 1 4.4645 5.072 4.5245 5.252 ;
      RECT MASK 1 4.6935 5.072 4.7535 5.252 ;
      RECT MASK 1 4.9225 5.072 4.9825 5.252 ;
      RECT MASK 1 5.6095 5.072 5.6695 5.252 ;
      RECT MASK 1 6.0675 5.072 6.1275 5.252 ;
      RECT MASK 1 6.5255 5.072 6.5855 5.252 ;
      RECT MASK 1 6.9835 5.072 7.0435 5.252 ;
      RECT MASK 1 7.4415 5.072 7.5015 5.252 ;
      RECT MASK 1 7.8995 5.072 7.9595 5.252 ;
      RECT MASK 1 8.3575 5.072 8.4175 5.252 ;
      RECT MASK 1 8.8155 5.072 8.8755 5.252 ;
      RECT MASK 1 9.0445 5.072 9.1045 5.252 ;
      RECT MASK 1 9.2735 5.072 9.3335 5.252 ;
      RECT MASK 1 9.5025 5.072 9.5625 5.252 ;
      RECT MASK 1 9.7315 5.072 9.7915 5.252 ;
      RECT MASK 1 11.3455 5.072 11.4055 5.252 ;
      RECT MASK 1 11.8035 5.072 11.8635 5.252 ;
      RECT MASK 1 12.2615 5.072 12.3215 5.252 ;
      RECT MASK 1 12.7195 5.072 12.7795 5.252 ;
      RECT MASK 1 14.5735 5.072 14.6335 5.252 ;
      RECT MASK 1 15.0315 5.072 15.0915 5.252 ;
      RECT MASK 1 15.4895 5.072 15.5495 5.252 ;
      RECT MASK 1 15.9475 5.072 16.0075 5.252 ;
      RECT MASK 1 16.4055 5.072 16.4655 5.252 ;
      RECT MASK 1 16.8635 5.072 16.9235 5.252 ;
      RECT MASK 1 17.3215 5.072 17.3815 5.252 ;
      RECT MASK 1 17.7795 5.072 17.8395 5.252 ;
      RECT MASK 1 18.2375 5.072 18.2975 5.252 ;
      RECT MASK 1 18.6955 5.072 18.7555 5.252 ;
      RECT MASK 1 19.1535 5.072 19.2135 5.252 ;
      RECT MASK 1 19.6115 5.072 19.6715 5.252 ;
      RECT MASK 1 20.0695 5.072 20.1295 5.252 ;
      RECT MASK 1 20.5275 5.072 20.5875 5.252 ;
      RECT MASK 1 20.9855 5.072 21.0455 5.252 ;
      RECT MASK 1 21.4435 5.072 21.5035 5.252 ;
      RECT MASK 1 25.4335 5.072 25.4935 5.252 ;
      RECT MASK 1 25.8915 5.072 25.9515 5.252 ;
      RECT MASK 1 26.3495 5.072 26.4095 5.252 ;
      RECT MASK 1 26.8075 5.072 26.8675 5.252 ;
      RECT MASK 1 27.2655 5.072 27.3255 5.252 ;
      RECT MASK 1 27.7235 5.072 27.7835 5.252 ;
      RECT MASK 1 28.1815 5.072 28.2415 5.252 ;
      RECT MASK 1 28.6395 5.072 28.6995 5.252 ;
      RECT MASK 1 29.0975 5.072 29.1575 5.252 ;
      RECT MASK 1 29.5555 5.072 29.6155 5.252 ;
      RECT MASK 1 30.0135 5.072 30.0735 5.252 ;
      RECT MASK 1 30.4715 5.072 30.5315 5.252 ;
      RECT MASK 1 30.9295 5.072 30.9895 5.252 ;
      RECT MASK 1 31.3875 5.072 31.4475 5.252 ;
      RECT MASK 1 31.8455 5.072 31.9055 5.252 ;
      RECT MASK 1 32.3035 5.072 32.3635 5.252 ;
      RECT MASK 1 34.1575 5.072 34.2175 5.252 ;
      RECT MASK 1 34.6155 5.072 34.6755 5.252 ;
      RECT MASK 1 35.0735 5.072 35.1335 5.252 ;
      RECT MASK 1 35.5315 5.072 35.5915 5.252 ;
      RECT MASK 1 37.1455 5.072 37.2055 5.252 ;
      RECT MASK 1 37.3745 5.072 37.4345 5.252 ;
      RECT MASK 1 37.6035 5.072 37.6635 5.252 ;
      RECT MASK 1 37.8325 5.072 37.8925 5.252 ;
      RECT MASK 1 38.0615 5.072 38.1215 5.252 ;
      RECT MASK 1 38.5195 5.072 38.5795 5.252 ;
      RECT MASK 1 38.9775 5.072 39.0375 5.252 ;
      RECT MASK 1 39.4355 5.072 39.4955 5.252 ;
      RECT MASK 1 39.8935 5.072 39.9535 5.252 ;
      RECT MASK 1 40.3515 5.072 40.4115 5.252 ;
      RECT MASK 1 40.8095 5.072 40.8695 5.252 ;
      RECT MASK 1 41.2675 5.072 41.3275 5.252 ;
      RECT MASK 1 41.9545 5.072 42.0145 5.252 ;
      RECT MASK 1 42.1835 5.072 42.2435 5.252 ;
      RECT MASK 1 42.4125 5.072 42.4725 5.252 ;
      RECT MASK 1 42.6415 5.072 42.7015 5.252 ;
      RECT MASK 1 42.8705 5.072 42.9305 5.252 ;
      RECT MASK 1 43.0995 5.072 43.1595 5.252 ;
      RECT MASK 1 43.3285 5.072 43.3885 5.252 ;
      RECT MASK 1 43.5575 5.072 43.6175 5.252 ;
      RECT MASK 1 44.4735 5.072 44.5335 5.252 ;
      RECT MASK 1 84.4855 5.098 88.2395 5.158 ;
      RECT MASK 1 88.6075 5.098 92.3615 5.158 ;
      RECT MASK 1 94.3435 5.098 98.0975 5.158 ;
      RECT MASK 1 98.4655 5.098 102.2195 5.158 ;
      RECT MASK 1 57.789 5.1025 57.969 5.1425 ;
      RECT MASK 1 22.4135 5.118 22.7135 5.142 ;
      RECT MASK 1 22.8235 5.118 23.1235 5.142 ;
      RECT MASK 1 23.8135 5.118 24.1135 5.142 ;
      RECT MASK 1 24.2235 5.118 24.5235 5.142 ;
      RECT MASK 1 58.536 5.222 58.596 5.402 ;
      RECT MASK 1 58.994 5.222 59.054 5.402 ;
      RECT MASK 1 59.452 5.222 59.512 5.402 ;
      RECT MASK 1 59.91 5.222 59.97 5.402 ;
      RECT MASK 1 60.368 5.222 60.428 5.402 ;
      RECT MASK 1 62.887 5.222 62.947 5.402 ;
      RECT MASK 1 63.345 5.222 63.405 5.402 ;
      RECT MASK 1 63.803 5.222 63.863 5.402 ;
      RECT MASK 1 64.261 5.222 64.321 5.402 ;
      RECT MASK 1 64.719 5.222 64.779 5.402 ;
      RECT MASK 1 65.177 5.222 65.237 5.402 ;
      RECT MASK 1 65.635 5.222 65.695 5.402 ;
      RECT MASK 1 60.995 5.2225 61.404 5.2625 ;
      RECT MASK 1 61.911 5.2225 62.091 5.2625 ;
      RECT MASK 1 46.8655 5.23 48.9595 5.27 ;
      RECT MASK 1 116.154 5.31 116.214 6.36 ;
      RECT MASK 1 116.428 5.31 116.488 6.36 ;
      RECT MASK 1 116.702 5.31 116.762 6.36 ;
      RECT MASK 1 116.976 5.31 117.036 6.36 ;
      RECT MASK 1 117.25 5.31 117.31 6.36 ;
      RECT MASK 1 117.524 5.31 117.584 6.36 ;
      RECT MASK 1 117.798 5.31 117.858 6.36 ;
      RECT MASK 1 118.072 5.31 118.132 6.36 ;
      RECT MASK 1 118.346 5.31 118.406 6.36 ;
      RECT MASK 1 118.62 5.31 118.68 6.36 ;
      RECT MASK 1 118.894 5.31 118.954 6.36 ;
      RECT MASK 1 119.168 5.31 119.228 6.36 ;
      RECT MASK 1 119.442 5.31 119.502 6.36 ;
      RECT MASK 1 119.716 5.31 119.776 6.36 ;
      RECT MASK 1 119.99 5.31 120.05 6.36 ;
      RECT MASK 1 120.264 5.31 120.324 6.36 ;
      RECT MASK 1 120.538 5.31 120.598 6.36 ;
      RECT MASK 1 120.812 5.31 120.872 6.36 ;
      RECT MASK 1 121.086 5.31 121.146 6.36 ;
      RECT MASK 1 121.36 5.31 121.42 6.36 ;
      RECT MASK 1 121.634 5.31 121.694 6.36 ;
      RECT MASK 1 121.908 5.31 121.968 6.36 ;
      RECT MASK 1 122.182 5.31 122.242 6.36 ;
      RECT MASK 1 122.456 5.31 122.516 6.36 ;
      RECT MASK 1 122.73 5.31 122.79 6.36 ;
      RECT MASK 1 123.004 5.31 123.064 6.36 ;
      RECT MASK 1 123.278 5.31 123.338 6.36 ;
      RECT MASK 1 123.552 5.31 123.612 6.36 ;
      RECT MASK 1 123.826 5.31 123.886 6.36 ;
      RECT MASK 1 124.1 5.31 124.16 6.36 ;
      RECT MASK 1 124.374 5.31 124.434 6.36 ;
      RECT MASK 1 124.648 5.31 124.708 6.36 ;
      RECT MASK 1 124.922 5.31 124.982 6.36 ;
      RECT MASK 1 125.196 5.31 125.256 6.36 ;
      RECT MASK 1 125.47 5.31 125.53 6.36 ;
      RECT MASK 1 125.744 5.31 125.804 6.36 ;
      RECT MASK 1 126.018 5.31 126.078 6.36 ;
      RECT MASK 1 126.292 5.31 126.352 6.36 ;
      RECT MASK 1 126.566 5.31 126.626 6.36 ;
      RECT MASK 1 126.84 5.31 126.9 6.36 ;
      RECT MASK 1 127.114 5.31 127.174 6.36 ;
      RECT MASK 1 127.388 5.31 127.448 6.36 ;
      RECT MASK 1 127.662 5.31 127.722 6.36 ;
      RECT MASK 1 127.936 5.31 127.996 6.36 ;
      RECT MASK 1 128.21 5.31 128.27 6.36 ;
      RECT MASK 1 84.1235 5.34 84.461 5.4 ;
      RECT MASK 1 84.6 5.34 88.125 5.4 ;
      RECT MASK 1 88.264 5.34 88.583 5.4 ;
      RECT MASK 1 88.722 5.34 92.247 5.4 ;
      RECT MASK 1 92.386 5.34 92.705 5.4 ;
      RECT MASK 1 94 5.34 94.319 5.4 ;
      RECT MASK 1 94.458 5.34 97.983 5.4 ;
      RECT MASK 1 98.122 5.34 98.441 5.4 ;
      RECT MASK 1 98.58 5.34 102.105 5.4 ;
      RECT MASK 1 102.244 5.34 102.5815 5.4 ;
      RECT MASK 1 53.9045 5.35 56.1725 5.39 ;
      RECT MASK 1 22.2235 5.478 23.3235 5.502 ;
      RECT MASK 1 23.6135 5.478 24.7135 5.502 ;
      RECT MASK 1 49.9465 5.49 52.7045 5.55 ;
      RECT MASK 1 62.5395 5.522 62.743 5.55 ;
      RECT MASK 1 65.839 5.522 66.042 5.55 ;
      RECT MASK 1 46.7465 5.551 49.0705 5.591 ;
      RECT MASK 1 53.7935 5.671 56.2835 5.711 ;
      RECT MASK 1 1.6805 5.71 10.7245 5.75 ;
      RECT MASK 1 11.1705 5.71 12.9295 5.75 ;
      RECT MASK 1 13.4005 5.71 21.7575 5.75 ;
      RECT MASK 1 25.1795 5.71 33.5365 5.75 ;
      RECT MASK 1 34.0075 5.71 35.7665 5.75 ;
      RECT MASK 1 36.2125 5.71 45.2565 5.75 ;
      RECT MASK 1 46.7465 5.726 49.0705 5.766 ;
      RECT MASK 1 50.0675 5.73 50.2475 5.79 ;
      RECT MASK 1 50.3895 5.73 50.5695 5.79 ;
      RECT MASK 1 50.7315 5.73 50.9115 5.79 ;
      RECT MASK 1 51.0535 5.73 51.2335 5.79 ;
      RECT MASK 1 51.3955 5.73 51.5755 5.79 ;
      RECT MASK 1 51.7175 5.73 51.8975 5.79 ;
      RECT MASK 1 52.0595 5.73 52.2395 5.79 ;
      RECT MASK 1 52.3815 5.73 52.5615 5.79 ;
      RECT MASK 1 65.0475 5.73 65.949 5.758 ;
      RECT MASK 1 84.4205 5.819 88.2955 5.879 ;
      RECT MASK 1 88.5605 5.819 88.9565 5.879 ;
      RECT MASK 1 89.2645 5.819 89.6485 5.879 ;
      RECT MASK 1 90.1785 5.819 90.4035 5.879 ;
      RECT MASK 1 90.6685 5.819 91.065 5.879 ;
      RECT MASK 1 95.64 5.819 96.0365 5.879 ;
      RECT MASK 1 96.3015 5.819 96.5265 5.879 ;
      RECT MASK 1 97.0565 5.819 97.4405 5.879 ;
      RECT MASK 1 97.7485 5.819 98.1445 5.879 ;
      RECT MASK 1 98.4095 5.819 102.2845 5.879 ;
      RECT MASK 1 53.7935 5.846 56.2835 5.886 ;
      RECT MASK 1 58.765 5.878 58.825 6.058 ;
      RECT MASK 1 59.223 5.878 59.283 6.058 ;
      RECT MASK 1 59.681 5.878 59.741 6.058 ;
      RECT MASK 1 60.826 5.878 60.886 6.058 ;
      RECT MASK 1 61.284 5.878 61.344 6.058 ;
      RECT MASK 1 61.742 5.878 61.802 6.058 ;
      RECT MASK 1 62.2 5.878 62.26 6.058 ;
      RECT MASK 1 62.658 5.878 62.718 6.058 ;
      RECT MASK 1 63.116 5.878 63.176 6.058 ;
      RECT MASK 1 63.803 5.878 63.863 6.058 ;
      RECT MASK 1 64.261 5.878 64.321 6.058 ;
      RECT MASK 1 64.719 5.878 64.779 6.058 ;
      RECT MASK 1 46.9055 5.893 47.1235 5.933 ;
      RECT MASK 1 47.2375 5.893 47.4555 5.933 ;
      RECT MASK 1 22.2235 5.958 23.3235 5.982 ;
      RECT MASK 1 23.6135 5.958 24.7135 5.982 ;
      RECT MASK 1 49.9465 5.97 52.7045 6.03 ;
      RECT MASK 1 48.8145 5.9875 48.9945 6.0275 ;
      RECT MASK 1 54.4505 6.013 54.6685 6.053 ;
      RECT MASK 1 55.2805 6.013 55.4985 6.053 ;
      RECT MASK 1 60.1675 6.0175 60.3475 6.0575 ;
      RECT MASK 1 65.575 6.0175 65.984 6.0575 ;
      RECT MASK 1 47.0715 6.077 47.2515 6.117 ;
      RECT MASK 1 47.4035 6.077 47.5835 6.117 ;
      RECT MASK 1 54.9485 6.096 55.1285 6.136 ;
      RECT MASK 1 53.8695 6.1075 54.0495 6.1475 ;
      RECT MASK 1 56.0275 6.1075 56.2075 6.1475 ;
      RECT MASK 1 57.789 6.1375 57.969 6.1775 ;
      RECT MASK 1 54.6165 6.197 54.7965 6.237 ;
      RECT MASK 1 55.4465 6.197 55.6265 6.237 ;
      RECT MASK 1 61.3835 6.198 62.743 6.238 ;
      RECT MASK 1 2.4035 6.208 2.4635 6.388 ;
      RECT MASK 1 2.8615 6.208 2.9215 6.389 ;
      RECT MASK 1 3.3195 6.208 3.3795 6.388 ;
      RECT MASK 1 3.5485 6.208 3.6085 6.388 ;
      RECT MASK 1 3.7775 6.208 3.8375 6.388 ;
      RECT MASK 1 4.0065 6.208 4.0665 6.388 ;
      RECT MASK 1 4.2355 6.208 4.2955 6.388 ;
      RECT MASK 1 4.4645 6.208 4.5245 6.388 ;
      RECT MASK 1 4.6935 6.208 4.7535 6.388 ;
      RECT MASK 1 4.9225 6.208 4.9825 6.388 ;
      RECT MASK 1 5.1515 6.208 5.2115 6.389 ;
      RECT MASK 1 5.6095 6.208 5.6695 6.388 ;
      RECT MASK 1 6.0675 6.208 6.1275 6.388 ;
      RECT MASK 1 6.5255 6.208 6.5855 6.388 ;
      RECT MASK 1 6.9835 6.208 7.0435 6.388 ;
      RECT MASK 1 7.4415 6.208 7.5015 6.388 ;
      RECT MASK 1 7.8995 6.208 7.9595 6.388 ;
      RECT MASK 1 8.3575 6.208 8.4175 6.388 ;
      RECT MASK 1 8.8155 6.208 8.8755 6.388 ;
      RECT MASK 1 9.0445 6.208 9.1045 6.388 ;
      RECT MASK 1 9.2735 6.208 9.3335 6.388 ;
      RECT MASK 1 9.5025 6.208 9.5625 6.388 ;
      RECT MASK 1 9.7315 6.208 9.7915 6.388 ;
      RECT MASK 1 11.3455 6.208 11.4055 6.388 ;
      RECT MASK 1 11.8035 6.208 11.8635 6.388 ;
      RECT MASK 1 12.2615 6.208 12.3215 6.388 ;
      RECT MASK 1 12.7195 6.208 12.7795 6.388 ;
      RECT MASK 1 14.5735 6.208 14.6335 6.388 ;
      RECT MASK 1 15.0315 6.208 15.0915 6.388 ;
      RECT MASK 1 15.4895 6.208 15.5495 6.388 ;
      RECT MASK 1 15.9475 6.208 16.0075 6.388 ;
      RECT MASK 1 16.4055 6.208 16.4655 6.388 ;
      RECT MASK 1 16.8635 6.208 16.9235 6.388 ;
      RECT MASK 1 17.3215 6.208 17.3815 6.388 ;
      RECT MASK 1 17.7795 6.208 17.8395 6.388 ;
      RECT MASK 1 18.2375 6.208 18.2975 6.388 ;
      RECT MASK 1 18.6955 6.208 18.7555 6.388 ;
      RECT MASK 1 19.1535 6.208 19.2135 6.388 ;
      RECT MASK 1 19.6115 6.208 19.6715 6.388 ;
      RECT MASK 1 20.0695 6.208 20.1295 6.388 ;
      RECT MASK 1 20.5275 6.208 20.5875 6.388 ;
      RECT MASK 1 20.9855 6.208 21.0455 6.388 ;
      RECT MASK 1 21.4435 6.208 21.5035 6.388 ;
      RECT MASK 1 25.4335 6.208 25.4935 6.388 ;
      RECT MASK 1 25.8915 6.208 25.9515 6.388 ;
      RECT MASK 1 26.3495 6.208 26.4095 6.388 ;
      RECT MASK 1 26.8075 6.208 26.8675 6.388 ;
      RECT MASK 1 27.2655 6.208 27.3255 6.388 ;
      RECT MASK 1 27.7235 6.208 27.7835 6.388 ;
      RECT MASK 1 28.1815 6.208 28.2415 6.388 ;
      RECT MASK 1 28.6395 6.208 28.6995 6.388 ;
      RECT MASK 1 29.0975 6.208 29.1575 6.388 ;
      RECT MASK 1 29.5555 6.208 29.6155 6.388 ;
      RECT MASK 1 30.0135 6.208 30.0735 6.388 ;
      RECT MASK 1 30.4715 6.208 30.5315 6.388 ;
      RECT MASK 1 30.9295 6.208 30.9895 6.388 ;
      RECT MASK 1 31.3875 6.208 31.4475 6.388 ;
      RECT MASK 1 31.8455 6.208 31.9055 6.388 ;
      RECT MASK 1 32.3035 6.208 32.3635 6.388 ;
      RECT MASK 1 34.1575 6.208 34.2175 6.388 ;
      RECT MASK 1 34.6155 6.208 34.6755 6.388 ;
      RECT MASK 1 35.0735 6.208 35.1335 6.388 ;
      RECT MASK 1 35.5315 6.208 35.5915 6.388 ;
      RECT MASK 1 37.1455 6.208 37.2055 6.388 ;
      RECT MASK 1 37.3745 6.208 37.4345 6.388 ;
      RECT MASK 1 37.6035 6.208 37.6635 6.388 ;
      RECT MASK 1 37.8325 6.208 37.8925 6.388 ;
      RECT MASK 1 38.0615 6.208 38.1215 6.388 ;
      RECT MASK 1 38.5195 6.208 38.5795 6.388 ;
      RECT MASK 1 38.9775 6.208 39.0375 6.388 ;
      RECT MASK 1 39.4355 6.208 39.4955 6.388 ;
      RECT MASK 1 39.8935 6.208 39.9535 6.388 ;
      RECT MASK 1 40.3515 6.208 40.4115 6.388 ;
      RECT MASK 1 40.8095 6.208 40.8695 6.388 ;
      RECT MASK 1 41.2675 6.208 41.3275 6.388 ;
      RECT MASK 1 41.7255 6.208 41.7855 6.389 ;
      RECT MASK 1 41.9545 6.208 42.0145 6.388 ;
      RECT MASK 1 42.1835 6.208 42.2435 6.388 ;
      RECT MASK 1 42.4125 6.208 42.4725 6.388 ;
      RECT MASK 1 42.6415 6.208 42.7015 6.388 ;
      RECT MASK 1 42.8705 6.208 42.9305 6.388 ;
      RECT MASK 1 43.0995 6.208 43.1595 6.388 ;
      RECT MASK 1 43.3285 6.208 43.3885 6.388 ;
      RECT MASK 1 43.5575 6.208 43.6175 6.388 ;
      RECT MASK 1 44.0155 6.208 44.0755 6.389 ;
      RECT MASK 1 44.4735 6.208 44.5335 6.388 ;
      RECT MASK 1 47.0715 6.303 47.2515 6.343 ;
      RECT MASK 1 47.4035 6.303 47.5835 6.343 ;
      RECT MASK 1 22.4135 6.318 22.7135 6.342 ;
      RECT MASK 1 22.8235 6.318 23.1235 6.342 ;
      RECT MASK 1 23.8135 6.318 24.1135 6.342 ;
      RECT MASK 1 24.2235 6.318 24.5235 6.342 ;
      RECT MASK 1 48.8145 6.3925 48.9945 6.4325 ;
      RECT MASK 1 58.74 6.4 64.804 6.44 ;
      RECT MASK 1 83.7885 6.4 93.0585 6.44 ;
      RECT MASK 1 93.6465 6.4 102.9165 6.44 ;
      RECT MASK 1 22.4135 6.408 22.7135 6.432 ;
      RECT MASK 1 22.8235 6.408 23.1235 6.432 ;
      RECT MASK 1 23.8135 6.408 24.1135 6.432 ;
      RECT MASK 1 24.2235 6.408 24.5235 6.432 ;
      RECT MASK 1 54.6165 6.423 54.7965 6.463 ;
      RECT MASK 1 55.4465 6.423 55.6265 6.463 ;
      RECT MASK 1 49.9395 6.43 52.6895 6.47 ;
      RECT MASK 1 10.3585 6.4675 10.5385 6.5075 ;
      RECT MASK 1 13.5865 6.4675 13.7665 6.5075 ;
      RECT MASK 1 33.1705 6.4675 33.3505 6.5075 ;
      RECT MASK 1 36.3985 6.4675 36.5785 6.5075 ;
      RECT MASK 1 46.9055 6.487 47.1235 6.527 ;
      RECT MASK 1 47.2375 6.487 47.4555 6.527 ;
      RECT MASK 1 22.4135 6.498 22.7135 6.522 ;
      RECT MASK 1 22.8235 6.498 23.1235 6.522 ;
      RECT MASK 1 23.8135 6.498 24.1135 6.522 ;
      RECT MASK 1 24.2235 6.498 24.5235 6.522 ;
      RECT MASK 1 53.8695 6.5125 54.0495 6.5525 ;
      RECT MASK 1 56.0275 6.5125 56.2075 6.5525 ;
      RECT MASK 1 54.9485 6.524 55.1285 6.564 ;
      RECT MASK 1 1.6135 6.5275 1.8575 6.5675 ;
      RECT MASK 1 45.0795 6.5275 45.3235 6.5675 ;
      RECT MASK 1 22.2135 6.588 23.3235 6.612 ;
      RECT MASK 1 23.6135 6.588 24.7235 6.612 ;
      RECT MASK 1 61.259 6.602 62.6185 6.642 ;
      RECT MASK 1 54.4505 6.607 54.6685 6.647 ;
      RECT MASK 1 55.2805 6.607 55.4985 6.647 ;
      RECT MASK 1 2.5025 6.629 2.7175 6.669 ;
      RECT MASK 1 2.8365 6.629 4.196 6.669 ;
      RECT MASK 1 5.7055 6.629 8.57 6.669 ;
      RECT MASK 1 9.373 6.629 10.0665 6.669 ;
      RECT MASK 1 11.0705 6.629 11.764 6.669 ;
      RECT MASK 1 12.361 6.629 13.0765 6.669 ;
      RECT MASK 1 14.663 6.629 21.414 6.669 ;
      RECT MASK 1 25.523 6.629 32.274 6.669 ;
      RECT MASK 1 33.8605 6.629 34.576 6.669 ;
      RECT MASK 1 35.173 6.629 35.8665 6.669 ;
      RECT MASK 1 36.8705 6.629 37.564 6.669 ;
      RECT MASK 1 38.367 6.629 41.2315 6.669 ;
      RECT MASK 1 42.741 6.629 44.1005 6.669 ;
      RECT MASK 1 44.2195 6.629 44.4345 6.669 ;
      RECT MASK 1 46.7465 6.654 49.0705 6.694 ;
      RECT MASK 1 57.789 6.6625 57.969 6.7025 ;
      RECT MASK 1 60.1675 6.6625 60.3475 6.7025 ;
      RECT MASK 1 65.575 6.6625 65.984 6.7025 ;
      RECT MASK 1 22.7735 6.678 23.4455 6.702 ;
      RECT MASK 1 23.667 6.678 24.1635 6.702 ;
      RECT MASK 1 53.7935 6.774 56.2835 6.814 ;
      RECT MASK 1 58.765 6.782 58.825 6.962 ;
      RECT MASK 1 59.223 6.782 59.283 6.962 ;
      RECT MASK 1 59.681 6.782 59.741 6.962 ;
      RECT MASK 1 60.826 6.782 60.886 6.962 ;
      RECT MASK 1 61.284 6.782 61.344 6.962 ;
      RECT MASK 1 61.742 6.782 61.802 6.962 ;
      RECT MASK 1 62.2 6.782 62.26 6.962 ;
      RECT MASK 1 62.658 6.782 62.718 6.962 ;
      RECT MASK 1 63.116 6.782 63.176 6.962 ;
      RECT MASK 1 63.803 6.782 63.863 6.962 ;
      RECT MASK 1 64.261 6.782 64.321 6.962 ;
      RECT MASK 1 64.719 6.782 64.779 6.962 ;
      RECT MASK 1 46.7465 6.829 49.0705 6.869 ;
      RECT MASK 1 2.5025 6.831 2.7175 6.871 ;
      RECT MASK 1 3.5235 6.831 9.692 6.871 ;
      RECT MASK 1 10.9455 6.831 11.764 6.871 ;
      RECT MASK 1 14.663 6.831 21.414 6.871 ;
      RECT MASK 1 25.523 6.831 32.274 6.871 ;
      RECT MASK 1 35.173 6.831 35.9915 6.871 ;
      RECT MASK 1 37.245 6.831 43.4135 6.871 ;
      RECT MASK 1 44.2195 6.831 44.4345 6.871 ;
      RECT MASK 1 49.9395 6.85 52.6895 6.89 ;
      RECT MASK 1 1.6135 6.9325 1.8575 6.9725 ;
      RECT MASK 1 45.0795 6.9325 45.3235 6.9725 ;
      RECT MASK 1 53.7935 6.949 56.2835 6.989 ;
      RECT MASK 1 46.7465 6.991 49.0705 7.031 ;
      RECT MASK 1 10.3585 6.9925 10.5385 7.0325 ;
      RECT MASK 1 13.5865 6.9925 13.7665 7.0325 ;
      RECT MASK 1 33.1705 6.9925 33.3505 7.0325 ;
      RECT MASK 1 36.3985 6.9925 36.5785 7.0325 ;
      RECT MASK 1 116.154 7.02 116.214 8.07 ;
      RECT MASK 1 116.428 7.02 116.488 8.07 ;
      RECT MASK 1 116.702 7.02 116.762 8.07 ;
      RECT MASK 1 116.976 7.02 117.036 8.07 ;
      RECT MASK 1 117.25 7.02 117.31 8.07 ;
      RECT MASK 1 117.524 7.02 117.584 8.07 ;
      RECT MASK 1 117.798 7.02 117.858 8.07 ;
      RECT MASK 1 118.072 7.02 118.132 8.07 ;
      RECT MASK 1 118.346 7.02 118.406 8.07 ;
      RECT MASK 1 118.62 7.02 118.68 8.07 ;
      RECT MASK 1 118.894 7.02 118.954 8.07 ;
      RECT MASK 1 119.168 7.02 119.228 8.07 ;
      RECT MASK 1 119.442 7.02 119.502 8.07 ;
      RECT MASK 1 119.716 7.02 119.776 8.07 ;
      RECT MASK 1 119.99 7.02 120.05 8.07 ;
      RECT MASK 1 120.264 7.02 120.324 8.07 ;
      RECT MASK 1 120.538 7.02 120.598 8.07 ;
      RECT MASK 1 120.812 7.02 120.872 8.07 ;
      RECT MASK 1 121.086 7.02 121.146 8.07 ;
      RECT MASK 1 121.36 7.02 121.42 8.07 ;
      RECT MASK 1 121.634 7.02 121.694 8.07 ;
      RECT MASK 1 121.908 7.02 121.968 8.07 ;
      RECT MASK 1 122.182 7.02 122.242 8.07 ;
      RECT MASK 1 122.456 7.02 122.516 8.07 ;
      RECT MASK 1 122.73 7.02 122.79 8.07 ;
      RECT MASK 1 123.004 7.02 123.064 8.07 ;
      RECT MASK 1 123.278 7.02 123.338 8.07 ;
      RECT MASK 1 123.552 7.02 123.612 8.07 ;
      RECT MASK 1 123.826 7.02 123.886 8.07 ;
      RECT MASK 1 124.1 7.02 124.16 8.07 ;
      RECT MASK 1 124.374 7.02 124.434 8.07 ;
      RECT MASK 1 124.648 7.02 124.708 8.07 ;
      RECT MASK 1 124.922 7.02 124.982 8.07 ;
      RECT MASK 1 125.196 7.02 125.256 8.07 ;
      RECT MASK 1 125.47 7.02 125.53 8.07 ;
      RECT MASK 1 125.744 7.02 125.804 8.07 ;
      RECT MASK 1 126.018 7.02 126.078 8.07 ;
      RECT MASK 1 126.292 7.02 126.352 8.07 ;
      RECT MASK 1 126.566 7.02 126.626 8.07 ;
      RECT MASK 1 126.84 7.02 126.9 8.07 ;
      RECT MASK 1 127.114 7.02 127.174 8.07 ;
      RECT MASK 1 127.388 7.02 127.448 8.07 ;
      RECT MASK 1 127.662 7.02 127.722 8.07 ;
      RECT MASK 1 127.936 7.02 127.996 8.07 ;
      RECT MASK 1 128.21 7.02 128.27 8.07 ;
      RECT MASK 1 22.2135 7.038 23.3235 7.062 ;
      RECT MASK 1 23.6135 7.038 24.7235 7.062 ;
      RECT MASK 1 83.7875 7.06 91.6835 7.1 ;
      RECT MASK 1 95.0215 7.06 102.9175 7.1 ;
      RECT MASK 1 65.0585 7.082 65.949 7.11 ;
      RECT MASK 1 2.4035 7.112 2.4635 7.292 ;
      RECT MASK 1 2.8615 7.112 2.9215 7.292 ;
      RECT MASK 1 3.3195 7.112 3.3795 7.292 ;
      RECT MASK 1 3.5485 7.112 3.6085 7.292 ;
      RECT MASK 1 3.7775 7.112 3.8375 7.292 ;
      RECT MASK 1 4.0065 7.112 4.0665 7.292 ;
      RECT MASK 1 4.2355 7.112 4.2955 7.292 ;
      RECT MASK 1 4.4645 7.112 4.5245 7.292 ;
      RECT MASK 1 4.6935 7.112 4.7535 7.292 ;
      RECT MASK 1 4.9225 7.112 4.9825 7.292 ;
      RECT MASK 1 5.1515 7.112 5.2115 7.292 ;
      RECT MASK 1 5.6095 7.112 5.6695 7.292 ;
      RECT MASK 1 6.0675 7.112 6.1275 7.292 ;
      RECT MASK 1 6.5255 7.112 6.5855 7.292 ;
      RECT MASK 1 6.9835 7.112 7.0435 7.292 ;
      RECT MASK 1 7.4415 7.112 7.5015 7.292 ;
      RECT MASK 1 7.8995 7.112 7.9595 7.292 ;
      RECT MASK 1 8.3575 7.112 8.4175 7.292 ;
      RECT MASK 1 8.8155 7.112 8.8755 7.292 ;
      RECT MASK 1 9.0445 7.112 9.1045 7.292 ;
      RECT MASK 1 9.2735 7.112 9.3335 7.292 ;
      RECT MASK 1 9.5025 7.112 9.5625 7.292 ;
      RECT MASK 1 9.7315 7.112 9.7915 7.292 ;
      RECT MASK 1 11.3455 7.112 11.4055 7.292 ;
      RECT MASK 1 11.8035 7.112 11.8635 7.292 ;
      RECT MASK 1 12.2615 7.112 12.3215 7.292 ;
      RECT MASK 1 12.7195 7.112 12.7795 7.292 ;
      RECT MASK 1 14.5735 7.112 14.6335 7.292 ;
      RECT MASK 1 15.0315 7.112 15.0915 7.292 ;
      RECT MASK 1 15.4895 7.112 15.5495 7.292 ;
      RECT MASK 1 15.9475 7.112 16.0075 7.292 ;
      RECT MASK 1 16.4055 7.112 16.4655 7.292 ;
      RECT MASK 1 16.8635 7.112 16.9235 7.292 ;
      RECT MASK 1 17.3215 7.112 17.3815 7.292 ;
      RECT MASK 1 17.7795 7.112 17.8395 7.292 ;
      RECT MASK 1 18.2375 7.112 18.2975 7.292 ;
      RECT MASK 1 18.6955 7.112 18.7555 7.292 ;
      RECT MASK 1 19.1535 7.112 19.2135 7.292 ;
      RECT MASK 1 19.6115 7.112 19.6715 7.292 ;
      RECT MASK 1 20.0695 7.112 20.1295 7.292 ;
      RECT MASK 1 20.5275 7.112 20.5875 7.292 ;
      RECT MASK 1 20.9855 7.112 21.0455 7.292 ;
      RECT MASK 1 21.4435 7.112 21.5035 7.292 ;
      RECT MASK 1 25.4335 7.112 25.4935 7.292 ;
      RECT MASK 1 25.8915 7.112 25.9515 7.292 ;
      RECT MASK 1 26.3495 7.112 26.4095 7.292 ;
      RECT MASK 1 26.8075 7.112 26.8675 7.292 ;
      RECT MASK 1 27.2655 7.112 27.3255 7.292 ;
      RECT MASK 1 27.7235 7.112 27.7835 7.292 ;
      RECT MASK 1 28.1815 7.112 28.2415 7.292 ;
      RECT MASK 1 28.6395 7.112 28.6995 7.292 ;
      RECT MASK 1 29.0975 7.112 29.1575 7.292 ;
      RECT MASK 1 29.5555 7.112 29.6155 7.292 ;
      RECT MASK 1 30.0135 7.112 30.0735 7.292 ;
      RECT MASK 1 30.4715 7.112 30.5315 7.292 ;
      RECT MASK 1 30.9295 7.112 30.9895 7.292 ;
      RECT MASK 1 31.3875 7.112 31.4475 7.292 ;
      RECT MASK 1 31.8455 7.112 31.9055 7.292 ;
      RECT MASK 1 32.3035 7.112 32.3635 7.292 ;
      RECT MASK 1 34.1575 7.112 34.2175 7.292 ;
      RECT MASK 1 34.6155 7.112 34.6755 7.292 ;
      RECT MASK 1 35.0735 7.112 35.1335 7.292 ;
      RECT MASK 1 35.5315 7.112 35.5915 7.292 ;
      RECT MASK 1 37.1455 7.112 37.2055 7.292 ;
      RECT MASK 1 37.3745 7.112 37.4345 7.292 ;
      RECT MASK 1 37.6035 7.112 37.6635 7.292 ;
      RECT MASK 1 37.8325 7.112 37.8925 7.292 ;
      RECT MASK 1 38.0615 7.112 38.1215 7.292 ;
      RECT MASK 1 38.5195 7.112 38.5795 7.292 ;
      RECT MASK 1 38.9775 7.112 39.0375 7.292 ;
      RECT MASK 1 39.4355 7.112 39.4955 7.292 ;
      RECT MASK 1 39.8935 7.112 39.9535 7.292 ;
      RECT MASK 1 40.3515 7.112 40.4115 7.292 ;
      RECT MASK 1 40.8095 7.112 40.8695 7.292 ;
      RECT MASK 1 41.2675 7.112 41.3275 7.292 ;
      RECT MASK 1 41.7255 7.112 41.7855 7.292 ;
      RECT MASK 1 41.9545 7.112 42.0145 7.292 ;
      RECT MASK 1 42.1835 7.112 42.2435 7.292 ;
      RECT MASK 1 42.4125 7.112 42.4725 7.292 ;
      RECT MASK 1 42.6415 7.112 42.7015 7.292 ;
      RECT MASK 1 42.8705 7.112 42.9305 7.292 ;
      RECT MASK 1 43.0995 7.112 43.1595 7.292 ;
      RECT MASK 1 43.3285 7.112 43.3885 7.292 ;
      RECT MASK 1 43.5575 7.112 43.6175 7.292 ;
      RECT MASK 1 44.0155 7.112 44.0755 7.292 ;
      RECT MASK 1 44.4735 7.112 44.5335 7.292 ;
      RECT MASK 1 22.2135 7.128 23.3235 7.152 ;
      RECT MASK 1 23.6135 7.128 24.7235 7.152 ;
      RECT MASK 1 46.7465 7.166 49.0705 7.206 ;
      RECT MASK 1 49.9495 7.17 50.1295 7.23 ;
      RECT MASK 1 50.2495 7.17 50.4695 7.23 ;
      RECT MASK 1 50.6135 7.17 50.7935 7.23 ;
      RECT MASK 1 50.9135 7.17 51.1335 7.23 ;
      RECT MASK 1 51.2775 7.17 51.4575 7.23 ;
      RECT MASK 1 51.5775 7.17 51.7975 7.23 ;
      RECT MASK 1 51.9415 7.17 52.1215 7.23 ;
      RECT MASK 1 52.2415 7.17 52.4615 7.23 ;
      RECT MASK 1 22.2135 7.218 23.3235 7.242 ;
      RECT MASK 1 23.6135 7.218 24.7235 7.242 ;
      RECT MASK 1 53.9045 7.27 56.1725 7.31 ;
      RECT MASK 1 65.0585 7.29 65.949 7.318 ;
      RECT MASK 1 83.8025 7.29 83.8825 8.13 ;
      RECT MASK 1 91.5885 7.29 91.6685 8.13 ;
      RECT MASK 1 95.0365 7.29 95.1165 8.13 ;
      RECT MASK 1 102.8225 7.29 102.9025 8.13 ;
      RECT MASK 1 46.9055 7.333 47.1235 7.373 ;
      RECT MASK 1 47.2375 7.333 47.4555 7.373 ;
      RECT MASK 1 47.5695 7.333 47.7875 7.373 ;
      RECT MASK 1 47.9365 7.333 48.2855 7.373 ;
      RECT MASK 1 50.1905 7.41 50.3705 7.47 ;
      RECT MASK 1 50.5105 7.41 50.6905 7.47 ;
      RECT MASK 1 50.8545 7.41 51.0345 7.47 ;
      RECT MASK 1 51.1745 7.41 51.3545 7.47 ;
      RECT MASK 1 51.5185 7.41 51.6985 7.47 ;
      RECT MASK 1 51.8385 7.41 52.0185 7.47 ;
      RECT MASK 1 52.1825 7.41 52.3625 7.47 ;
      RECT MASK 1 52.5025 7.41 52.6825 7.47 ;
      RECT MASK 1 48.8145 7.4275 48.9945 7.4675 ;
      RECT MASK 1 58.765 7.438 58.825 7.618 ;
      RECT MASK 1 59.223 7.438 59.283 7.618 ;
      RECT MASK 1 59.681 7.438 59.741 7.618 ;
      RECT MASK 1 60.826 7.438 60.886 7.618 ;
      RECT MASK 1 61.284 7.438 61.344 7.618 ;
      RECT MASK 1 61.742 7.438 61.802 7.618 ;
      RECT MASK 1 62.2 7.438 62.26 7.618 ;
      RECT MASK 1 62.658 7.438 62.718 7.618 ;
      RECT MASK 1 63.116 7.438 63.176 7.618 ;
      RECT MASK 1 63.803 7.438 63.863 7.618 ;
      RECT MASK 1 64.261 7.438 64.321 7.618 ;
      RECT MASK 1 64.719 7.438 64.779 7.618 ;
      RECT MASK 1 47.0715 7.517 47.2515 7.557 ;
      RECT MASK 1 47.4035 7.517 47.5835 7.557 ;
      RECT MASK 1 47.7355 7.517 47.9155 7.557 ;
      RECT MASK 1 48.2335 7.517 48.4135 7.557 ;
      RECT MASK 1 84.1235 7.53 84.461 7.59 ;
      RECT MASK 1 84.6 7.53 86.2935 7.59 ;
      RECT MASK 1 86.4285 7.53 88.125 7.59 ;
      RECT MASK 1 88.264 7.53 88.6045 7.59 ;
      RECT MASK 1 88.722 7.53 89.041 7.59 ;
      RECT MASK 1 89.18 7.53 89.499 7.59 ;
      RECT MASK 1 89.608 7.53 89.957 7.59 ;
      RECT MASK 1 90.0845 7.53 90.415 7.59 ;
      RECT MASK 1 90.554 7.53 90.904 7.59 ;
      RECT MASK 1 91.012 7.53 91.4125 7.59 ;
      RECT MASK 1 95.2925 7.53 95.693 7.59 ;
      RECT MASK 1 95.801 7.53 96.151 7.59 ;
      RECT MASK 1 96.29 7.53 96.6205 7.59 ;
      RECT MASK 1 96.748 7.53 97.097 7.59 ;
      RECT MASK 1 97.206 7.53 97.525 7.59 ;
      RECT MASK 1 97.664 7.53 97.983 7.59 ;
      RECT MASK 1 98.1005 7.53 98.441 7.59 ;
      RECT MASK 1 98.58 7.53 100.2765 7.59 ;
      RECT MASK 1 100.4115 7.53 102.105 7.59 ;
      RECT MASK 1 102.244 7.53 102.5815 7.59 ;
      RECT MASK 1 50.1675 7.65 50.3475 7.71 ;
      RECT MASK 1 50.5105 7.65 50.6905 7.71 ;
      RECT MASK 1 50.8315 7.65 51.0115 7.71 ;
      RECT MASK 1 51.1745 7.65 51.3545 7.71 ;
      RECT MASK 1 51.4955 7.65 51.6755 7.71 ;
      RECT MASK 1 51.8385 7.65 52.0185 7.71 ;
      RECT MASK 1 52.1595 7.65 52.3395 7.71 ;
      RECT MASK 1 52.5025 7.65 52.6825 7.71 ;
      RECT MASK 1 57.789 7.6975 57.969 7.7375 ;
      RECT MASK 1 60.1675 7.6975 60.3475 7.7375 ;
      RECT MASK 1 65.575 7.6975 65.984 7.7375 ;
      RECT MASK 1 47.0715 7.743 47.2515 7.783 ;
      RECT MASK 1 47.4035 7.743 47.5835 7.783 ;
      RECT MASK 1 47.7355 7.743 47.9155 7.783 ;
      RECT MASK 1 48.2335 7.743 48.4135 7.783 ;
      RECT MASK 1 1.6805 7.75 13.9525 7.79 ;
      RECT MASK 1 14.3195 7.75 21.7575 7.79 ;
      RECT MASK 1 25.1795 7.75 32.6175 7.79 ;
      RECT MASK 1 32.9845 7.75 45.2565 7.79 ;
      RECT MASK 1 61.259 7.758 62.6185 7.798 ;
      RECT MASK 1 86.5465 7.772 91.4125 7.832 ;
      RECT MASK 1 95.2925 7.772 100.1585 7.832 ;
      RECT MASK 1 48.8145 7.8325 48.9945 7.8725 ;
      RECT MASK 1 49.9465 7.89 50.1265 7.95 ;
      RECT MASK 1 50.2665 7.89 50.4465 7.95 ;
      RECT MASK 1 50.6105 7.89 50.7905 7.95 ;
      RECT MASK 1 50.9305 7.89 51.1105 7.95 ;
      RECT MASK 1 51.2745 7.89 51.4545 7.95 ;
      RECT MASK 1 51.5945 7.89 51.7745 7.95 ;
      RECT MASK 1 51.9385 7.89 52.1185 7.95 ;
      RECT MASK 1 52.2585 7.89 52.4385 7.95 ;
      RECT MASK 1 46.9055 7.927 47.1235 7.967 ;
      RECT MASK 1 47.2375 7.927 47.4555 7.967 ;
      RECT MASK 1 47.5695 7.927 47.7875 7.967 ;
      RECT MASK 1 47.9365 7.927 48.1465 7.967 ;
      RECT MASK 1 58.74 7.96 64.804 8 ;
      RECT MASK 1 46.7465 8.094 49.0705 8.134 ;
      RECT MASK 1 49.8465 8.13 52.7825 8.19 ;
      RECT MASK 1 61.3835 8.162 62.743 8.202 ;
      RECT MASK 1 1.6805 8.17 13.9525 8.21 ;
      RECT MASK 1 14.3195 8.17 21.7575 8.21 ;
      RECT MASK 1 57.789 8.2225 57.969 8.2625 ;
      RECT MASK 1 46.7465 8.269 49.0705 8.309 ;
      RECT MASK 1 83.7875 8.32 91.6835 8.36 ;
      RECT MASK 1 95.0215 8.32 102.9175 8.36 ;
      RECT MASK 1 58.765 8.342 58.825 8.522 ;
      RECT MASK 1 59.223 8.342 59.283 8.522 ;
      RECT MASK 1 59.681 8.342 59.741 8.522 ;
      RECT MASK 1 60.826 8.342 60.886 8.522 ;
      RECT MASK 1 61.284 8.342 61.344 8.522 ;
      RECT MASK 1 61.742 8.342 61.802 8.522 ;
      RECT MASK 1 62.2 8.342 62.26 8.522 ;
      RECT MASK 1 62.658 8.342 62.718 8.522 ;
      RECT MASK 1 63.116 8.342 63.176 8.522 ;
      RECT MASK 1 63.803 8.342 63.863 8.522 ;
      RECT MASK 1 64.261 8.342 64.321 8.522 ;
      RECT MASK 1 64.719 8.342 64.779 8.522 ;
      RECT MASK 1 60.1675 8.3425 60.3475 8.3825 ;
      RECT MASK 1 65.575 8.3425 65.984 8.3825 ;
      RECT MASK 1 49.9415 8.37 52.7045 8.43 ;
      RECT MASK 1 46.7465 8.431 49.0705 8.471 ;
      RECT MASK 1 67.634 8.59 70.721 8.63 ;
      RECT MASK 1 46.7465 8.606 49.0705 8.646 ;
      RECT MASK 1 50.1675 8.61 50.4465 8.67 ;
      RECT MASK 1 50.8315 8.61 51.1105 8.67 ;
      RECT MASK 1 51.4955 8.61 51.7745 8.67 ;
      RECT MASK 1 52.1595 8.61 52.4385 8.67 ;
      RECT MASK 1 31.5485 8.62 39.1995 8.66 ;
      RECT MASK 1 53.7665 8.62 56.1665 8.66 ;
      RECT MASK 1 65.0475 8.642 65.949 8.67 ;
      RECT MASK 1 2.4035 8.668 2.4635 8.848 ;
      RECT MASK 1 2.8615 8.668 2.9215 8.848 ;
      RECT MASK 1 3.3195 8.668 3.3795 8.848 ;
      RECT MASK 1 3.5485 8.668 3.6085 8.848 ;
      RECT MASK 1 3.7775 8.668 3.8375 8.848 ;
      RECT MASK 1 4.0065 8.668 4.0665 8.848 ;
      RECT MASK 1 4.2355 8.668 4.2955 8.848 ;
      RECT MASK 1 4.4645 8.668 4.5245 8.848 ;
      RECT MASK 1 4.6935 8.668 4.7535 8.848 ;
      RECT MASK 1 4.9225 8.668 4.9825 8.848 ;
      RECT MASK 1 5.1515 8.668 5.2115 8.848 ;
      RECT MASK 1 5.6095 8.668 5.6695 8.848 ;
      RECT MASK 1 6.0675 8.668 6.1275 8.848 ;
      RECT MASK 1 6.5255 8.668 6.5855 8.848 ;
      RECT MASK 1 6.9835 8.668 7.0435 8.848 ;
      RECT MASK 1 7.4415 8.668 7.5015 8.848 ;
      RECT MASK 1 7.8995 8.668 7.9595 8.848 ;
      RECT MASK 1 8.3575 8.668 8.4175 8.848 ;
      RECT MASK 1 8.8155 8.668 8.8755 8.848 ;
      RECT MASK 1 9.0445 8.668 9.1045 8.848 ;
      RECT MASK 1 9.2735 8.668 9.3335 8.848 ;
      RECT MASK 1 9.5025 8.668 9.5625 8.848 ;
      RECT MASK 1 9.7315 8.668 9.7915 8.848 ;
      RECT MASK 1 11.3455 8.668 11.4055 8.848 ;
      RECT MASK 1 11.8035 8.668 11.8635 8.848 ;
      RECT MASK 1 12.2615 8.668 12.3215 8.848 ;
      RECT MASK 1 12.7195 8.668 12.7795 8.848 ;
      RECT MASK 1 14.5735 8.668 14.6335 8.848 ;
      RECT MASK 1 15.0315 8.668 15.0915 8.848 ;
      RECT MASK 1 15.4895 8.668 15.5495 8.848 ;
      RECT MASK 1 15.9475 8.668 16.0075 8.848 ;
      RECT MASK 1 16.4055 8.668 16.4655 8.848 ;
      RECT MASK 1 16.8635 8.668 16.9235 8.848 ;
      RECT MASK 1 17.3215 8.668 17.3815 8.848 ;
      RECT MASK 1 17.7795 8.668 17.8395 8.848 ;
      RECT MASK 1 18.2375 8.668 18.2975 8.848 ;
      RECT MASK 1 18.6955 8.668 18.7555 8.848 ;
      RECT MASK 1 19.1535 8.668 19.2135 8.848 ;
      RECT MASK 1 19.6115 8.668 19.6715 8.848 ;
      RECT MASK 1 20.0695 8.668 20.1295 8.848 ;
      RECT MASK 1 20.5275 8.668 20.5875 8.848 ;
      RECT MASK 1 20.9855 8.668 21.0455 8.848 ;
      RECT MASK 1 21.4435 8.668 21.5035 8.848 ;
      RECT MASK 1 72.7245 8.68 76.9845 8.72 ;
      RECT MASK 1 109.7205 8.68 113.9805 8.72 ;
      RECT MASK 1 22.2135 8.718 23.3235 8.742 ;
      RECT MASK 1 116.154 8.73 116.214 9.78 ;
      RECT MASK 1 116.428 8.73 116.488 9.78 ;
      RECT MASK 1 116.702 8.73 116.762 9.78 ;
      RECT MASK 1 116.976 8.73 117.036 9.78 ;
      RECT MASK 1 117.25 8.73 117.31 9.78 ;
      RECT MASK 1 117.524 8.73 117.584 9.78 ;
      RECT MASK 1 117.798 8.73 117.858 9.78 ;
      RECT MASK 1 118.072 8.73 118.132 9.78 ;
      RECT MASK 1 118.346 8.73 118.406 9.78 ;
      RECT MASK 1 118.62 8.73 118.68 9.78 ;
      RECT MASK 1 118.894 8.73 118.954 9.78 ;
      RECT MASK 1 119.168 8.73 119.228 9.78 ;
      RECT MASK 1 119.442 8.73 119.502 9.78 ;
      RECT MASK 1 119.716 8.73 119.776 9.78 ;
      RECT MASK 1 119.99 8.73 120.05 9.78 ;
      RECT MASK 1 120.264 8.73 120.324 9.78 ;
      RECT MASK 1 120.538 8.73 120.598 9.78 ;
      RECT MASK 1 120.812 8.73 120.872 9.78 ;
      RECT MASK 1 121.086 8.73 121.146 9.78 ;
      RECT MASK 1 121.36 8.73 121.42 9.78 ;
      RECT MASK 1 121.634 8.73 121.694 9.78 ;
      RECT MASK 1 121.908 8.73 121.968 9.78 ;
      RECT MASK 1 122.182 8.73 122.242 9.78 ;
      RECT MASK 1 122.456 8.73 122.516 9.78 ;
      RECT MASK 1 122.73 8.73 122.79 9.78 ;
      RECT MASK 1 123.004 8.73 123.064 9.78 ;
      RECT MASK 1 123.278 8.73 123.338 9.78 ;
      RECT MASK 1 123.552 8.73 123.612 9.78 ;
      RECT MASK 1 123.826 8.73 123.886 9.78 ;
      RECT MASK 1 124.1 8.73 124.16 9.78 ;
      RECT MASK 1 124.374 8.73 124.434 9.78 ;
      RECT MASK 1 124.648 8.73 124.708 9.78 ;
      RECT MASK 1 124.922 8.73 124.982 9.78 ;
      RECT MASK 1 125.196 8.73 125.256 9.78 ;
      RECT MASK 1 125.47 8.73 125.53 9.78 ;
      RECT MASK 1 125.744 8.73 125.804 9.78 ;
      RECT MASK 1 126.018 8.73 126.078 9.78 ;
      RECT MASK 1 126.292 8.73 126.352 9.78 ;
      RECT MASK 1 126.566 8.73 126.626 9.78 ;
      RECT MASK 1 126.84 8.73 126.9 9.78 ;
      RECT MASK 1 127.114 8.73 127.174 9.78 ;
      RECT MASK 1 127.388 8.73 127.448 9.78 ;
      RECT MASK 1 127.662 8.73 127.722 9.78 ;
      RECT MASK 1 127.936 8.73 127.996 9.78 ;
      RECT MASK 1 128.21 8.73 128.27 9.78 ;
      RECT MASK 1 46.9055 8.773 47.1235 8.813 ;
      RECT MASK 1 47.2375 8.773 47.4555 8.813 ;
      RECT MASK 1 47.6045 8.773 47.8145 8.813 ;
      RECT MASK 1 48.0675 8.773 48.2855 8.813 ;
      RECT MASK 1 22.2135 8.808 23.3235 8.832 ;
      RECT MASK 1 62.5395 8.85 62.743 8.878 ;
      RECT MASK 1 65.839 8.85 66.042 8.878 ;
      RECT MASK 1 48.8145 8.8675 48.9945 8.9075 ;
      RECT MASK 1 22.2135 8.898 23.3235 8.922 ;
      RECT MASK 1 67.46 8.911 70.895 8.951 ;
      RECT MASK 1 10.3585 8.9275 10.5385 8.9675 ;
      RECT MASK 1 13.5865 8.9275 13.7665 8.9675 ;
      RECT MASK 1 31.3665 8.941 39.3815 8.981 ;
      RECT MASK 1 53.5925 8.941 56.3405 8.981 ;
      RECT MASK 1 47.0715 8.957 47.2515 8.997 ;
      RECT MASK 1 47.4035 8.957 47.5835 8.997 ;
      RECT MASK 1 47.9015 8.957 48.0815 8.997 ;
      RECT MASK 1 48.2335 8.957 48.4135 8.997 ;
      RECT MASK 1 49.9395 8.98 52.6895 9.02 ;
      RECT MASK 1 1.6135 8.9875 1.8575 9.0275 ;
      RECT MASK 1 58.536 8.998 58.596 9.178 ;
      RECT MASK 1 58.994 8.998 59.054 9.178 ;
      RECT MASK 1 59.452 8.998 59.512 9.178 ;
      RECT MASK 1 59.91 8.998 59.97 9.178 ;
      RECT MASK 1 60.368 8.998 60.428 9.178 ;
      RECT MASK 1 62.887 8.998 62.947 9.178 ;
      RECT MASK 1 63.345 8.998 63.405 9.178 ;
      RECT MASK 1 63.803 8.998 63.863 9.178 ;
      RECT MASK 1 64.261 8.998 64.321 9.178 ;
      RECT MASK 1 64.719 8.998 64.779 9.178 ;
      RECT MASK 1 65.177 8.998 65.237 9.178 ;
      RECT MASK 1 65.635 8.998 65.695 9.178 ;
      RECT MASK 1 68.346 9.071 68.406 9.292 ;
      RECT MASK 1 68.575 9.071 68.635 9.292 ;
      RECT MASK 1 68.804 9.071 68.864 9.292 ;
      RECT MASK 1 69.033 9.071 69.093 9.292 ;
      RECT MASK 1 69.262 9.071 69.322 9.292 ;
      RECT MASK 1 69.491 9.071 69.551 9.292 ;
      RECT MASK 1 69.949 9.071 70.009 9.292 ;
      RECT MASK 1 2.5025 9.089 2.7175 9.129 ;
      RECT MASK 1 3.5235 9.089 9.692 9.129 ;
      RECT MASK 1 10.9455 9.089 11.764 9.129 ;
      RECT MASK 1 14.663 9.089 21.414 9.129 ;
      RECT MASK 1 54.4785 9.101 54.5385 9.322 ;
      RECT MASK 1 54.7075 9.101 54.7675 9.322 ;
      RECT MASK 1 54.9365 9.101 54.9965 9.322 ;
      RECT MASK 1 55.1655 9.101 55.2255 9.322 ;
      RECT MASK 1 55.3945 9.101 55.4545 9.322 ;
      RECT MASK 1 32.0535 9.116 38.6945 9.156 ;
      RECT MASK 1 60.995 9.1375 61.404 9.1775 ;
      RECT MASK 1 61.911 9.1375 62.091 9.1775 ;
      RECT MASK 1 47.0715 9.183 47.2515 9.223 ;
      RECT MASK 1 47.4035 9.183 47.5835 9.223 ;
      RECT MASK 1 47.9015 9.183 48.0815 9.223 ;
      RECT MASK 1 48.2335 9.183 48.4135 9.223 ;
      RECT MASK 1 57.789 9.2575 57.969 9.2975 ;
      RECT MASK 1 21.99 9.258 23.1635 9.282 ;
      RECT MASK 1 48.8145 9.2725 48.9945 9.3125 ;
      RECT MASK 1 2.5025 9.291 2.7175 9.331 ;
      RECT MASK 1 2.8365 9.291 4.196 9.331 ;
      RECT MASK 1 5.7055 9.291 8.57 9.331 ;
      RECT MASK 1 9.373 9.291 10.0665 9.331 ;
      RECT MASK 1 11.0705 9.291 11.764 9.331 ;
      RECT MASK 1 12.361 9.291 13.0765 9.331 ;
      RECT MASK 1 14.663 9.291 21.414 9.331 ;
      RECT MASK 1 62.633 9.318 63.0765 9.358 ;
      RECT MASK 1 63.6735 9.318 65.3665 9.358 ;
      RECT MASK 1 65.5055 9.318 65.949 9.358 ;
      RECT MASK 1 67.567 9.3475 67.811 9.3875 ;
      RECT MASK 1 70.544 9.3475 70.788 9.3875 ;
      RECT MASK 1 22.2135 9.348 23.3235 9.372 ;
      RECT MASK 1 32.536 9.366 32.7855 9.406 ;
      RECT MASK 1 33.452 9.366 33.7015 9.406 ;
      RECT MASK 1 34.368 9.366 34.6175 9.406 ;
      RECT MASK 1 35.284 9.366 35.5335 9.406 ;
      RECT MASK 1 36.2 9.366 36.4495 9.406 ;
      RECT MASK 1 37.116 9.366 37.3655 9.406 ;
      RECT MASK 1 38.032 9.366 38.2815 9.406 ;
      RECT MASK 1 46.9055 9.367 47.1235 9.407 ;
      RECT MASK 1 47.2375 9.367 47.4555 9.407 ;
      RECT MASK 1 47.6045 9.367 47.9535 9.407 ;
      RECT MASK 1 48.0675 9.367 48.2855 9.407 ;
      RECT MASK 1 31.4735 9.3775 31.7175 9.4175 ;
      RECT MASK 1 39.0305 9.3775 39.2745 9.4175 ;
      RECT MASK 1 53.6995 9.3775 53.9435 9.4175 ;
      RECT MASK 1 55.9895 9.3775 56.2335 9.4175 ;
      RECT MASK 1 1.6135 9.3925 1.8575 9.4325 ;
      RECT MASK 1 49.9395 9.4 52.6895 9.44 ;
      RECT MASK 1 22.4135 9.438 22.7135 9.462 ;
      RECT MASK 1 22.8235 9.438 23.1235 9.462 ;
      RECT MASK 1 10.3585 9.4525 10.5385 9.4925 ;
      RECT MASK 1 13.5865 9.4525 13.7665 9.4925 ;
      RECT MASK 1 22.4135 9.528 22.7135 9.552 ;
      RECT MASK 1 22.8235 9.528 23.1235 9.552 ;
      RECT MASK 1 46.7465 9.534 49.0705 9.574 ;
      RECT MASK 1 2.8615 9.571 2.9215 9.752 ;
      RECT MASK 1 5.1515 9.571 5.2115 9.752 ;
      RECT MASK 1 2.4035 9.572 2.4635 9.752 ;
      RECT MASK 1 3.3195 9.572 3.3795 9.752 ;
      RECT MASK 1 3.5485 9.572 3.6085 9.752 ;
      RECT MASK 1 3.7775 9.572 3.8375 9.752 ;
      RECT MASK 1 4.0065 9.572 4.0665 9.752 ;
      RECT MASK 1 4.2355 9.572 4.2955 9.752 ;
      RECT MASK 1 4.4645 9.572 4.5245 9.752 ;
      RECT MASK 1 4.6935 9.572 4.7535 9.752 ;
      RECT MASK 1 4.9225 9.572 4.9825 9.752 ;
      RECT MASK 1 5.6095 9.572 5.6695 9.752 ;
      RECT MASK 1 6.0675 9.572 6.1275 9.752 ;
      RECT MASK 1 6.5255 9.572 6.5855 9.752 ;
      RECT MASK 1 6.9835 9.572 7.0435 9.752 ;
      RECT MASK 1 7.4415 9.572 7.5015 9.752 ;
      RECT MASK 1 7.8995 9.572 7.9595 9.752 ;
      RECT MASK 1 8.3575 9.572 8.4175 9.752 ;
      RECT MASK 1 8.8155 9.572 8.8755 9.752 ;
      RECT MASK 1 9.0445 9.572 9.1045 9.752 ;
      RECT MASK 1 9.2735 9.572 9.3335 9.752 ;
      RECT MASK 1 9.5025 9.572 9.5625 9.752 ;
      RECT MASK 1 9.7315 9.572 9.7915 9.752 ;
      RECT MASK 1 11.3455 9.572 11.4055 9.752 ;
      RECT MASK 1 11.8035 9.572 11.8635 9.752 ;
      RECT MASK 1 12.2615 9.572 12.3215 9.752 ;
      RECT MASK 1 12.7195 9.572 12.7795 9.752 ;
      RECT MASK 1 14.5735 9.572 14.6335 9.752 ;
      RECT MASK 1 15.0315 9.572 15.0915 9.752 ;
      RECT MASK 1 15.4895 9.572 15.5495 9.752 ;
      RECT MASK 1 15.9475 9.572 16.0075 9.752 ;
      RECT MASK 1 16.4055 9.572 16.4655 9.752 ;
      RECT MASK 1 16.8635 9.572 16.9235 9.752 ;
      RECT MASK 1 17.3215 9.572 17.3815 9.752 ;
      RECT MASK 1 17.7795 9.572 17.8395 9.752 ;
      RECT MASK 1 18.2375 9.572 18.2975 9.752 ;
      RECT MASK 1 18.6955 9.572 18.7555 9.752 ;
      RECT MASK 1 19.1535 9.572 19.2135 9.752 ;
      RECT MASK 1 19.6115 9.572 19.6715 9.752 ;
      RECT MASK 1 20.0695 9.572 20.1295 9.752 ;
      RECT MASK 1 20.5275 9.572 20.5875 9.752 ;
      RECT MASK 1 20.9855 9.572 21.0455 9.752 ;
      RECT MASK 1 21.4435 9.572 21.5035 9.752 ;
      RECT MASK 1 22.4135 9.618 22.7135 9.642 ;
      RECT MASK 1 22.8235 9.618 23.1235 9.642 ;
      RECT MASK 1 46.7465 9.709 49.0705 9.749 ;
      RECT MASK 1 49.8415 9.71 50.0265 9.77 ;
      RECT MASK 1 62.633 9.722 63.0765 9.762 ;
      RECT MASK 1 63.549 9.722 64.2215 9.762 ;
      RECT MASK 1 64.465 9.722 65.8245 9.762 ;
      RECT MASK 1 67.567 9.7525 67.811 9.7925 ;
      RECT MASK 1 70.544 9.7525 70.788 9.7925 ;
      RECT MASK 1 31.4735 9.7825 31.7175 9.8225 ;
      RECT MASK 1 39.0305 9.7825 39.2745 9.8225 ;
      RECT MASK 1 53.6995 9.7825 53.9435 9.8225 ;
      RECT MASK 1 55.9895 9.7825 56.2335 9.8225 ;
      RECT MASK 1 57.789 9.7825 57.969 9.8225 ;
      RECT MASK 1 60.995 9.7825 61.404 9.8225 ;
      RECT MASK 1 61.911 9.7825 62.091 9.8225 ;
      RECT MASK 1 32.536 9.794 32.7855 9.834 ;
      RECT MASK 1 33.452 9.794 33.7015 9.834 ;
      RECT MASK 1 34.368 9.794 34.6175 9.834 ;
      RECT MASK 1 35.284 9.794 35.5335 9.834 ;
      RECT MASK 1 36.2 9.794 36.4495 9.834 ;
      RECT MASK 1 37.116 9.794 37.3655 9.834 ;
      RECT MASK 1 38.032 9.794 38.2815 9.834 ;
      RECT MASK 1 68.346 9.848 68.406 10.069 ;
      RECT MASK 1 68.575 9.848 68.635 10.069 ;
      RECT MASK 1 68.804 9.848 68.864 10.069 ;
      RECT MASK 1 69.033 9.848 69.093 10.069 ;
      RECT MASK 1 69.262 9.848 69.322 10.069 ;
      RECT MASK 1 69.491 9.848 69.551 10.069 ;
      RECT MASK 1 69.72 9.848 69.78 10.069 ;
      RECT MASK 1 69.949 9.848 70.009 10.069 ;
      RECT MASK 1 54.4785 9.878 54.5385 10.099 ;
      RECT MASK 1 54.7075 9.878 54.7675 10.099 ;
      RECT MASK 1 54.9365 9.878 54.9965 10.099 ;
      RECT MASK 1 55.1655 9.878 55.2255 10.099 ;
      RECT MASK 1 55.3945 9.878 55.4545 10.099 ;
      RECT MASK 1 58.536 9.902 58.596 10.082 ;
      RECT MASK 1 58.994 9.902 59.054 10.082 ;
      RECT MASK 1 59.452 9.902 59.512 10.082 ;
      RECT MASK 1 59.91 9.902 59.97 10.082 ;
      RECT MASK 1 60.368 9.902 60.428 10.082 ;
      RECT MASK 1 62.887 9.902 62.947 10.082 ;
      RECT MASK 1 63.345 9.902 63.405 10.082 ;
      RECT MASK 1 63.803 9.902 63.863 10.082 ;
      RECT MASK 1 64.261 9.902 64.321 10.082 ;
      RECT MASK 1 64.719 9.902 64.779 10.082 ;
      RECT MASK 1 65.177 9.902 65.237 10.082 ;
      RECT MASK 1 65.635 9.902 65.695 10.082 ;
      RECT MASK 1 49.9465 9.93 52.6825 9.99 ;
      RECT MASK 1 22.2235 9.978 23.3235 10.002 ;
      RECT MASK 1 46.8655 10.03 48.9595 10.07 ;
      RECT MASK 1 32.0535 10.044 38.6945 10.084 ;
      RECT MASK 1 50.1525 10.17 50.4695 10.23 ;
      RECT MASK 1 50.8165 10.17 51.1335 10.23 ;
      RECT MASK 1 51.4805 10.17 51.7975 10.23 ;
      RECT MASK 1 52.1445 10.17 52.4615 10.23 ;
      RECT MASK 1 67.46 10.189 70.895 10.229 ;
      RECT MASK 1 62.5395 10.1995 62.743 10.2275 ;
      RECT MASK 1 65.839 10.1995 66.042 10.2275 ;
      RECT MASK 1 1.6805 10.21 10.7245 10.25 ;
      RECT MASK 1 11.1705 10.21 12.9295 10.25 ;
      RECT MASK 1 13.4005 10.21 21.7575 10.25 ;
      RECT MASK 1 31.3665 10.219 39.3815 10.259 ;
      RECT MASK 1 53.5925 10.219 56.3405 10.259 ;
      RECT MASK 1 77.4385 10.39 82.3625 10.43 ;
      RECT MASK 1 104.3425 10.39 109.2665 10.43 ;
      RECT MASK 1 116.154 10.44 116.214 11.49 ;
      RECT MASK 1 116.428 10.44 116.488 11.49 ;
      RECT MASK 1 116.702 10.44 116.762 11.49 ;
      RECT MASK 1 116.976 10.44 117.036 11.49 ;
      RECT MASK 1 117.25 10.44 117.31 11.49 ;
      RECT MASK 1 117.524 10.44 117.584 11.49 ;
      RECT MASK 1 117.798 10.44 117.858 11.49 ;
      RECT MASK 1 118.072 10.44 118.132 11.49 ;
      RECT MASK 1 118.346 10.44 118.406 11.49 ;
      RECT MASK 1 118.62 10.44 118.68 11.49 ;
      RECT MASK 1 118.894 10.44 118.954 11.49 ;
      RECT MASK 1 119.168 10.44 119.228 11.49 ;
      RECT MASK 1 119.442 10.44 119.502 11.49 ;
      RECT MASK 1 119.716 10.44 119.776 11.49 ;
      RECT MASK 1 119.99 10.44 120.05 11.49 ;
      RECT MASK 1 120.264 10.44 120.324 11.49 ;
      RECT MASK 1 120.538 10.44 120.598 11.49 ;
      RECT MASK 1 120.812 10.44 120.872 11.49 ;
      RECT MASK 1 121.086 10.44 121.146 11.49 ;
      RECT MASK 1 121.36 10.44 121.42 11.49 ;
      RECT MASK 1 121.634 10.44 121.694 11.49 ;
      RECT MASK 1 121.908 10.44 121.968 11.49 ;
      RECT MASK 1 122.182 10.44 122.242 11.49 ;
      RECT MASK 1 122.456 10.44 122.516 11.49 ;
      RECT MASK 1 122.73 10.44 122.79 11.49 ;
      RECT MASK 1 123.004 10.44 123.064 11.49 ;
      RECT MASK 1 123.278 10.44 123.338 11.49 ;
      RECT MASK 1 123.552 10.44 123.612 11.49 ;
      RECT MASK 1 123.826 10.44 123.886 11.49 ;
      RECT MASK 1 124.1 10.44 124.16 11.49 ;
      RECT MASK 1 124.374 10.44 124.434 11.49 ;
      RECT MASK 1 124.648 10.44 124.708 11.49 ;
      RECT MASK 1 124.922 10.44 124.982 11.49 ;
      RECT MASK 1 125.196 10.44 125.256 11.49 ;
      RECT MASK 1 125.47 10.44 125.53 11.49 ;
      RECT MASK 1 125.744 10.44 125.804 11.49 ;
      RECT MASK 1 126.018 10.44 126.078 11.49 ;
      RECT MASK 1 126.292 10.44 126.352 11.49 ;
      RECT MASK 1 126.566 10.44 126.626 11.49 ;
      RECT MASK 1 126.84 10.44 126.9 11.49 ;
      RECT MASK 1 127.114 10.44 127.174 11.49 ;
      RECT MASK 1 127.388 10.44 127.448 11.49 ;
      RECT MASK 1 127.662 10.44 127.722 11.49 ;
      RECT MASK 1 127.936 10.44 127.996 11.49 ;
      RECT MASK 1 128.21 10.44 128.27 11.49 ;
      RECT MASK 1 67.634 10.51 70.721 10.55 ;
      RECT MASK 1 31.5485 10.54 39.1995 10.58 ;
      RECT MASK 1 53.7665 10.54 56.1665 10.58 ;
      RECT MASK 1 57.824 10.54 60.453 10.58 ;
      RECT MASK 1 61.946 10.54 65.984 10.58 ;
      RECT MASK 1 49.9395 10.63 52.6895 10.67 ;
      RECT MASK 1 4.362 11.86 111.8085 11.9 ;
      RECT MASK 1 116.154 12.15 116.214 13.2 ;
      RECT MASK 1 116.428 12.15 116.488 13.2 ;
      RECT MASK 1 116.702 12.15 116.762 13.2 ;
      RECT MASK 1 116.976 12.15 117.036 13.2 ;
      RECT MASK 1 117.25 12.15 117.31 13.2 ;
      RECT MASK 1 117.524 12.15 117.584 13.2 ;
      RECT MASK 1 117.798 12.15 117.858 13.2 ;
      RECT MASK 1 118.072 12.15 118.132 13.2 ;
      RECT MASK 1 118.346 12.15 118.406 13.2 ;
      RECT MASK 1 118.62 12.15 118.68 13.2 ;
      RECT MASK 1 118.894 12.15 118.954 13.2 ;
      RECT MASK 1 119.168 12.15 119.228 13.2 ;
      RECT MASK 1 119.442 12.15 119.502 13.2 ;
      RECT MASK 1 119.716 12.15 119.776 13.2 ;
      RECT MASK 1 119.99 12.15 120.05 13.2 ;
      RECT MASK 1 120.264 12.15 120.324 13.2 ;
      RECT MASK 1 120.538 12.15 120.598 13.2 ;
      RECT MASK 1 120.812 12.15 120.872 13.2 ;
      RECT MASK 1 121.086 12.15 121.146 13.2 ;
      RECT MASK 1 121.36 12.15 121.42 13.2 ;
      RECT MASK 1 121.634 12.15 121.694 13.2 ;
      RECT MASK 1 121.908 12.15 121.968 13.2 ;
      RECT MASK 1 122.182 12.15 122.242 13.2 ;
      RECT MASK 1 122.456 12.15 122.516 13.2 ;
      RECT MASK 1 122.73 12.15 122.79 13.2 ;
      RECT MASK 1 123.004 12.15 123.064 13.2 ;
      RECT MASK 1 123.278 12.15 123.338 13.2 ;
      RECT MASK 1 123.552 12.15 123.612 13.2 ;
      RECT MASK 1 123.826 12.15 123.886 13.2 ;
      RECT MASK 1 124.1 12.15 124.16 13.2 ;
      RECT MASK 1 124.374 12.15 124.434 13.2 ;
      RECT MASK 1 124.648 12.15 124.708 13.2 ;
      RECT MASK 1 124.922 12.15 124.982 13.2 ;
      RECT MASK 1 125.196 12.15 125.256 13.2 ;
      RECT MASK 1 125.47 12.15 125.53 13.2 ;
      RECT MASK 1 125.744 12.15 125.804 13.2 ;
      RECT MASK 1 126.018 12.15 126.078 13.2 ;
      RECT MASK 1 126.292 12.15 126.352 13.2 ;
      RECT MASK 1 126.566 12.15 126.626 13.2 ;
      RECT MASK 1 126.84 12.15 126.9 13.2 ;
      RECT MASK 1 127.114 12.15 127.174 13.2 ;
      RECT MASK 1 127.388 12.15 127.448 13.2 ;
      RECT MASK 1 127.662 12.15 127.722 13.2 ;
      RECT MASK 1 127.936 12.15 127.996 13.2 ;
      RECT MASK 1 128.21 12.15 128.27 13.2 ;
      RECT MASK 1 4.251 12.181 111.819 12.221 ;
      RECT MASK 1 4.251 12.356 111.819 12.396 ;
      RECT MASK 1 8.356 12.523 8.871 12.563 ;
      RECT MASK 1 9.093 12.523 9.608 12.563 ;
      RECT MASK 1 10.016 12.523 10.531 12.563 ;
      RECT MASK 1 10.753 12.523 11.268 12.563 ;
      RECT MASK 1 22.373 12.523 22.888 12.563 ;
      RECT MASK 1 23.296 12.523 23.811 12.563 ;
      RECT MASK 1 24.033 12.523 24.548 12.563 ;
      RECT MASK 1 24.956 12.523 25.471 12.563 ;
      RECT MASK 1 25.651 12.523 26.081 12.563 ;
      RECT MASK 1 26.743 12.523 27.173 12.563 ;
      RECT MASK 1 27.446 12.523 27.629 12.563 ;
      RECT MASK 1 28.403 12.523 28.833 12.563 ;
      RECT MASK 1 28.971 12.523 29.401 12.563 ;
      RECT MASK 1 30.009 12.523 30.192 12.563 ;
      RECT MASK 1 30.631 12.523 31.061 12.563 ;
      RECT MASK 1 31.723 12.523 32.153 12.563 ;
      RECT MASK 1 32.291 12.523 32.721 12.563 ;
      RECT MASK 1 33.383 12.523 33.813 12.563 ;
      RECT MASK 1 34.086 12.523 34.601 12.563 ;
      RECT MASK 1 34.823 12.523 35.338 12.563 ;
      RECT MASK 1 35.653 12.523 36.168 12.563 ;
      RECT MASK 1 36.576 12.523 37.091 12.563 ;
      RECT MASK 1 37.271 12.523 37.701 12.563 ;
      RECT MASK 1 38.363 12.523 38.793 12.563 ;
      RECT MASK 1 38.931 12.523 39.361 12.563 ;
      RECT MASK 1 40.023 12.523 40.453 12.563 ;
      RECT MASK 1 40.726 12.523 40.909 12.563 ;
      RECT MASK 1 41.556 12.523 41.739 12.563 ;
      RECT MASK 1 42.251 12.523 42.681 12.563 ;
      RECT MASK 1 43.343 12.523 43.773 12.563 ;
      RECT MASK 1 43.953 12.523 44.468 12.563 ;
      RECT MASK 1 44.876 12.523 45.391 12.563 ;
      RECT MASK 1 45.706 12.523 46.221 12.563 ;
      RECT MASK 1 46.536 12.523 47.051 12.563 ;
      RECT MASK 1 47.231 12.523 47.661 12.563 ;
      RECT MASK 1 48.323 12.523 48.753 12.563 ;
      RECT MASK 1 48.933 12.523 49.448 12.563 ;
      RECT MASK 1 49.856 12.523 50.371 12.563 ;
      RECT MASK 1 50.593 12.523 51.108 12.563 ;
      RECT MASK 1 51.516 12.523 52.031 12.563 ;
      RECT MASK 1 52.253 12.523 52.768 12.563 ;
      RECT MASK 1 53.176 12.523 53.691 12.563 ;
      RECT MASK 1 53.871 12.523 54.301 12.563 ;
      RECT MASK 1 54.963 12.523 55.393 12.563 ;
      RECT MASK 1 55.573 12.523 55.756 12.563 ;
      RECT MASK 1 56.789 12.523 57.219 12.563 ;
      RECT MASK 1 57.357 12.523 57.787 12.563 ;
      RECT MASK 1 58.322 12.523 58.837 12.563 ;
      RECT MASK 1 59.059 12.523 59.574 12.563 ;
      RECT MASK 1 60.055 12.523 60.238 12.563 ;
      RECT MASK 1 60.719 12.523 61.234 12.563 ;
      RECT MASK 1 61.642 12.523 62.157 12.563 ;
      RECT MASK 1 62.472 12.523 62.655 12.563 ;
      RECT MASK 1 63.429 12.523 63.859 12.563 ;
      RECT MASK 1 63.997 12.523 64.427 12.563 ;
      RECT MASK 1 64.962 12.523 65.477 12.563 ;
      RECT MASK 1 65.699 12.523 66.214 12.563 ;
      RECT MASK 1 66.622 12.523 67.137 12.563 ;
      RECT MASK 1 67.359 12.523 67.874 12.563 ;
      RECT MASK 1 68.282 12.523 68.797 12.563 ;
      RECT MASK 1 69.019 12.523 69.534 12.563 ;
      RECT MASK 1 69.942 12.523 70.457 12.563 ;
      RECT MASK 1 70.679 12.523 71.194 12.563 ;
      RECT MASK 1 71.602 12.523 72.117 12.563 ;
      RECT MASK 1 72.339 12.523 72.854 12.563 ;
      RECT MASK 1 77.319 12.523 77.834 12.563 ;
      RECT MASK 1 78.242 12.523 78.757 12.563 ;
      RECT MASK 1 78.979 12.523 79.494 12.563 ;
      RECT MASK 1 79.902 12.523 80.417 12.563 ;
      RECT MASK 1 83.349 12.523 83.779 12.563 ;
      RECT MASK 1 83.917 12.523 84.347 12.563 ;
      RECT MASK 1 88.939 12.523 89.454 12.563 ;
      RECT MASK 1 89.862 12.523 90.377 12.563 ;
      RECT MASK 1 90.599 12.523 91.114 12.563 ;
      RECT MASK 1 91.522 12.523 92.037 12.563 ;
      RECT MASK 1 101.482 12.523 101.997 12.563 ;
      RECT MASK 1 102.219 12.523 102.734 12.563 ;
      RECT MASK 1 103.142 12.523 103.657 12.563 ;
      RECT MASK 1 103.879 12.523 104.394 12.563 ;
      RECT MASK 1 4.327 12.6175 4.507 12.6575 ;
      RECT MASK 1 111.563 12.6175 111.743 12.6575 ;
      RECT MASK 1 8.228 12.707 8.574 12.747 ;
      RECT MASK 1 9.39 12.707 9.736 12.747 ;
      RECT MASK 1 9.888 12.707 10.234 12.747 ;
      RECT MASK 1 11.05 12.707 11.396 12.747 ;
      RECT MASK 1 22.67 12.707 23.016 12.747 ;
      RECT MASK 1 23.168 12.707 23.514 12.747 ;
      RECT MASK 1 24.33 12.707 24.676 12.747 ;
      RECT MASK 1 24.828 12.707 25.174 12.747 ;
      RECT MASK 1 25.658 12.707 26.336 12.747 ;
      RECT MASK 1 26.488 12.707 27.166 12.747 ;
      RECT MASK 1 27.318 12.707 27.664 12.747 ;
      RECT MASK 1 28.148 12.707 28.826 12.747 ;
      RECT MASK 1 28.978 12.707 29.656 12.747 ;
      RECT MASK 1 29.974 12.707 30.32 12.747 ;
      RECT MASK 1 30.638 12.707 31.316 12.747 ;
      RECT MASK 1 31.468 12.707 32.146 12.747 ;
      RECT MASK 1 32.298 12.707 32.976 12.747 ;
      RECT MASK 1 33.128 12.707 33.806 12.747 ;
      RECT MASK 1 33.958 12.707 34.304 12.747 ;
      RECT MASK 1 35.12 12.707 35.466 12.747 ;
      RECT MASK 1 35.95 12.707 36.296 12.747 ;
      RECT MASK 1 36.448 12.707 36.794 12.747 ;
      RECT MASK 1 37.278 12.707 37.956 12.747 ;
      RECT MASK 1 38.108 12.707 38.786 12.747 ;
      RECT MASK 1 38.938 12.707 39.616 12.747 ;
      RECT MASK 1 39.768 12.707 40.446 12.747 ;
      RECT MASK 1 40.598 12.707 40.944 12.747 ;
      RECT MASK 1 41.428 12.707 41.774 12.747 ;
      RECT MASK 1 42.258 12.707 42.936 12.747 ;
      RECT MASK 1 43.088 12.707 43.766 12.747 ;
      RECT MASK 1 44.25 12.707 44.596 12.747 ;
      RECT MASK 1 44.748 12.707 45.094 12.747 ;
      RECT MASK 1 45.578 12.707 45.924 12.747 ;
      RECT MASK 1 46.408 12.707 46.754 12.747 ;
      RECT MASK 1 47.238 12.707 47.916 12.747 ;
      RECT MASK 1 48.068 12.707 48.746 12.747 ;
      RECT MASK 1 49.23 12.707 49.576 12.747 ;
      RECT MASK 1 49.728 12.707 50.074 12.747 ;
      RECT MASK 1 50.89 12.707 51.236 12.747 ;
      RECT MASK 1 51.388 12.707 51.734 12.747 ;
      RECT MASK 1 52.55 12.707 52.896 12.747 ;
      RECT MASK 1 53.048 12.707 53.394 12.747 ;
      RECT MASK 1 53.878 12.707 54.556 12.747 ;
      RECT MASK 1 54.708 12.707 55.386 12.747 ;
      RECT MASK 1 55.538 12.707 55.884 12.747 ;
      RECT MASK 1 56.534 12.707 57.212 12.747 ;
      RECT MASK 1 57.364 12.707 58.042 12.747 ;
      RECT MASK 1 58.194 12.707 58.54 12.747 ;
      RECT MASK 1 59.356 12.707 59.702 12.747 ;
      RECT MASK 1 60.02 12.707 60.366 12.747 ;
      RECT MASK 1 61.016 12.707 61.362 12.747 ;
      RECT MASK 1 61.514 12.707 61.86 12.747 ;
      RECT MASK 1 62.344 12.707 62.69 12.747 ;
      RECT MASK 1 63.174 12.707 63.852 12.747 ;
      RECT MASK 1 64.004 12.707 64.682 12.747 ;
      RECT MASK 1 64.834 12.707 65.18 12.747 ;
      RECT MASK 1 65.996 12.707 66.342 12.747 ;
      RECT MASK 1 66.494 12.707 66.84 12.747 ;
      RECT MASK 1 67.656 12.707 68.002 12.747 ;
      RECT MASK 1 68.154 12.707 68.5 12.747 ;
      RECT MASK 1 69.316 12.707 69.662 12.747 ;
      RECT MASK 1 69.814 12.707 70.16 12.747 ;
      RECT MASK 1 70.976 12.707 71.322 12.747 ;
      RECT MASK 1 71.474 12.707 71.82 12.747 ;
      RECT MASK 1 72.636 12.707 72.982 12.747 ;
      RECT MASK 1 77.616 12.707 77.962 12.747 ;
      RECT MASK 1 78.114 12.707 78.46 12.747 ;
      RECT MASK 1 79.276 12.707 79.622 12.747 ;
      RECT MASK 1 79.774 12.707 80.12 12.747 ;
      RECT MASK 1 83.094 12.707 83.772 12.747 ;
      RECT MASK 1 83.924 12.707 84.602 12.747 ;
      RECT MASK 1 89.236 12.707 89.582 12.747 ;
      RECT MASK 1 89.734 12.707 90.08 12.747 ;
      RECT MASK 1 90.896 12.707 91.242 12.747 ;
      RECT MASK 1 91.394 12.707 91.74 12.747 ;
      RECT MASK 1 101.354 12.707 101.7 12.747 ;
      RECT MASK 1 102.516 12.707 102.862 12.747 ;
      RECT MASK 1 103.014 12.707 103.36 12.747 ;
      RECT MASK 1 104.176 12.707 104.522 12.747 ;
      RECT MASK 1 8.228 12.933 8.906 12.973 ;
      RECT MASK 1 9.058 12.933 9.736 12.973 ;
      RECT MASK 1 9.888 12.933 10.566 12.973 ;
      RECT MASK 1 10.718 12.933 11.396 12.973 ;
      RECT MASK 1 22.338 12.933 23.016 12.973 ;
      RECT MASK 1 23.168 12.933 23.846 12.973 ;
      RECT MASK 1 23.998 12.933 24.676 12.973 ;
      RECT MASK 1 24.828 12.933 25.506 12.973 ;
      RECT MASK 1 25.658 12.933 26.336 12.973 ;
      RECT MASK 1 26.488 12.933 27.166 12.973 ;
      RECT MASK 1 27.318 12.933 27.664 12.973 ;
      RECT MASK 1 28.148 12.933 28.826 12.973 ;
      RECT MASK 1 28.978 12.933 29.656 12.973 ;
      RECT MASK 1 29.974 12.933 30.32 12.973 ;
      RECT MASK 1 30.638 12.933 31.316 12.973 ;
      RECT MASK 1 31.468 12.933 32.146 12.973 ;
      RECT MASK 1 32.298 12.933 32.976 12.973 ;
      RECT MASK 1 33.128 12.933 33.806 12.973 ;
      RECT MASK 1 33.958 12.933 34.636 12.973 ;
      RECT MASK 1 34.788 12.933 35.466 12.973 ;
      RECT MASK 1 35.618 12.933 36.296 12.973 ;
      RECT MASK 1 36.448 12.933 37.126 12.973 ;
      RECT MASK 1 37.278 12.933 37.956 12.973 ;
      RECT MASK 1 38.108 12.933 38.786 12.973 ;
      RECT MASK 1 38.938 12.933 39.616 12.973 ;
      RECT MASK 1 39.768 12.933 40.446 12.973 ;
      RECT MASK 1 40.598 12.933 40.944 12.973 ;
      RECT MASK 1 41.428 12.933 41.774 12.973 ;
      RECT MASK 1 42.258 12.933 42.936 12.973 ;
      RECT MASK 1 43.088 12.933 43.766 12.973 ;
      RECT MASK 1 43.918 12.933 44.596 12.973 ;
      RECT MASK 1 44.748 12.933 45.426 12.973 ;
      RECT MASK 1 45.578 12.933 46.256 12.973 ;
      RECT MASK 1 46.408 12.933 47.086 12.973 ;
      RECT MASK 1 47.238 12.933 47.916 12.973 ;
      RECT MASK 1 48.068 12.933 48.746 12.973 ;
      RECT MASK 1 48.898 12.933 49.576 12.973 ;
      RECT MASK 1 49.728 12.933 50.406 12.973 ;
      RECT MASK 1 50.558 12.933 51.236 12.973 ;
      RECT MASK 1 51.388 12.933 52.066 12.973 ;
      RECT MASK 1 52.218 12.933 52.896 12.973 ;
      RECT MASK 1 53.048 12.933 53.726 12.973 ;
      RECT MASK 1 53.878 12.933 54.556 12.973 ;
      RECT MASK 1 54.708 12.933 55.386 12.973 ;
      RECT MASK 1 55.538 12.933 55.884 12.973 ;
      RECT MASK 1 56.534 12.933 57.212 12.973 ;
      RECT MASK 1 57.364 12.933 58.042 12.973 ;
      RECT MASK 1 58.194 12.933 58.872 12.973 ;
      RECT MASK 1 59.024 12.933 59.702 12.973 ;
      RECT MASK 1 60.02 12.933 60.366 12.973 ;
      RECT MASK 1 60.684 12.933 61.362 12.973 ;
      RECT MASK 1 61.514 12.933 62.192 12.973 ;
      RECT MASK 1 62.344 12.933 62.69 12.973 ;
      RECT MASK 1 63.174 12.933 63.852 12.973 ;
      RECT MASK 1 64.004 12.933 64.682 12.973 ;
      RECT MASK 1 64.834 12.933 65.512 12.973 ;
      RECT MASK 1 65.664 12.933 66.342 12.973 ;
      RECT MASK 1 66.494 12.933 67.172 12.973 ;
      RECT MASK 1 67.324 12.933 68.002 12.973 ;
      RECT MASK 1 68.154 12.933 68.832 12.973 ;
      RECT MASK 1 68.984 12.933 69.662 12.973 ;
      RECT MASK 1 69.814 12.933 70.492 12.973 ;
      RECT MASK 1 70.644 12.933 71.322 12.973 ;
      RECT MASK 1 71.474 12.933 72.152 12.973 ;
      RECT MASK 1 72.304 12.933 72.982 12.973 ;
      RECT MASK 1 77.284 12.933 77.962 12.973 ;
      RECT MASK 1 78.114 12.933 78.792 12.973 ;
      RECT MASK 1 78.944 12.933 79.622 12.973 ;
      RECT MASK 1 79.774 12.933 80.452 12.973 ;
      RECT MASK 1 83.094 12.933 83.772 12.973 ;
      RECT MASK 1 83.924 12.933 84.602 12.973 ;
      RECT MASK 1 88.904 12.933 89.582 12.973 ;
      RECT MASK 1 89.734 12.933 90.412 12.973 ;
      RECT MASK 1 90.564 12.933 91.242 12.973 ;
      RECT MASK 1 91.394 12.933 92.072 12.973 ;
      RECT MASK 1 101.354 12.933 102.032 12.973 ;
      RECT MASK 1 102.184 12.933 102.862 12.973 ;
      RECT MASK 1 103.014 12.933 103.692 12.973 ;
      RECT MASK 1 103.844 12.933 104.522 12.973 ;
      RECT MASK 1 4.327 13.0225 4.507 13.0625 ;
      RECT MASK 1 111.563 13.0225 111.743 13.0625 ;
      RECT MASK 1 8.522 13.117 8.871 13.157 ;
      RECT MASK 1 9.093 13.117 9.442 13.157 ;
      RECT MASK 1 10.182 13.117 10.531 13.157 ;
      RECT MASK 1 10.753 13.117 11.102 13.157 ;
      RECT MASK 1 22.373 13.117 22.722 13.157 ;
      RECT MASK 1 23.462 13.117 23.811 13.157 ;
      RECT MASK 1 24.033 13.117 24.382 13.157 ;
      RECT MASK 1 25.122 13.117 25.471 13.157 ;
      RECT MASK 1 25.658 13.117 26.208 13.157 ;
      RECT MASK 1 26.616 13.117 27.166 13.157 ;
      RECT MASK 1 27.446 13.117 27.629 13.157 ;
      RECT MASK 1 28.276 13.117 28.826 13.157 ;
      RECT MASK 1 28.978 13.117 29.528 13.157 ;
      RECT MASK 1 30.009 13.117 30.192 13.157 ;
      RECT MASK 1 30.638 13.117 31.188 13.157 ;
      RECT MASK 1 31.596 13.117 32.146 13.157 ;
      RECT MASK 1 32.298 13.117 32.848 13.157 ;
      RECT MASK 1 33.256 13.117 33.806 13.157 ;
      RECT MASK 1 34.252 13.117 34.601 13.157 ;
      RECT MASK 1 34.823 13.117 35.172 13.157 ;
      RECT MASK 1 35.653 13.117 36.002 13.157 ;
      RECT MASK 1 36.742 13.117 37.091 13.157 ;
      RECT MASK 1 37.278 13.117 37.828 13.157 ;
      RECT MASK 1 38.236 13.117 38.786 13.157 ;
      RECT MASK 1 38.938 13.117 39.488 13.157 ;
      RECT MASK 1 39.896 13.117 40.446 13.157 ;
      RECT MASK 1 40.726 13.117 40.909 13.157 ;
      RECT MASK 1 41.556 13.117 41.739 13.157 ;
      RECT MASK 1 42.258 13.117 42.808 13.157 ;
      RECT MASK 1 43.216 13.117 43.766 13.157 ;
      RECT MASK 1 43.953 13.117 44.302 13.157 ;
      RECT MASK 1 45.042 13.117 45.391 13.157 ;
      RECT MASK 1 45.872 13.117 46.221 13.157 ;
      RECT MASK 1 46.702 13.117 47.051 13.157 ;
      RECT MASK 1 47.238 13.117 47.788 13.157 ;
      RECT MASK 1 48.196 13.117 48.746 13.157 ;
      RECT MASK 1 48.933 13.117 49.282 13.157 ;
      RECT MASK 1 50.022 13.117 50.371 13.157 ;
      RECT MASK 1 50.593 13.117 50.942 13.157 ;
      RECT MASK 1 51.682 13.117 52.031 13.157 ;
      RECT MASK 1 52.253 13.117 52.602 13.157 ;
      RECT MASK 1 53.342 13.117 53.691 13.157 ;
      RECT MASK 1 53.878 13.117 54.428 13.157 ;
      RECT MASK 1 54.836 13.117 55.386 13.157 ;
      RECT MASK 1 55.573 13.117 55.756 13.157 ;
      RECT MASK 1 56.662 13.117 57.212 13.157 ;
      RECT MASK 1 57.364 13.117 57.914 13.157 ;
      RECT MASK 1 58.488 13.117 58.837 13.157 ;
      RECT MASK 1 59.059 13.117 59.408 13.157 ;
      RECT MASK 1 60.055 13.117 60.238 13.157 ;
      RECT MASK 1 60.719 13.117 61.068 13.157 ;
      RECT MASK 1 61.808 13.117 62.157 13.157 ;
      RECT MASK 1 62.472 13.117 62.655 13.157 ;
      RECT MASK 1 63.302 13.117 63.852 13.157 ;
      RECT MASK 1 64.004 13.117 64.554 13.157 ;
      RECT MASK 1 65.128 13.117 65.477 13.157 ;
      RECT MASK 1 65.699 13.117 66.048 13.157 ;
      RECT MASK 1 66.788 13.117 67.137 13.157 ;
      RECT MASK 1 67.359 13.117 67.708 13.157 ;
      RECT MASK 1 68.448 13.117 68.797 13.157 ;
      RECT MASK 1 69.019 13.117 69.368 13.157 ;
      RECT MASK 1 70.108 13.117 70.457 13.157 ;
      RECT MASK 1 70.679 13.117 71.028 13.157 ;
      RECT MASK 1 71.768 13.117 72.117 13.157 ;
      RECT MASK 1 72.339 13.117 72.688 13.157 ;
      RECT MASK 1 77.319 13.117 77.668 13.157 ;
      RECT MASK 1 78.408 13.117 78.757 13.157 ;
      RECT MASK 1 78.979 13.117 79.328 13.157 ;
      RECT MASK 1 80.068 13.117 80.417 13.157 ;
      RECT MASK 1 83.222 13.117 83.772 13.157 ;
      RECT MASK 1 83.924 13.117 84.474 13.157 ;
      RECT MASK 1 88.939 13.117 89.288 13.157 ;
      RECT MASK 1 90.028 13.117 90.377 13.157 ;
      RECT MASK 1 90.599 13.117 90.948 13.157 ;
      RECT MASK 1 91.688 13.117 92.037 13.157 ;
      RECT MASK 1 101.648 13.117 101.997 13.157 ;
      RECT MASK 1 102.219 13.117 102.568 13.157 ;
      RECT MASK 1 103.308 13.117 103.657 13.157 ;
      RECT MASK 1 103.879 13.117 104.228 13.157 ;
      RECT MASK 1 4.251 13.284 111.819 13.324 ;
      RECT MASK 1 4.251 13.459 111.819 13.499 ;
      RECT MASK 1 4.362 13.78 111.708 13.82 ;
      RECT MASK 1 116.154 13.86 116.214 14.91 ;
      RECT MASK 1 116.428 13.86 116.488 14.91 ;
      RECT MASK 1 116.702 13.86 116.762 14.91 ;
      RECT MASK 1 116.976 13.86 117.036 14.91 ;
      RECT MASK 1 117.25 13.86 117.31 14.91 ;
      RECT MASK 1 117.524 13.86 117.584 14.91 ;
      RECT MASK 1 117.798 13.86 117.858 14.91 ;
      RECT MASK 1 118.072 13.86 118.132 14.91 ;
      RECT MASK 1 118.346 13.86 118.406 14.91 ;
      RECT MASK 1 118.62 13.86 118.68 14.91 ;
      RECT MASK 1 118.894 13.86 118.954 14.91 ;
      RECT MASK 1 119.168 13.86 119.228 14.91 ;
      RECT MASK 1 119.442 13.86 119.502 14.91 ;
      RECT MASK 1 119.716 13.86 119.776 14.91 ;
      RECT MASK 1 119.99 13.86 120.05 14.91 ;
      RECT MASK 1 120.264 13.86 120.324 14.91 ;
      RECT MASK 1 120.538 13.86 120.598 14.91 ;
      RECT MASK 1 120.812 13.86 120.872 14.91 ;
      RECT MASK 1 121.086 13.86 121.146 14.91 ;
      RECT MASK 1 121.36 13.86 121.42 14.91 ;
      RECT MASK 1 121.634 13.86 121.694 14.91 ;
      RECT MASK 1 121.908 13.86 121.968 14.91 ;
      RECT MASK 1 122.182 13.86 122.242 14.91 ;
      RECT MASK 1 122.456 13.86 122.516 14.91 ;
      RECT MASK 1 122.73 13.86 122.79 14.91 ;
      RECT MASK 1 123.004 13.86 123.064 14.91 ;
      RECT MASK 1 123.278 13.86 123.338 14.91 ;
      RECT MASK 1 123.552 13.86 123.612 14.91 ;
      RECT MASK 1 123.826 13.86 123.886 14.91 ;
      RECT MASK 1 124.1 13.86 124.16 14.91 ;
      RECT MASK 1 124.374 13.86 124.434 14.91 ;
      RECT MASK 1 124.648 13.86 124.708 14.91 ;
      RECT MASK 1 124.922 13.86 124.982 14.91 ;
      RECT MASK 1 125.196 13.86 125.256 14.91 ;
      RECT MASK 1 125.47 13.86 125.53 14.91 ;
      RECT MASK 1 125.744 13.86 125.804 14.91 ;
      RECT MASK 1 126.018 13.86 126.078 14.91 ;
      RECT MASK 1 126.292 13.86 126.352 14.91 ;
      RECT MASK 1 126.566 13.86 126.626 14.91 ;
      RECT MASK 1 126.84 13.86 126.9 14.91 ;
      RECT MASK 1 127.114 13.86 127.174 14.91 ;
      RECT MASK 1 127.388 13.86 127.448 14.91 ;
      RECT MASK 1 127.662 13.86 127.722 14.91 ;
      RECT MASK 1 127.936 13.86 127.996 14.91 ;
      RECT MASK 1 128.21 13.86 128.27 14.91 ;
      RECT MASK 1 4.251 14.101 111.819 14.141 ;
      RECT MASK 1 4.251 14.276 111.819 14.316 ;
      RECT MASK 1 5.036 14.443 5.586 14.483 ;
      RECT MASK 1 5.738 14.443 6.288 14.483 ;
      RECT MASK 1 6.696 14.443 7.246 14.483 ;
      RECT MASK 1 7.398 14.443 7.948 14.483 ;
      RECT MASK 1 8.356 14.443 8.906 14.483 ;
      RECT MASK 1 9.058 14.443 9.608 14.483 ;
      RECT MASK 1 10.016 14.443 10.566 14.483 ;
      RECT MASK 1 10.718 14.443 11.268 14.483 ;
      RECT MASK 1 11.676 14.443 12.226 14.483 ;
      RECT MASK 1 12.378 14.443 12.928 14.483 ;
      RECT MASK 1 13.336 14.443 13.886 14.483 ;
      RECT MASK 1 14.038 14.443 14.588 14.483 ;
      RECT MASK 1 14.996 14.443 15.546 14.483 ;
      RECT MASK 1 15.698 14.443 16.248 14.483 ;
      RECT MASK 1 16.656 14.443 17.206 14.483 ;
      RECT MASK 1 17.358 14.443 17.908 14.483 ;
      RECT MASK 1 18.316 14.443 18.866 14.483 ;
      RECT MASK 1 19.018 14.443 19.568 14.483 ;
      RECT MASK 1 19.976 14.443 20.526 14.483 ;
      RECT MASK 1 20.678 14.443 21.228 14.483 ;
      RECT MASK 1 21.636 14.443 22.186 14.483 ;
      RECT MASK 1 22.338 14.443 22.888 14.483 ;
      RECT MASK 1 23.296 14.443 23.846 14.483 ;
      RECT MASK 1 23.998 14.443 24.548 14.483 ;
      RECT MASK 1 24.956 14.443 25.506 14.483 ;
      RECT MASK 1 25.658 14.443 26.208 14.483 ;
      RECT MASK 1 26.616 14.443 27.166 14.483 ;
      RECT MASK 1 27.318 14.443 27.868 14.483 ;
      RECT MASK 1 28.276 14.443 28.826 14.483 ;
      RECT MASK 1 28.978 14.443 29.528 14.483 ;
      RECT MASK 1 29.936 14.443 30.486 14.483 ;
      RECT MASK 1 30.638 14.443 31.188 14.483 ;
      RECT MASK 1 31.596 14.443 32.146 14.483 ;
      RECT MASK 1 32.298 14.443 32.848 14.483 ;
      RECT MASK 1 33.256 14.443 33.806 14.483 ;
      RECT MASK 1 33.958 14.443 34.508 14.483 ;
      RECT MASK 1 34.916 14.443 35.466 14.483 ;
      RECT MASK 1 35.618 14.443 36.168 14.483 ;
      RECT MASK 1 36.576 14.443 37.126 14.483 ;
      RECT MASK 1 37.278 14.443 37.828 14.483 ;
      RECT MASK 1 38.236 14.443 38.786 14.483 ;
      RECT MASK 1 38.938 14.443 39.488 14.483 ;
      RECT MASK 1 39.896 14.443 40.446 14.483 ;
      RECT MASK 1 40.598 14.443 41.148 14.483 ;
      RECT MASK 1 41.556 14.443 42.106 14.483 ;
      RECT MASK 1 42.258 14.443 42.808 14.483 ;
      RECT MASK 1 43.216 14.443 43.766 14.483 ;
      RECT MASK 1 43.918 14.443 44.468 14.483 ;
      RECT MASK 1 44.876 14.443 45.426 14.483 ;
      RECT MASK 1 45.578 14.443 46.128 14.483 ;
      RECT MASK 1 46.536 14.443 47.086 14.483 ;
      RECT MASK 1 47.238 14.443 47.788 14.483 ;
      RECT MASK 1 48.196 14.443 48.746 14.483 ;
      RECT MASK 1 48.898 14.443 49.448 14.483 ;
      RECT MASK 1 49.856 14.443 50.406 14.483 ;
      RECT MASK 1 50.558 14.443 51.108 14.483 ;
      RECT MASK 1 51.516 14.443 52.066 14.483 ;
      RECT MASK 1 52.218 14.443 52.768 14.483 ;
      RECT MASK 1 53.176 14.443 53.726 14.483 ;
      RECT MASK 1 53.878 14.443 54.428 14.483 ;
      RECT MASK 1 54.836 14.443 55.386 14.483 ;
      RECT MASK 1 55.538 14.443 56.088 14.483 ;
      RECT MASK 1 56.662 14.443 57.212 14.483 ;
      RECT MASK 1 57.364 14.443 57.914 14.483 ;
      RECT MASK 1 58.322 14.443 58.872 14.483 ;
      RECT MASK 1 59.024 14.443 59.574 14.483 ;
      RECT MASK 1 59.982 14.443 60.532 14.483 ;
      RECT MASK 1 60.684 14.443 61.234 14.483 ;
      RECT MASK 1 61.642 14.443 62.192 14.483 ;
      RECT MASK 1 62.344 14.443 62.894 14.483 ;
      RECT MASK 1 63.302 14.443 63.852 14.483 ;
      RECT MASK 1 64.004 14.443 64.554 14.483 ;
      RECT MASK 1 64.962 14.443 65.512 14.483 ;
      RECT MASK 1 65.664 14.443 66.214 14.483 ;
      RECT MASK 1 66.622 14.443 67.172 14.483 ;
      RECT MASK 1 67.324 14.443 67.874 14.483 ;
      RECT MASK 1 68.282 14.443 68.832 14.483 ;
      RECT MASK 1 68.984 14.443 69.534 14.483 ;
      RECT MASK 1 69.942 14.443 70.492 14.483 ;
      RECT MASK 1 70.644 14.443 71.194 14.483 ;
      RECT MASK 1 71.602 14.443 72.152 14.483 ;
      RECT MASK 1 72.304 14.443 72.854 14.483 ;
      RECT MASK 1 73.262 14.443 73.812 14.483 ;
      RECT MASK 1 73.964 14.443 74.514 14.483 ;
      RECT MASK 1 74.922 14.443 75.472 14.483 ;
      RECT MASK 1 75.624 14.443 76.174 14.483 ;
      RECT MASK 1 76.582 14.443 77.132 14.483 ;
      RECT MASK 1 77.284 14.443 77.834 14.483 ;
      RECT MASK 1 78.242 14.443 78.792 14.483 ;
      RECT MASK 1 78.944 14.443 79.494 14.483 ;
      RECT MASK 1 79.902 14.443 80.452 14.483 ;
      RECT MASK 1 80.604 14.443 81.154 14.483 ;
      RECT MASK 1 81.562 14.443 82.112 14.483 ;
      RECT MASK 1 82.264 14.443 82.814 14.483 ;
      RECT MASK 1 83.222 14.443 83.772 14.483 ;
      RECT MASK 1 83.924 14.443 84.474 14.483 ;
      RECT MASK 1 84.882 14.443 85.432 14.483 ;
      RECT MASK 1 85.584 14.443 86.134 14.483 ;
      RECT MASK 1 86.542 14.443 87.092 14.483 ;
      RECT MASK 1 87.244 14.443 87.794 14.483 ;
      RECT MASK 1 88.202 14.443 88.752 14.483 ;
      RECT MASK 1 88.904 14.443 89.454 14.483 ;
      RECT MASK 1 89.862 14.443 90.412 14.483 ;
      RECT MASK 1 90.564 14.443 91.114 14.483 ;
      RECT MASK 1 91.522 14.443 92.072 14.483 ;
      RECT MASK 1 92.224 14.443 92.774 14.483 ;
      RECT MASK 1 93.182 14.443 93.732 14.483 ;
      RECT MASK 1 93.884 14.443 94.434 14.483 ;
      RECT MASK 1 94.842 14.443 95.392 14.483 ;
      RECT MASK 1 95.544 14.443 96.094 14.483 ;
      RECT MASK 1 96.502 14.443 97.052 14.483 ;
      RECT MASK 1 97.204 14.443 97.754 14.483 ;
      RECT MASK 1 98.162 14.443 98.712 14.483 ;
      RECT MASK 1 98.864 14.443 99.414 14.483 ;
      RECT MASK 1 99.822 14.443 100.372 14.483 ;
      RECT MASK 1 100.524 14.443 101.074 14.483 ;
      RECT MASK 1 101.482 14.443 102.032 14.483 ;
      RECT MASK 1 102.184 14.443 102.734 14.483 ;
      RECT MASK 1 103.142 14.443 103.692 14.483 ;
      RECT MASK 1 103.844 14.443 104.394 14.483 ;
      RECT MASK 1 104.802 14.443 105.352 14.483 ;
      RECT MASK 1 105.504 14.443 106.054 14.483 ;
      RECT MASK 1 106.462 14.443 107.012 14.483 ;
      RECT MASK 1 107.164 14.443 107.714 14.483 ;
      RECT MASK 1 108.122 14.443 108.672 14.483 ;
      RECT MASK 1 108.824 14.443 109.374 14.483 ;
      RECT MASK 1 109.782 14.443 110.332 14.483 ;
      RECT MASK 1 110.484 14.443 111.034 14.483 ;
      RECT MASK 1 4.327 14.5375 4.507 14.5775 ;
      RECT MASK 1 111.563 14.5375 111.743 14.5775 ;
      RECT MASK 1 4.908 14.627 5.586 14.667 ;
      RECT MASK 1 5.738 14.627 6.416 14.667 ;
      RECT MASK 1 6.568 14.627 7.246 14.667 ;
      RECT MASK 1 7.398 14.627 8.076 14.667 ;
      RECT MASK 1 8.228 14.627 8.906 14.667 ;
      RECT MASK 1 9.058 14.627 9.736 14.667 ;
      RECT MASK 1 9.888 14.627 10.566 14.667 ;
      RECT MASK 1 10.718 14.627 11.396 14.667 ;
      RECT MASK 1 11.548 14.627 12.226 14.667 ;
      RECT MASK 1 12.378 14.627 13.056 14.667 ;
      RECT MASK 1 13.208 14.627 13.886 14.667 ;
      RECT MASK 1 14.038 14.627 14.716 14.667 ;
      RECT MASK 1 14.868 14.627 15.546 14.667 ;
      RECT MASK 1 15.698 14.627 16.376 14.667 ;
      RECT MASK 1 16.528 14.627 17.206 14.667 ;
      RECT MASK 1 17.358 14.627 18.036 14.667 ;
      RECT MASK 1 18.188 14.627 18.866 14.667 ;
      RECT MASK 1 19.018 14.627 19.696 14.667 ;
      RECT MASK 1 19.848 14.627 20.526 14.667 ;
      RECT MASK 1 20.678 14.627 21.356 14.667 ;
      RECT MASK 1 21.508 14.627 22.186 14.667 ;
      RECT MASK 1 22.338 14.627 23.016 14.667 ;
      RECT MASK 1 23.168 14.627 23.846 14.667 ;
      RECT MASK 1 23.998 14.627 24.676 14.667 ;
      RECT MASK 1 24.828 14.627 25.506 14.667 ;
      RECT MASK 1 25.658 14.627 26.336 14.667 ;
      RECT MASK 1 26.488 14.627 27.166 14.667 ;
      RECT MASK 1 27.318 14.627 27.996 14.667 ;
      RECT MASK 1 28.148 14.627 28.826 14.667 ;
      RECT MASK 1 28.978 14.627 29.656 14.667 ;
      RECT MASK 1 29.808 14.627 30.486 14.667 ;
      RECT MASK 1 30.638 14.627 31.316 14.667 ;
      RECT MASK 1 31.468 14.627 32.146 14.667 ;
      RECT MASK 1 32.298 14.627 32.976 14.667 ;
      RECT MASK 1 33.128 14.627 33.806 14.667 ;
      RECT MASK 1 33.958 14.627 34.636 14.667 ;
      RECT MASK 1 34.788 14.627 35.466 14.667 ;
      RECT MASK 1 35.618 14.627 36.296 14.667 ;
      RECT MASK 1 36.448 14.627 37.126 14.667 ;
      RECT MASK 1 37.278 14.627 37.956 14.667 ;
      RECT MASK 1 38.108 14.627 38.786 14.667 ;
      RECT MASK 1 38.938 14.627 39.616 14.667 ;
      RECT MASK 1 39.768 14.627 40.446 14.667 ;
      RECT MASK 1 40.598 14.627 41.276 14.667 ;
      RECT MASK 1 41.428 14.627 42.106 14.667 ;
      RECT MASK 1 42.258 14.627 42.936 14.667 ;
      RECT MASK 1 43.088 14.627 43.766 14.667 ;
      RECT MASK 1 43.918 14.627 44.596 14.667 ;
      RECT MASK 1 44.748 14.627 45.426 14.667 ;
      RECT MASK 1 45.578 14.627 46.256 14.667 ;
      RECT MASK 1 46.408 14.627 47.086 14.667 ;
      RECT MASK 1 47.238 14.627 47.916 14.667 ;
      RECT MASK 1 48.068 14.627 48.746 14.667 ;
      RECT MASK 1 48.898 14.627 49.576 14.667 ;
      RECT MASK 1 49.728 14.627 50.406 14.667 ;
      RECT MASK 1 50.558 14.627 51.236 14.667 ;
      RECT MASK 1 51.388 14.627 52.066 14.667 ;
      RECT MASK 1 52.218 14.627 52.896 14.667 ;
      RECT MASK 1 53.048 14.627 53.726 14.667 ;
      RECT MASK 1 53.878 14.627 54.556 14.667 ;
      RECT MASK 1 54.708 14.627 55.386 14.667 ;
      RECT MASK 1 55.538 14.627 56.216 14.667 ;
      RECT MASK 1 56.534 14.627 57.212 14.667 ;
      RECT MASK 1 57.364 14.627 58.042 14.667 ;
      RECT MASK 1 58.194 14.627 58.872 14.667 ;
      RECT MASK 1 59.024 14.627 59.702 14.667 ;
      RECT MASK 1 59.854 14.627 60.532 14.667 ;
      RECT MASK 1 60.684 14.627 61.362 14.667 ;
      RECT MASK 1 61.514 14.627 62.192 14.667 ;
      RECT MASK 1 62.344 14.627 63.022 14.667 ;
      RECT MASK 1 63.174 14.627 63.852 14.667 ;
      RECT MASK 1 64.004 14.627 64.682 14.667 ;
      RECT MASK 1 64.834 14.627 65.512 14.667 ;
      RECT MASK 1 65.664 14.627 66.342 14.667 ;
      RECT MASK 1 66.494 14.627 67.172 14.667 ;
      RECT MASK 1 67.324 14.627 68.002 14.667 ;
      RECT MASK 1 68.154 14.627 68.832 14.667 ;
      RECT MASK 1 68.984 14.627 69.662 14.667 ;
      RECT MASK 1 69.814 14.627 70.492 14.667 ;
      RECT MASK 1 70.644 14.627 71.322 14.667 ;
      RECT MASK 1 71.474 14.627 72.152 14.667 ;
      RECT MASK 1 72.304 14.627 72.982 14.667 ;
      RECT MASK 1 73.134 14.627 73.812 14.667 ;
      RECT MASK 1 73.964 14.627 74.642 14.667 ;
      RECT MASK 1 74.794 14.627 75.472 14.667 ;
      RECT MASK 1 75.624 14.627 76.302 14.667 ;
      RECT MASK 1 76.454 14.627 77.132 14.667 ;
      RECT MASK 1 77.284 14.627 77.962 14.667 ;
      RECT MASK 1 78.114 14.627 78.792 14.667 ;
      RECT MASK 1 78.944 14.627 79.622 14.667 ;
      RECT MASK 1 79.774 14.627 80.452 14.667 ;
      RECT MASK 1 80.604 14.627 81.282 14.667 ;
      RECT MASK 1 81.434 14.627 82.112 14.667 ;
      RECT MASK 1 82.264 14.627 82.942 14.667 ;
      RECT MASK 1 83.094 14.627 83.772 14.667 ;
      RECT MASK 1 83.924 14.627 84.602 14.667 ;
      RECT MASK 1 84.754 14.627 85.432 14.667 ;
      RECT MASK 1 85.584 14.627 86.262 14.667 ;
      RECT MASK 1 86.414 14.627 87.092 14.667 ;
      RECT MASK 1 87.244 14.627 87.922 14.667 ;
      RECT MASK 1 88.074 14.627 88.752 14.667 ;
      RECT MASK 1 88.904 14.627 89.582 14.667 ;
      RECT MASK 1 89.734 14.627 90.412 14.667 ;
      RECT MASK 1 90.564 14.627 91.242 14.667 ;
      RECT MASK 1 91.394 14.627 92.072 14.667 ;
      RECT MASK 1 92.224 14.627 92.902 14.667 ;
      RECT MASK 1 93.054 14.627 93.732 14.667 ;
      RECT MASK 1 93.884 14.627 94.562 14.667 ;
      RECT MASK 1 94.714 14.627 95.392 14.667 ;
      RECT MASK 1 95.544 14.627 96.222 14.667 ;
      RECT MASK 1 96.374 14.627 97.052 14.667 ;
      RECT MASK 1 97.204 14.627 97.882 14.667 ;
      RECT MASK 1 98.034 14.627 98.712 14.667 ;
      RECT MASK 1 98.864 14.627 99.542 14.667 ;
      RECT MASK 1 99.694 14.627 100.372 14.667 ;
      RECT MASK 1 100.524 14.627 101.202 14.667 ;
      RECT MASK 1 101.354 14.627 102.032 14.667 ;
      RECT MASK 1 102.184 14.627 102.862 14.667 ;
      RECT MASK 1 103.014 14.627 103.692 14.667 ;
      RECT MASK 1 103.844 14.627 104.522 14.667 ;
      RECT MASK 1 104.674 14.627 105.352 14.667 ;
      RECT MASK 1 105.504 14.627 106.182 14.667 ;
      RECT MASK 1 106.334 14.627 107.012 14.667 ;
      RECT MASK 1 107.164 14.627 107.842 14.667 ;
      RECT MASK 1 107.994 14.627 108.672 14.667 ;
      RECT MASK 1 108.824 14.627 109.502 14.667 ;
      RECT MASK 1 109.654 14.627 110.332 14.667 ;
      RECT MASK 1 110.484 14.627 111.162 14.667 ;
      RECT MASK 1 4.908 14.853 5.586 14.893 ;
      RECT MASK 1 5.738 14.853 6.416 14.893 ;
      RECT MASK 1 6.568 14.853 7.246 14.893 ;
      RECT MASK 1 7.398 14.853 8.076 14.893 ;
      RECT MASK 1 8.228 14.853 8.906 14.893 ;
      RECT MASK 1 9.058 14.853 9.736 14.893 ;
      RECT MASK 1 9.888 14.853 10.566 14.893 ;
      RECT MASK 1 10.718 14.853 11.396 14.893 ;
      RECT MASK 1 11.548 14.853 12.226 14.893 ;
      RECT MASK 1 12.378 14.853 13.056 14.893 ;
      RECT MASK 1 13.208 14.853 13.886 14.893 ;
      RECT MASK 1 14.038 14.853 14.716 14.893 ;
      RECT MASK 1 14.868 14.853 15.546 14.893 ;
      RECT MASK 1 15.698 14.853 16.376 14.893 ;
      RECT MASK 1 16.528 14.853 17.206 14.893 ;
      RECT MASK 1 17.358 14.853 18.036 14.893 ;
      RECT MASK 1 18.188 14.853 18.866 14.893 ;
      RECT MASK 1 19.018 14.853 19.696 14.893 ;
      RECT MASK 1 19.848 14.853 20.526 14.893 ;
      RECT MASK 1 20.678 14.853 21.356 14.893 ;
      RECT MASK 1 21.508 14.853 22.186 14.893 ;
      RECT MASK 1 22.338 14.853 23.016 14.893 ;
      RECT MASK 1 23.168 14.853 23.846 14.893 ;
      RECT MASK 1 23.998 14.853 24.676 14.893 ;
      RECT MASK 1 24.828 14.853 25.506 14.893 ;
      RECT MASK 1 25.658 14.853 26.336 14.893 ;
      RECT MASK 1 26.488 14.853 27.166 14.893 ;
      RECT MASK 1 27.318 14.853 27.996 14.893 ;
      RECT MASK 1 28.148 14.853 28.826 14.893 ;
      RECT MASK 1 28.978 14.853 29.656 14.893 ;
      RECT MASK 1 29.808 14.853 30.486 14.893 ;
      RECT MASK 1 30.638 14.853 31.316 14.893 ;
      RECT MASK 1 31.468 14.853 32.146 14.893 ;
      RECT MASK 1 32.298 14.853 32.976 14.893 ;
      RECT MASK 1 33.128 14.853 33.806 14.893 ;
      RECT MASK 1 33.958 14.853 34.636 14.893 ;
      RECT MASK 1 34.788 14.853 35.466 14.893 ;
      RECT MASK 1 35.618 14.853 36.296 14.893 ;
      RECT MASK 1 36.448 14.853 37.126 14.893 ;
      RECT MASK 1 37.278 14.853 37.956 14.893 ;
      RECT MASK 1 38.108 14.853 38.786 14.893 ;
      RECT MASK 1 38.938 14.853 39.616 14.893 ;
      RECT MASK 1 39.768 14.853 40.446 14.893 ;
      RECT MASK 1 40.598 14.853 41.276 14.893 ;
      RECT MASK 1 41.428 14.853 42.106 14.893 ;
      RECT MASK 1 42.258 14.853 42.936 14.893 ;
      RECT MASK 1 43.088 14.853 43.766 14.893 ;
      RECT MASK 1 43.918 14.853 44.596 14.893 ;
      RECT MASK 1 44.748 14.853 45.426 14.893 ;
      RECT MASK 1 45.578 14.853 46.256 14.893 ;
      RECT MASK 1 46.408 14.853 47.086 14.893 ;
      RECT MASK 1 47.238 14.853 47.916 14.893 ;
      RECT MASK 1 48.068 14.853 48.746 14.893 ;
      RECT MASK 1 48.898 14.853 49.576 14.893 ;
      RECT MASK 1 49.728 14.853 50.406 14.893 ;
      RECT MASK 1 50.558 14.853 51.236 14.893 ;
      RECT MASK 1 51.388 14.853 52.066 14.893 ;
      RECT MASK 1 52.218 14.853 52.896 14.893 ;
      RECT MASK 1 53.048 14.853 53.726 14.893 ;
      RECT MASK 1 53.878 14.853 54.556 14.893 ;
      RECT MASK 1 54.708 14.853 55.386 14.893 ;
      RECT MASK 1 55.538 14.853 56.216 14.893 ;
      RECT MASK 1 56.534 14.853 57.212 14.893 ;
      RECT MASK 1 57.364 14.853 58.042 14.893 ;
      RECT MASK 1 58.194 14.853 58.872 14.893 ;
      RECT MASK 1 59.024 14.853 59.702 14.893 ;
      RECT MASK 1 59.854 14.853 60.532 14.893 ;
      RECT MASK 1 60.684 14.853 61.362 14.893 ;
      RECT MASK 1 61.514 14.853 62.192 14.893 ;
      RECT MASK 1 62.344 14.853 63.022 14.893 ;
      RECT MASK 1 63.174 14.853 63.852 14.893 ;
      RECT MASK 1 64.004 14.853 64.682 14.893 ;
      RECT MASK 1 64.834 14.853 65.512 14.893 ;
      RECT MASK 1 65.664 14.853 66.342 14.893 ;
      RECT MASK 1 66.494 14.853 67.172 14.893 ;
      RECT MASK 1 67.324 14.853 68.002 14.893 ;
      RECT MASK 1 68.154 14.853 68.832 14.893 ;
      RECT MASK 1 68.984 14.853 69.662 14.893 ;
      RECT MASK 1 69.814 14.853 70.492 14.893 ;
      RECT MASK 1 70.644 14.853 71.322 14.893 ;
      RECT MASK 1 71.474 14.853 72.152 14.893 ;
      RECT MASK 1 72.304 14.853 72.982 14.893 ;
      RECT MASK 1 73.134 14.853 73.812 14.893 ;
      RECT MASK 1 73.964 14.853 74.642 14.893 ;
      RECT MASK 1 74.794 14.853 75.472 14.893 ;
      RECT MASK 1 75.624 14.853 76.302 14.893 ;
      RECT MASK 1 76.454 14.853 77.132 14.893 ;
      RECT MASK 1 77.284 14.853 77.962 14.893 ;
      RECT MASK 1 78.114 14.853 78.792 14.893 ;
      RECT MASK 1 78.944 14.853 79.622 14.893 ;
      RECT MASK 1 79.774 14.853 80.452 14.893 ;
      RECT MASK 1 80.604 14.853 81.282 14.893 ;
      RECT MASK 1 81.434 14.853 82.112 14.893 ;
      RECT MASK 1 82.264 14.853 82.942 14.893 ;
      RECT MASK 1 83.094 14.853 83.772 14.893 ;
      RECT MASK 1 83.924 14.853 84.602 14.893 ;
      RECT MASK 1 84.754 14.853 85.432 14.893 ;
      RECT MASK 1 85.584 14.853 86.262 14.893 ;
      RECT MASK 1 86.414 14.853 87.092 14.893 ;
      RECT MASK 1 87.244 14.853 87.922 14.893 ;
      RECT MASK 1 88.074 14.853 88.752 14.893 ;
      RECT MASK 1 88.904 14.853 89.582 14.893 ;
      RECT MASK 1 89.734 14.853 90.412 14.893 ;
      RECT MASK 1 90.564 14.853 91.242 14.893 ;
      RECT MASK 1 91.394 14.853 92.072 14.893 ;
      RECT MASK 1 92.224 14.853 92.902 14.893 ;
      RECT MASK 1 93.054 14.853 93.732 14.893 ;
      RECT MASK 1 93.884 14.853 94.562 14.893 ;
      RECT MASK 1 94.714 14.853 95.392 14.893 ;
      RECT MASK 1 95.544 14.853 96.222 14.893 ;
      RECT MASK 1 96.374 14.853 97.052 14.893 ;
      RECT MASK 1 97.204 14.853 97.882 14.893 ;
      RECT MASK 1 98.034 14.853 98.712 14.893 ;
      RECT MASK 1 98.864 14.853 99.542 14.893 ;
      RECT MASK 1 99.694 14.853 100.372 14.893 ;
      RECT MASK 1 100.524 14.853 101.202 14.893 ;
      RECT MASK 1 101.354 14.853 102.032 14.893 ;
      RECT MASK 1 102.184 14.853 102.862 14.893 ;
      RECT MASK 1 103.014 14.853 103.692 14.893 ;
      RECT MASK 1 103.844 14.853 104.522 14.893 ;
      RECT MASK 1 104.674 14.853 105.352 14.893 ;
      RECT MASK 1 105.504 14.853 106.182 14.893 ;
      RECT MASK 1 106.334 14.853 107.012 14.893 ;
      RECT MASK 1 107.164 14.853 107.842 14.893 ;
      RECT MASK 1 107.994 14.853 108.672 14.893 ;
      RECT MASK 1 108.824 14.853 109.502 14.893 ;
      RECT MASK 1 109.654 14.853 110.332 14.893 ;
      RECT MASK 1 110.484 14.853 111.162 14.893 ;
      RECT MASK 1 4.327 14.9425 4.507 14.9825 ;
      RECT MASK 1 111.563 14.9425 111.743 14.9825 ;
      RECT MASK 1 5.163 15.037 5.593 15.077 ;
      RECT MASK 1 5.731 15.037 6.161 15.077 ;
      RECT MASK 1 6.823 15.037 7.253 15.077 ;
      RECT MASK 1 7.391 15.037 7.821 15.077 ;
      RECT MASK 1 8.483 15.037 8.913 15.077 ;
      RECT MASK 1 9.051 15.037 9.481 15.077 ;
      RECT MASK 1 10.143 15.037 10.573 15.077 ;
      RECT MASK 1 10.711 15.037 11.141 15.077 ;
      RECT MASK 1 11.803 15.037 12.233 15.077 ;
      RECT MASK 1 12.371 15.037 12.801 15.077 ;
      RECT MASK 1 13.463 15.037 13.893 15.077 ;
      RECT MASK 1 14.031 15.037 14.461 15.077 ;
      RECT MASK 1 15.123 15.037 15.553 15.077 ;
      RECT MASK 1 15.691 15.037 16.121 15.077 ;
      RECT MASK 1 16.783 15.037 17.213 15.077 ;
      RECT MASK 1 17.351 15.037 17.781 15.077 ;
      RECT MASK 1 18.443 15.037 18.873 15.077 ;
      RECT MASK 1 19.011 15.037 19.441 15.077 ;
      RECT MASK 1 20.103 15.037 20.533 15.077 ;
      RECT MASK 1 20.671 15.037 21.101 15.077 ;
      RECT MASK 1 21.763 15.037 22.193 15.077 ;
      RECT MASK 1 22.331 15.037 22.761 15.077 ;
      RECT MASK 1 23.423 15.037 23.853 15.077 ;
      RECT MASK 1 23.991 15.037 24.421 15.077 ;
      RECT MASK 1 25.083 15.037 25.513 15.077 ;
      RECT MASK 1 25.651 15.037 26.081 15.077 ;
      RECT MASK 1 26.743 15.037 27.173 15.077 ;
      RECT MASK 1 27.311 15.037 27.741 15.077 ;
      RECT MASK 1 28.403 15.037 28.833 15.077 ;
      RECT MASK 1 28.971 15.037 29.401 15.077 ;
      RECT MASK 1 30.063 15.037 30.493 15.077 ;
      RECT MASK 1 30.631 15.037 31.061 15.077 ;
      RECT MASK 1 31.723 15.037 32.153 15.077 ;
      RECT MASK 1 32.291 15.037 32.721 15.077 ;
      RECT MASK 1 33.383 15.037 33.813 15.077 ;
      RECT MASK 1 33.951 15.037 34.381 15.077 ;
      RECT MASK 1 35.043 15.037 35.473 15.077 ;
      RECT MASK 1 35.611 15.037 36.041 15.077 ;
      RECT MASK 1 36.703 15.037 37.133 15.077 ;
      RECT MASK 1 37.271 15.037 37.701 15.077 ;
      RECT MASK 1 38.363 15.037 38.793 15.077 ;
      RECT MASK 1 38.931 15.037 39.361 15.077 ;
      RECT MASK 1 40.023 15.037 40.453 15.077 ;
      RECT MASK 1 40.591 15.037 41.021 15.077 ;
      RECT MASK 1 41.683 15.037 42.113 15.077 ;
      RECT MASK 1 42.251 15.037 42.681 15.077 ;
      RECT MASK 1 43.343 15.037 43.773 15.077 ;
      RECT MASK 1 43.911 15.037 44.341 15.077 ;
      RECT MASK 1 45.003 15.037 45.433 15.077 ;
      RECT MASK 1 45.571 15.037 46.001 15.077 ;
      RECT MASK 1 46.663 15.037 47.093 15.077 ;
      RECT MASK 1 47.231 15.037 47.661 15.077 ;
      RECT MASK 1 48.323 15.037 48.753 15.077 ;
      RECT MASK 1 48.891 15.037 49.321 15.077 ;
      RECT MASK 1 49.983 15.037 50.413 15.077 ;
      RECT MASK 1 50.551 15.037 50.981 15.077 ;
      RECT MASK 1 51.643 15.037 52.073 15.077 ;
      RECT MASK 1 52.211 15.037 52.641 15.077 ;
      RECT MASK 1 53.303 15.037 53.733 15.077 ;
      RECT MASK 1 53.871 15.037 54.301 15.077 ;
      RECT MASK 1 54.963 15.037 55.393 15.077 ;
      RECT MASK 1 55.531 15.037 55.961 15.077 ;
      RECT MASK 1 56.789 15.037 57.219 15.077 ;
      RECT MASK 1 57.357 15.037 57.787 15.077 ;
      RECT MASK 1 58.449 15.037 58.879 15.077 ;
      RECT MASK 1 59.017 15.037 59.447 15.077 ;
      RECT MASK 1 60.109 15.037 60.539 15.077 ;
      RECT MASK 1 60.677 15.037 61.107 15.077 ;
      RECT MASK 1 61.769 15.037 62.199 15.077 ;
      RECT MASK 1 62.337 15.037 62.767 15.077 ;
      RECT MASK 1 63.429 15.037 63.859 15.077 ;
      RECT MASK 1 63.997 15.037 64.427 15.077 ;
      RECT MASK 1 65.089 15.037 65.519 15.077 ;
      RECT MASK 1 65.657 15.037 66.087 15.077 ;
      RECT MASK 1 66.749 15.037 67.179 15.077 ;
      RECT MASK 1 67.317 15.037 67.747 15.077 ;
      RECT MASK 1 68.409 15.037 68.839 15.077 ;
      RECT MASK 1 68.977 15.037 69.407 15.077 ;
      RECT MASK 1 70.069 15.037 70.499 15.077 ;
      RECT MASK 1 70.637 15.037 71.067 15.077 ;
      RECT MASK 1 71.729 15.037 72.159 15.077 ;
      RECT MASK 1 72.297 15.037 72.727 15.077 ;
      RECT MASK 1 73.389 15.037 73.819 15.077 ;
      RECT MASK 1 73.957 15.037 74.387 15.077 ;
      RECT MASK 1 75.049 15.037 75.479 15.077 ;
      RECT MASK 1 75.617 15.037 76.047 15.077 ;
      RECT MASK 1 76.709 15.037 77.139 15.077 ;
      RECT MASK 1 77.277 15.037 77.707 15.077 ;
      RECT MASK 1 78.369 15.037 78.799 15.077 ;
      RECT MASK 1 78.937 15.037 79.367 15.077 ;
      RECT MASK 1 80.029 15.037 80.459 15.077 ;
      RECT MASK 1 80.597 15.037 81.027 15.077 ;
      RECT MASK 1 81.689 15.037 82.119 15.077 ;
      RECT MASK 1 82.257 15.037 82.687 15.077 ;
      RECT MASK 1 83.349 15.037 83.779 15.077 ;
      RECT MASK 1 83.917 15.037 84.347 15.077 ;
      RECT MASK 1 85.009 15.037 85.439 15.077 ;
      RECT MASK 1 85.577 15.037 86.007 15.077 ;
      RECT MASK 1 86.669 15.037 87.099 15.077 ;
      RECT MASK 1 87.237 15.037 87.667 15.077 ;
      RECT MASK 1 88.329 15.037 88.759 15.077 ;
      RECT MASK 1 88.897 15.037 89.327 15.077 ;
      RECT MASK 1 89.989 15.037 90.419 15.077 ;
      RECT MASK 1 90.557 15.037 90.987 15.077 ;
      RECT MASK 1 91.649 15.037 92.079 15.077 ;
      RECT MASK 1 92.217 15.037 92.647 15.077 ;
      RECT MASK 1 93.309 15.037 93.739 15.077 ;
      RECT MASK 1 93.877 15.037 94.307 15.077 ;
      RECT MASK 1 94.969 15.037 95.399 15.077 ;
      RECT MASK 1 95.537 15.037 95.967 15.077 ;
      RECT MASK 1 96.629 15.037 97.059 15.077 ;
      RECT MASK 1 97.197 15.037 97.627 15.077 ;
      RECT MASK 1 98.289 15.037 98.719 15.077 ;
      RECT MASK 1 98.857 15.037 99.287 15.077 ;
      RECT MASK 1 99.949 15.037 100.379 15.077 ;
      RECT MASK 1 100.517 15.037 100.947 15.077 ;
      RECT MASK 1 101.609 15.037 102.039 15.077 ;
      RECT MASK 1 102.177 15.037 102.607 15.077 ;
      RECT MASK 1 103.269 15.037 103.699 15.077 ;
      RECT MASK 1 103.837 15.037 104.267 15.077 ;
      RECT MASK 1 104.929 15.037 105.359 15.077 ;
      RECT MASK 1 105.497 15.037 105.927 15.077 ;
      RECT MASK 1 106.589 15.037 107.019 15.077 ;
      RECT MASK 1 107.157 15.037 107.587 15.077 ;
      RECT MASK 1 108.249 15.037 108.679 15.077 ;
      RECT MASK 1 108.817 15.037 109.247 15.077 ;
      RECT MASK 1 109.909 15.037 110.339 15.077 ;
      RECT MASK 1 110.477 15.037 110.907 15.077 ;
      RECT MASK 1 4.251 15.204 111.819 15.244 ;
      RECT MASK 1 4.251 15.379 111.819 15.419 ;
      RECT MASK 1 116.154 15.57 116.214 16.62 ;
      RECT MASK 1 116.428 15.57 116.488 16.62 ;
      RECT MASK 1 116.702 15.57 116.762 16.62 ;
      RECT MASK 1 116.976 15.57 117.036 16.62 ;
      RECT MASK 1 117.25 15.57 117.31 16.62 ;
      RECT MASK 1 117.524 15.57 117.584 16.62 ;
      RECT MASK 1 117.798 15.57 117.858 16.62 ;
      RECT MASK 1 118.072 15.57 118.132 16.62 ;
      RECT MASK 1 118.346 15.57 118.406 16.62 ;
      RECT MASK 1 118.62 15.57 118.68 16.62 ;
      RECT MASK 1 118.894 15.57 118.954 16.62 ;
      RECT MASK 1 119.168 15.57 119.228 16.62 ;
      RECT MASK 1 119.442 15.57 119.502 16.62 ;
      RECT MASK 1 119.716 15.57 119.776 16.62 ;
      RECT MASK 1 119.99 15.57 120.05 16.62 ;
      RECT MASK 1 120.264 15.57 120.324 16.62 ;
      RECT MASK 1 120.538 15.57 120.598 16.62 ;
      RECT MASK 1 120.812 15.57 120.872 16.62 ;
      RECT MASK 1 121.086 15.57 121.146 16.62 ;
      RECT MASK 1 121.36 15.57 121.42 16.62 ;
      RECT MASK 1 121.634 15.57 121.694 16.62 ;
      RECT MASK 1 121.908 15.57 121.968 16.62 ;
      RECT MASK 1 122.182 15.57 122.242 16.62 ;
      RECT MASK 1 122.456 15.57 122.516 16.62 ;
      RECT MASK 1 122.73 15.57 122.79 16.62 ;
      RECT MASK 1 123.004 15.57 123.064 16.62 ;
      RECT MASK 1 123.278 15.57 123.338 16.62 ;
      RECT MASK 1 123.552 15.57 123.612 16.62 ;
      RECT MASK 1 123.826 15.57 123.886 16.62 ;
      RECT MASK 1 124.1 15.57 124.16 16.62 ;
      RECT MASK 1 124.374 15.57 124.434 16.62 ;
      RECT MASK 1 124.648 15.57 124.708 16.62 ;
      RECT MASK 1 124.922 15.57 124.982 16.62 ;
      RECT MASK 1 125.196 15.57 125.256 16.62 ;
      RECT MASK 1 125.47 15.57 125.53 16.62 ;
      RECT MASK 1 125.744 15.57 125.804 16.62 ;
      RECT MASK 1 126.018 15.57 126.078 16.62 ;
      RECT MASK 1 126.292 15.57 126.352 16.62 ;
      RECT MASK 1 126.566 15.57 126.626 16.62 ;
      RECT MASK 1 126.84 15.57 126.9 16.62 ;
      RECT MASK 1 127.114 15.57 127.174 16.62 ;
      RECT MASK 1 127.388 15.57 127.448 16.62 ;
      RECT MASK 1 127.662 15.57 127.722 16.62 ;
      RECT MASK 1 127.936 15.57 127.996 16.62 ;
      RECT MASK 1 128.21 15.57 128.27 16.62 ;
      RECT MASK 1 4.362 15.7 111.708 15.74 ;
      RECT MASK 1 4.251 16.021 111.819 16.061 ;
      RECT MASK 1 4.251 16.196 111.819 16.236 ;
      RECT MASK 1 5.163 16.363 5.593 16.403 ;
      RECT MASK 1 5.731 16.363 6.161 16.403 ;
      RECT MASK 1 6.823 16.363 7.253 16.403 ;
      RECT MASK 1 7.391 16.363 7.821 16.403 ;
      RECT MASK 1 8.483 16.363 8.913 16.403 ;
      RECT MASK 1 9.051 16.363 9.481 16.403 ;
      RECT MASK 1 10.143 16.363 10.573 16.403 ;
      RECT MASK 1 10.711 16.363 11.141 16.403 ;
      RECT MASK 1 11.803 16.363 12.233 16.403 ;
      RECT MASK 1 12.371 16.363 12.801 16.403 ;
      RECT MASK 1 13.463 16.363 13.893 16.403 ;
      RECT MASK 1 14.031 16.363 14.461 16.403 ;
      RECT MASK 1 15.123 16.363 15.553 16.403 ;
      RECT MASK 1 15.691 16.363 16.121 16.403 ;
      RECT MASK 1 16.783 16.363 17.213 16.403 ;
      RECT MASK 1 17.351 16.363 17.781 16.403 ;
      RECT MASK 1 18.443 16.363 18.873 16.403 ;
      RECT MASK 1 19.011 16.363 19.441 16.403 ;
      RECT MASK 1 20.103 16.363 20.533 16.403 ;
      RECT MASK 1 20.671 16.363 21.101 16.403 ;
      RECT MASK 1 21.763 16.363 22.193 16.403 ;
      RECT MASK 1 22.331 16.363 22.761 16.403 ;
      RECT MASK 1 23.423 16.363 23.853 16.403 ;
      RECT MASK 1 23.991 16.363 24.421 16.403 ;
      RECT MASK 1 25.083 16.363 25.513 16.403 ;
      RECT MASK 1 25.651 16.363 26.081 16.403 ;
      RECT MASK 1 26.743 16.363 27.173 16.403 ;
      RECT MASK 1 27.311 16.363 27.741 16.403 ;
      RECT MASK 1 28.403 16.363 28.833 16.403 ;
      RECT MASK 1 28.971 16.363 29.401 16.403 ;
      RECT MASK 1 30.063 16.363 30.493 16.403 ;
      RECT MASK 1 30.631 16.363 31.061 16.403 ;
      RECT MASK 1 31.723 16.363 32.153 16.403 ;
      RECT MASK 1 32.291 16.363 32.721 16.403 ;
      RECT MASK 1 33.383 16.363 33.813 16.403 ;
      RECT MASK 1 33.951 16.363 34.381 16.403 ;
      RECT MASK 1 35.043 16.363 35.473 16.403 ;
      RECT MASK 1 35.611 16.363 36.041 16.403 ;
      RECT MASK 1 36.703 16.363 37.133 16.403 ;
      RECT MASK 1 37.271 16.363 37.701 16.403 ;
      RECT MASK 1 38.363 16.363 38.793 16.403 ;
      RECT MASK 1 38.931 16.363 39.361 16.403 ;
      RECT MASK 1 40.023 16.363 40.453 16.403 ;
      RECT MASK 1 40.591 16.363 41.021 16.403 ;
      RECT MASK 1 41.683 16.363 42.113 16.403 ;
      RECT MASK 1 42.251 16.363 42.681 16.403 ;
      RECT MASK 1 43.343 16.363 43.773 16.403 ;
      RECT MASK 1 43.911 16.363 44.341 16.403 ;
      RECT MASK 1 45.003 16.363 45.433 16.403 ;
      RECT MASK 1 45.571 16.363 46.001 16.403 ;
      RECT MASK 1 46.663 16.363 47.093 16.403 ;
      RECT MASK 1 47.231 16.363 47.661 16.403 ;
      RECT MASK 1 48.323 16.363 48.753 16.403 ;
      RECT MASK 1 48.891 16.363 49.321 16.403 ;
      RECT MASK 1 49.983 16.363 50.413 16.403 ;
      RECT MASK 1 50.551 16.363 50.981 16.403 ;
      RECT MASK 1 51.643 16.363 52.073 16.403 ;
      RECT MASK 1 52.211 16.363 52.641 16.403 ;
      RECT MASK 1 53.303 16.363 53.733 16.403 ;
      RECT MASK 1 53.871 16.363 54.301 16.403 ;
      RECT MASK 1 54.963 16.363 55.393 16.403 ;
      RECT MASK 1 55.531 16.363 55.961 16.403 ;
      RECT MASK 1 56.789 16.363 57.219 16.403 ;
      RECT MASK 1 57.357 16.363 57.787 16.403 ;
      RECT MASK 1 58.449 16.363 58.879 16.403 ;
      RECT MASK 1 59.017 16.363 59.447 16.403 ;
      RECT MASK 1 60.109 16.363 60.539 16.403 ;
      RECT MASK 1 60.677 16.363 61.107 16.403 ;
      RECT MASK 1 61.769 16.363 62.199 16.403 ;
      RECT MASK 1 62.337 16.363 62.767 16.403 ;
      RECT MASK 1 63.429 16.363 63.859 16.403 ;
      RECT MASK 1 63.997 16.363 64.427 16.403 ;
      RECT MASK 1 65.089 16.363 65.519 16.403 ;
      RECT MASK 1 65.657 16.363 66.087 16.403 ;
      RECT MASK 1 66.749 16.363 67.179 16.403 ;
      RECT MASK 1 67.317 16.363 67.747 16.403 ;
      RECT MASK 1 68.409 16.363 68.839 16.403 ;
      RECT MASK 1 68.977 16.363 69.407 16.403 ;
      RECT MASK 1 70.069 16.363 70.499 16.403 ;
      RECT MASK 1 70.637 16.363 71.067 16.403 ;
      RECT MASK 1 71.729 16.363 72.159 16.403 ;
      RECT MASK 1 72.297 16.363 72.727 16.403 ;
      RECT MASK 1 73.389 16.363 73.819 16.403 ;
      RECT MASK 1 73.957 16.363 74.387 16.403 ;
      RECT MASK 1 75.049 16.363 75.479 16.403 ;
      RECT MASK 1 75.617 16.363 76.047 16.403 ;
      RECT MASK 1 76.709 16.363 77.139 16.403 ;
      RECT MASK 1 77.277 16.363 77.707 16.403 ;
      RECT MASK 1 78.369 16.363 78.799 16.403 ;
      RECT MASK 1 78.937 16.363 79.367 16.403 ;
      RECT MASK 1 80.029 16.363 80.459 16.403 ;
      RECT MASK 1 80.597 16.363 81.027 16.403 ;
      RECT MASK 1 81.689 16.363 82.119 16.403 ;
      RECT MASK 1 82.257 16.363 82.687 16.403 ;
      RECT MASK 1 83.349 16.363 83.779 16.403 ;
      RECT MASK 1 83.917 16.363 84.347 16.403 ;
      RECT MASK 1 85.009 16.363 85.439 16.403 ;
      RECT MASK 1 85.577 16.363 86.007 16.403 ;
      RECT MASK 1 86.669 16.363 87.099 16.403 ;
      RECT MASK 1 87.237 16.363 87.667 16.403 ;
      RECT MASK 1 88.329 16.363 88.759 16.403 ;
      RECT MASK 1 88.897 16.363 89.327 16.403 ;
      RECT MASK 1 89.989 16.363 90.419 16.403 ;
      RECT MASK 1 90.557 16.363 90.987 16.403 ;
      RECT MASK 1 91.649 16.363 92.079 16.403 ;
      RECT MASK 1 92.217 16.363 92.647 16.403 ;
      RECT MASK 1 93.309 16.363 93.739 16.403 ;
      RECT MASK 1 93.877 16.363 94.307 16.403 ;
      RECT MASK 1 94.969 16.363 95.399 16.403 ;
      RECT MASK 1 95.537 16.363 95.967 16.403 ;
      RECT MASK 1 96.629 16.363 97.059 16.403 ;
      RECT MASK 1 97.197 16.363 97.627 16.403 ;
      RECT MASK 1 98.289 16.363 98.719 16.403 ;
      RECT MASK 1 98.857 16.363 99.287 16.403 ;
      RECT MASK 1 99.949 16.363 100.379 16.403 ;
      RECT MASK 1 100.517 16.363 100.947 16.403 ;
      RECT MASK 1 101.609 16.363 102.039 16.403 ;
      RECT MASK 1 102.177 16.363 102.607 16.403 ;
      RECT MASK 1 103.269 16.363 103.699 16.403 ;
      RECT MASK 1 103.837 16.363 104.267 16.403 ;
      RECT MASK 1 104.929 16.363 105.359 16.403 ;
      RECT MASK 1 105.497 16.363 105.927 16.403 ;
      RECT MASK 1 106.589 16.363 107.019 16.403 ;
      RECT MASK 1 107.157 16.363 107.587 16.403 ;
      RECT MASK 1 108.249 16.363 108.679 16.403 ;
      RECT MASK 1 108.817 16.363 109.247 16.403 ;
      RECT MASK 1 109.909 16.363 110.339 16.403 ;
      RECT MASK 1 110.477 16.363 110.907 16.403 ;
      RECT MASK 1 4.327 16.4575 4.507 16.4975 ;
      RECT MASK 1 111.563 16.4575 111.743 16.4975 ;
      RECT MASK 1 4.908 16.547 5.586 16.587 ;
      RECT MASK 1 5.738 16.547 6.416 16.587 ;
      RECT MASK 1 6.568 16.547 7.246 16.587 ;
      RECT MASK 1 7.398 16.547 8.076 16.587 ;
      RECT MASK 1 8.228 16.547 8.906 16.587 ;
      RECT MASK 1 9.058 16.547 9.736 16.587 ;
      RECT MASK 1 9.888 16.547 10.566 16.587 ;
      RECT MASK 1 10.718 16.547 11.396 16.587 ;
      RECT MASK 1 11.548 16.547 12.226 16.587 ;
      RECT MASK 1 12.378 16.547 13.056 16.587 ;
      RECT MASK 1 13.208 16.547 13.886 16.587 ;
      RECT MASK 1 14.038 16.547 14.716 16.587 ;
      RECT MASK 1 14.868 16.547 15.546 16.587 ;
      RECT MASK 1 15.698 16.547 16.376 16.587 ;
      RECT MASK 1 16.528 16.547 17.206 16.587 ;
      RECT MASK 1 17.358 16.547 18.036 16.587 ;
      RECT MASK 1 18.188 16.547 18.866 16.587 ;
      RECT MASK 1 19.018 16.547 19.696 16.587 ;
      RECT MASK 1 19.848 16.547 20.526 16.587 ;
      RECT MASK 1 20.678 16.547 21.356 16.587 ;
      RECT MASK 1 21.508 16.547 22.186 16.587 ;
      RECT MASK 1 22.338 16.547 23.016 16.587 ;
      RECT MASK 1 23.168 16.547 23.846 16.587 ;
      RECT MASK 1 23.998 16.547 24.676 16.587 ;
      RECT MASK 1 24.828 16.547 25.506 16.587 ;
      RECT MASK 1 25.658 16.547 26.336 16.587 ;
      RECT MASK 1 26.488 16.547 27.166 16.587 ;
      RECT MASK 1 27.318 16.547 27.996 16.587 ;
      RECT MASK 1 28.148 16.547 28.826 16.587 ;
      RECT MASK 1 28.978 16.547 29.656 16.587 ;
      RECT MASK 1 29.808 16.547 30.486 16.587 ;
      RECT MASK 1 30.638 16.547 31.316 16.587 ;
      RECT MASK 1 31.468 16.547 32.146 16.587 ;
      RECT MASK 1 32.298 16.547 32.976 16.587 ;
      RECT MASK 1 33.128 16.547 33.806 16.587 ;
      RECT MASK 1 33.958 16.547 34.636 16.587 ;
      RECT MASK 1 34.788 16.547 35.466 16.587 ;
      RECT MASK 1 35.618 16.547 36.296 16.587 ;
      RECT MASK 1 36.448 16.547 37.126 16.587 ;
      RECT MASK 1 37.278 16.547 37.956 16.587 ;
      RECT MASK 1 38.108 16.547 38.786 16.587 ;
      RECT MASK 1 38.938 16.547 39.616 16.587 ;
      RECT MASK 1 39.768 16.547 40.446 16.587 ;
      RECT MASK 1 40.598 16.547 41.276 16.587 ;
      RECT MASK 1 41.428 16.547 42.106 16.587 ;
      RECT MASK 1 42.258 16.547 42.936 16.587 ;
      RECT MASK 1 43.088 16.547 43.766 16.587 ;
      RECT MASK 1 43.918 16.547 44.596 16.587 ;
      RECT MASK 1 44.748 16.547 45.426 16.587 ;
      RECT MASK 1 45.578 16.547 46.256 16.587 ;
      RECT MASK 1 46.408 16.547 47.086 16.587 ;
      RECT MASK 1 47.238 16.547 47.916 16.587 ;
      RECT MASK 1 48.068 16.547 48.746 16.587 ;
      RECT MASK 1 48.898 16.547 49.576 16.587 ;
      RECT MASK 1 49.728 16.547 50.406 16.587 ;
      RECT MASK 1 50.558 16.547 51.236 16.587 ;
      RECT MASK 1 51.388 16.547 52.066 16.587 ;
      RECT MASK 1 52.218 16.547 52.896 16.587 ;
      RECT MASK 1 53.048 16.547 53.726 16.587 ;
      RECT MASK 1 53.878 16.547 54.556 16.587 ;
      RECT MASK 1 54.708 16.547 55.386 16.587 ;
      RECT MASK 1 55.538 16.547 56.216 16.587 ;
      RECT MASK 1 56.534 16.547 57.212 16.587 ;
      RECT MASK 1 57.364 16.547 58.042 16.587 ;
      RECT MASK 1 58.194 16.547 58.872 16.587 ;
      RECT MASK 1 59.024 16.547 59.702 16.587 ;
      RECT MASK 1 59.854 16.547 60.532 16.587 ;
      RECT MASK 1 60.684 16.547 61.362 16.587 ;
      RECT MASK 1 61.514 16.547 62.192 16.587 ;
      RECT MASK 1 62.344 16.547 63.022 16.587 ;
      RECT MASK 1 63.174 16.547 63.852 16.587 ;
      RECT MASK 1 64.004 16.547 64.682 16.587 ;
      RECT MASK 1 64.834 16.547 65.512 16.587 ;
      RECT MASK 1 65.664 16.547 66.342 16.587 ;
      RECT MASK 1 66.494 16.547 67.172 16.587 ;
      RECT MASK 1 67.324 16.547 68.002 16.587 ;
      RECT MASK 1 68.154 16.547 68.832 16.587 ;
      RECT MASK 1 68.984 16.547 69.662 16.587 ;
      RECT MASK 1 69.814 16.547 70.492 16.587 ;
      RECT MASK 1 70.644 16.547 71.322 16.587 ;
      RECT MASK 1 71.474 16.547 72.152 16.587 ;
      RECT MASK 1 72.304 16.547 72.982 16.587 ;
      RECT MASK 1 73.134 16.547 73.812 16.587 ;
      RECT MASK 1 73.964 16.547 74.642 16.587 ;
      RECT MASK 1 74.794 16.547 75.472 16.587 ;
      RECT MASK 1 75.624 16.547 76.302 16.587 ;
      RECT MASK 1 76.454 16.547 77.132 16.587 ;
      RECT MASK 1 77.284 16.547 77.962 16.587 ;
      RECT MASK 1 78.114 16.547 78.792 16.587 ;
      RECT MASK 1 78.944 16.547 79.622 16.587 ;
      RECT MASK 1 79.774 16.547 80.452 16.587 ;
      RECT MASK 1 80.604 16.547 81.282 16.587 ;
      RECT MASK 1 81.434 16.547 82.112 16.587 ;
      RECT MASK 1 82.264 16.547 82.942 16.587 ;
      RECT MASK 1 83.094 16.547 83.772 16.587 ;
      RECT MASK 1 83.924 16.547 84.602 16.587 ;
      RECT MASK 1 84.754 16.547 85.432 16.587 ;
      RECT MASK 1 85.584 16.547 86.262 16.587 ;
      RECT MASK 1 86.414 16.547 87.092 16.587 ;
      RECT MASK 1 87.244 16.547 87.922 16.587 ;
      RECT MASK 1 88.074 16.547 88.752 16.587 ;
      RECT MASK 1 88.904 16.547 89.582 16.587 ;
      RECT MASK 1 89.734 16.547 90.412 16.587 ;
      RECT MASK 1 90.564 16.547 91.242 16.587 ;
      RECT MASK 1 91.394 16.547 92.072 16.587 ;
      RECT MASK 1 92.224 16.547 92.902 16.587 ;
      RECT MASK 1 93.054 16.547 93.732 16.587 ;
      RECT MASK 1 93.884 16.547 94.562 16.587 ;
      RECT MASK 1 94.714 16.547 95.392 16.587 ;
      RECT MASK 1 95.544 16.547 96.222 16.587 ;
      RECT MASK 1 96.374 16.547 97.052 16.587 ;
      RECT MASK 1 97.204 16.547 97.882 16.587 ;
      RECT MASK 1 98.034 16.547 98.712 16.587 ;
      RECT MASK 1 98.864 16.547 99.542 16.587 ;
      RECT MASK 1 99.694 16.547 100.372 16.587 ;
      RECT MASK 1 100.524 16.547 101.202 16.587 ;
      RECT MASK 1 101.354 16.547 102.032 16.587 ;
      RECT MASK 1 102.184 16.547 102.862 16.587 ;
      RECT MASK 1 103.014 16.547 103.692 16.587 ;
      RECT MASK 1 103.844 16.547 104.522 16.587 ;
      RECT MASK 1 104.674 16.547 105.352 16.587 ;
      RECT MASK 1 105.504 16.547 106.182 16.587 ;
      RECT MASK 1 106.334 16.547 107.012 16.587 ;
      RECT MASK 1 107.164 16.547 107.842 16.587 ;
      RECT MASK 1 107.994 16.547 108.672 16.587 ;
      RECT MASK 1 108.824 16.547 109.502 16.587 ;
      RECT MASK 1 109.654 16.547 110.332 16.587 ;
      RECT MASK 1 110.484 16.547 111.162 16.587 ;
      RECT MASK 1 4.908 16.773 5.586 16.813 ;
      RECT MASK 1 5.738 16.773 6.416 16.813 ;
      RECT MASK 1 6.568 16.773 7.246 16.813 ;
      RECT MASK 1 7.398 16.773 8.076 16.813 ;
      RECT MASK 1 8.228 16.773 8.906 16.813 ;
      RECT MASK 1 9.058 16.773 9.736 16.813 ;
      RECT MASK 1 9.888 16.773 10.566 16.813 ;
      RECT MASK 1 10.718 16.773 11.396 16.813 ;
      RECT MASK 1 11.548 16.773 12.226 16.813 ;
      RECT MASK 1 12.378 16.773 13.056 16.813 ;
      RECT MASK 1 13.208 16.773 13.886 16.813 ;
      RECT MASK 1 14.038 16.773 14.716 16.813 ;
      RECT MASK 1 14.868 16.773 15.546 16.813 ;
      RECT MASK 1 15.698 16.773 16.376 16.813 ;
      RECT MASK 1 16.528 16.773 17.206 16.813 ;
      RECT MASK 1 17.358 16.773 18.036 16.813 ;
      RECT MASK 1 18.188 16.773 18.866 16.813 ;
      RECT MASK 1 19.018 16.773 19.696 16.813 ;
      RECT MASK 1 19.848 16.773 20.526 16.813 ;
      RECT MASK 1 20.678 16.773 21.356 16.813 ;
      RECT MASK 1 21.508 16.773 22.186 16.813 ;
      RECT MASK 1 22.338 16.773 23.016 16.813 ;
      RECT MASK 1 23.168 16.773 23.846 16.813 ;
      RECT MASK 1 23.998 16.773 24.676 16.813 ;
      RECT MASK 1 24.828 16.773 25.506 16.813 ;
      RECT MASK 1 25.658 16.773 26.336 16.813 ;
      RECT MASK 1 26.488 16.773 27.166 16.813 ;
      RECT MASK 1 27.318 16.773 27.996 16.813 ;
      RECT MASK 1 28.148 16.773 28.826 16.813 ;
      RECT MASK 1 28.978 16.773 29.656 16.813 ;
      RECT MASK 1 29.808 16.773 30.486 16.813 ;
      RECT MASK 1 30.638 16.773 31.316 16.813 ;
      RECT MASK 1 31.468 16.773 32.146 16.813 ;
      RECT MASK 1 32.298 16.773 32.976 16.813 ;
      RECT MASK 1 33.128 16.773 33.806 16.813 ;
      RECT MASK 1 33.958 16.773 34.636 16.813 ;
      RECT MASK 1 34.788 16.773 35.466 16.813 ;
      RECT MASK 1 35.618 16.773 36.296 16.813 ;
      RECT MASK 1 36.448 16.773 37.126 16.813 ;
      RECT MASK 1 37.278 16.773 37.956 16.813 ;
      RECT MASK 1 38.108 16.773 38.786 16.813 ;
      RECT MASK 1 38.938 16.773 39.616 16.813 ;
      RECT MASK 1 39.768 16.773 40.446 16.813 ;
      RECT MASK 1 40.598 16.773 41.276 16.813 ;
      RECT MASK 1 41.428 16.773 42.106 16.813 ;
      RECT MASK 1 42.258 16.773 42.936 16.813 ;
      RECT MASK 1 43.088 16.773 43.766 16.813 ;
      RECT MASK 1 43.918 16.773 44.596 16.813 ;
      RECT MASK 1 44.748 16.773 45.426 16.813 ;
      RECT MASK 1 45.578 16.773 46.256 16.813 ;
      RECT MASK 1 46.408 16.773 47.086 16.813 ;
      RECT MASK 1 47.238 16.773 47.916 16.813 ;
      RECT MASK 1 48.068 16.773 48.746 16.813 ;
      RECT MASK 1 48.898 16.773 49.576 16.813 ;
      RECT MASK 1 49.728 16.773 50.406 16.813 ;
      RECT MASK 1 50.558 16.773 51.236 16.813 ;
      RECT MASK 1 51.388 16.773 52.066 16.813 ;
      RECT MASK 1 52.218 16.773 52.896 16.813 ;
      RECT MASK 1 53.048 16.773 53.726 16.813 ;
      RECT MASK 1 53.878 16.773 54.556 16.813 ;
      RECT MASK 1 54.708 16.773 55.386 16.813 ;
      RECT MASK 1 55.538 16.773 56.216 16.813 ;
      RECT MASK 1 56.534 16.773 57.212 16.813 ;
      RECT MASK 1 57.364 16.773 58.042 16.813 ;
      RECT MASK 1 58.194 16.773 58.872 16.813 ;
      RECT MASK 1 59.024 16.773 59.702 16.813 ;
      RECT MASK 1 59.854 16.773 60.532 16.813 ;
      RECT MASK 1 60.684 16.773 61.362 16.813 ;
      RECT MASK 1 61.514 16.773 62.192 16.813 ;
      RECT MASK 1 62.344 16.773 63.022 16.813 ;
      RECT MASK 1 63.174 16.773 63.852 16.813 ;
      RECT MASK 1 64.004 16.773 64.682 16.813 ;
      RECT MASK 1 64.834 16.773 65.512 16.813 ;
      RECT MASK 1 65.664 16.773 66.342 16.813 ;
      RECT MASK 1 66.494 16.773 67.172 16.813 ;
      RECT MASK 1 67.324 16.773 68.002 16.813 ;
      RECT MASK 1 68.154 16.773 68.832 16.813 ;
      RECT MASK 1 68.984 16.773 69.662 16.813 ;
      RECT MASK 1 69.814 16.773 70.492 16.813 ;
      RECT MASK 1 70.644 16.773 71.322 16.813 ;
      RECT MASK 1 71.474 16.773 72.152 16.813 ;
      RECT MASK 1 72.304 16.773 72.982 16.813 ;
      RECT MASK 1 73.134 16.773 73.812 16.813 ;
      RECT MASK 1 73.964 16.773 74.642 16.813 ;
      RECT MASK 1 74.794 16.773 75.472 16.813 ;
      RECT MASK 1 75.624 16.773 76.302 16.813 ;
      RECT MASK 1 76.454 16.773 77.132 16.813 ;
      RECT MASK 1 77.284 16.773 77.962 16.813 ;
      RECT MASK 1 78.114 16.773 78.792 16.813 ;
      RECT MASK 1 78.944 16.773 79.622 16.813 ;
      RECT MASK 1 79.774 16.773 80.452 16.813 ;
      RECT MASK 1 80.604 16.773 81.282 16.813 ;
      RECT MASK 1 81.434 16.773 82.112 16.813 ;
      RECT MASK 1 82.264 16.773 82.942 16.813 ;
      RECT MASK 1 83.094 16.773 83.772 16.813 ;
      RECT MASK 1 83.924 16.773 84.602 16.813 ;
      RECT MASK 1 84.754 16.773 85.432 16.813 ;
      RECT MASK 1 85.584 16.773 86.262 16.813 ;
      RECT MASK 1 86.414 16.773 87.092 16.813 ;
      RECT MASK 1 87.244 16.773 87.922 16.813 ;
      RECT MASK 1 88.074 16.773 88.752 16.813 ;
      RECT MASK 1 88.904 16.773 89.582 16.813 ;
      RECT MASK 1 89.734 16.773 90.412 16.813 ;
      RECT MASK 1 90.564 16.773 91.242 16.813 ;
      RECT MASK 1 91.394 16.773 92.072 16.813 ;
      RECT MASK 1 92.224 16.773 92.902 16.813 ;
      RECT MASK 1 93.054 16.773 93.732 16.813 ;
      RECT MASK 1 93.884 16.773 94.562 16.813 ;
      RECT MASK 1 94.714 16.773 95.392 16.813 ;
      RECT MASK 1 95.544 16.773 96.222 16.813 ;
      RECT MASK 1 96.374 16.773 97.052 16.813 ;
      RECT MASK 1 97.204 16.773 97.882 16.813 ;
      RECT MASK 1 98.034 16.773 98.712 16.813 ;
      RECT MASK 1 98.864 16.773 99.542 16.813 ;
      RECT MASK 1 99.694 16.773 100.372 16.813 ;
      RECT MASK 1 100.524 16.773 101.202 16.813 ;
      RECT MASK 1 101.354 16.773 102.032 16.813 ;
      RECT MASK 1 102.184 16.773 102.862 16.813 ;
      RECT MASK 1 103.014 16.773 103.692 16.813 ;
      RECT MASK 1 103.844 16.773 104.522 16.813 ;
      RECT MASK 1 104.674 16.773 105.352 16.813 ;
      RECT MASK 1 105.504 16.773 106.182 16.813 ;
      RECT MASK 1 106.334 16.773 107.012 16.813 ;
      RECT MASK 1 107.164 16.773 107.842 16.813 ;
      RECT MASK 1 107.994 16.773 108.672 16.813 ;
      RECT MASK 1 108.824 16.773 109.502 16.813 ;
      RECT MASK 1 109.654 16.773 110.332 16.813 ;
      RECT MASK 1 110.484 16.773 111.162 16.813 ;
      RECT MASK 1 4.327 16.8625 4.507 16.9025 ;
      RECT MASK 1 111.563 16.8625 111.743 16.9025 ;
      RECT MASK 1 5.036 16.957 5.586 16.997 ;
      RECT MASK 1 5.738 16.957 6.288 16.997 ;
      RECT MASK 1 6.696 16.957 7.246 16.997 ;
      RECT MASK 1 7.398 16.957 7.948 16.997 ;
      RECT MASK 1 8.356 16.957 8.906 16.997 ;
      RECT MASK 1 9.058 16.957 9.608 16.997 ;
      RECT MASK 1 10.016 16.957 10.566 16.997 ;
      RECT MASK 1 10.718 16.957 11.268 16.997 ;
      RECT MASK 1 11.676 16.957 12.226 16.997 ;
      RECT MASK 1 12.378 16.957 12.928 16.997 ;
      RECT MASK 1 13.336 16.957 13.886 16.997 ;
      RECT MASK 1 14.038 16.957 14.588 16.997 ;
      RECT MASK 1 14.996 16.957 15.546 16.997 ;
      RECT MASK 1 15.698 16.957 16.248 16.997 ;
      RECT MASK 1 16.656 16.957 17.206 16.997 ;
      RECT MASK 1 17.358 16.957 17.908 16.997 ;
      RECT MASK 1 18.316 16.957 18.866 16.997 ;
      RECT MASK 1 19.018 16.957 19.568 16.997 ;
      RECT MASK 1 19.976 16.957 20.526 16.997 ;
      RECT MASK 1 20.678 16.957 21.228 16.997 ;
      RECT MASK 1 21.636 16.957 22.186 16.997 ;
      RECT MASK 1 22.338 16.957 22.888 16.997 ;
      RECT MASK 1 23.296 16.957 23.846 16.997 ;
      RECT MASK 1 23.998 16.957 24.548 16.997 ;
      RECT MASK 1 24.956 16.957 25.506 16.997 ;
      RECT MASK 1 25.658 16.957 26.208 16.997 ;
      RECT MASK 1 26.616 16.957 27.166 16.997 ;
      RECT MASK 1 27.318 16.957 27.868 16.997 ;
      RECT MASK 1 28.276 16.957 28.826 16.997 ;
      RECT MASK 1 28.978 16.957 29.528 16.997 ;
      RECT MASK 1 29.936 16.957 30.486 16.997 ;
      RECT MASK 1 30.638 16.957 31.188 16.997 ;
      RECT MASK 1 31.596 16.957 32.146 16.997 ;
      RECT MASK 1 32.298 16.957 32.848 16.997 ;
      RECT MASK 1 33.256 16.957 33.806 16.997 ;
      RECT MASK 1 33.958 16.957 34.508 16.997 ;
      RECT MASK 1 34.916 16.957 35.466 16.997 ;
      RECT MASK 1 35.618 16.957 36.168 16.997 ;
      RECT MASK 1 36.576 16.957 37.126 16.997 ;
      RECT MASK 1 37.278 16.957 37.828 16.997 ;
      RECT MASK 1 38.236 16.957 38.786 16.997 ;
      RECT MASK 1 38.938 16.957 39.488 16.997 ;
      RECT MASK 1 39.896 16.957 40.446 16.997 ;
      RECT MASK 1 40.598 16.957 41.148 16.997 ;
      RECT MASK 1 41.556 16.957 42.106 16.997 ;
      RECT MASK 1 42.258 16.957 42.808 16.997 ;
      RECT MASK 1 43.216 16.957 43.766 16.997 ;
      RECT MASK 1 43.918 16.957 44.468 16.997 ;
      RECT MASK 1 44.876 16.957 45.426 16.997 ;
      RECT MASK 1 45.578 16.957 46.128 16.997 ;
      RECT MASK 1 46.536 16.957 47.086 16.997 ;
      RECT MASK 1 47.238 16.957 47.788 16.997 ;
      RECT MASK 1 48.196 16.957 48.746 16.997 ;
      RECT MASK 1 48.898 16.957 49.448 16.997 ;
      RECT MASK 1 49.856 16.957 50.406 16.997 ;
      RECT MASK 1 50.558 16.957 51.108 16.997 ;
      RECT MASK 1 51.516 16.957 52.066 16.997 ;
      RECT MASK 1 52.218 16.957 52.768 16.997 ;
      RECT MASK 1 53.176 16.957 53.726 16.997 ;
      RECT MASK 1 53.878 16.957 54.428 16.997 ;
      RECT MASK 1 54.836 16.957 55.386 16.997 ;
      RECT MASK 1 55.538 16.957 56.088 16.997 ;
      RECT MASK 1 56.662 16.957 57.212 16.997 ;
      RECT MASK 1 57.364 16.957 57.914 16.997 ;
      RECT MASK 1 58.322 16.957 58.872 16.997 ;
      RECT MASK 1 59.024 16.957 59.574 16.997 ;
      RECT MASK 1 59.982 16.957 60.532 16.997 ;
      RECT MASK 1 60.684 16.957 61.234 16.997 ;
      RECT MASK 1 61.642 16.957 62.192 16.997 ;
      RECT MASK 1 62.344 16.957 62.894 16.997 ;
      RECT MASK 1 63.302 16.957 63.852 16.997 ;
      RECT MASK 1 64.004 16.957 64.554 16.997 ;
      RECT MASK 1 64.962 16.957 65.512 16.997 ;
      RECT MASK 1 65.664 16.957 66.214 16.997 ;
      RECT MASK 1 66.622 16.957 67.172 16.997 ;
      RECT MASK 1 67.324 16.957 67.874 16.997 ;
      RECT MASK 1 68.282 16.957 68.832 16.997 ;
      RECT MASK 1 68.984 16.957 69.534 16.997 ;
      RECT MASK 1 69.942 16.957 70.492 16.997 ;
      RECT MASK 1 70.644 16.957 71.194 16.997 ;
      RECT MASK 1 71.602 16.957 72.152 16.997 ;
      RECT MASK 1 72.304 16.957 72.854 16.997 ;
      RECT MASK 1 73.262 16.957 73.812 16.997 ;
      RECT MASK 1 73.964 16.957 74.514 16.997 ;
      RECT MASK 1 74.922 16.957 75.472 16.997 ;
      RECT MASK 1 75.624 16.957 76.174 16.997 ;
      RECT MASK 1 76.582 16.957 77.132 16.997 ;
      RECT MASK 1 77.284 16.957 77.834 16.997 ;
      RECT MASK 1 78.242 16.957 78.792 16.997 ;
      RECT MASK 1 78.944 16.957 79.494 16.997 ;
      RECT MASK 1 79.902 16.957 80.452 16.997 ;
      RECT MASK 1 80.604 16.957 81.154 16.997 ;
      RECT MASK 1 81.562 16.957 82.112 16.997 ;
      RECT MASK 1 82.264 16.957 82.814 16.997 ;
      RECT MASK 1 83.222 16.957 83.772 16.997 ;
      RECT MASK 1 83.924 16.957 84.474 16.997 ;
      RECT MASK 1 84.882 16.957 85.432 16.997 ;
      RECT MASK 1 85.584 16.957 86.134 16.997 ;
      RECT MASK 1 86.542 16.957 87.092 16.997 ;
      RECT MASK 1 87.244 16.957 87.794 16.997 ;
      RECT MASK 1 88.202 16.957 88.752 16.997 ;
      RECT MASK 1 88.904 16.957 89.454 16.997 ;
      RECT MASK 1 89.862 16.957 90.412 16.997 ;
      RECT MASK 1 90.564 16.957 91.114 16.997 ;
      RECT MASK 1 91.522 16.957 92.072 16.997 ;
      RECT MASK 1 92.224 16.957 92.774 16.997 ;
      RECT MASK 1 93.182 16.957 93.732 16.997 ;
      RECT MASK 1 93.884 16.957 94.434 16.997 ;
      RECT MASK 1 94.842 16.957 95.392 16.997 ;
      RECT MASK 1 95.544 16.957 96.094 16.997 ;
      RECT MASK 1 96.502 16.957 97.052 16.997 ;
      RECT MASK 1 97.204 16.957 97.754 16.997 ;
      RECT MASK 1 98.162 16.957 98.712 16.997 ;
      RECT MASK 1 98.864 16.957 99.414 16.997 ;
      RECT MASK 1 99.822 16.957 100.372 16.997 ;
      RECT MASK 1 100.524 16.957 101.074 16.997 ;
      RECT MASK 1 101.482 16.957 102.032 16.997 ;
      RECT MASK 1 102.184 16.957 102.734 16.997 ;
      RECT MASK 1 103.142 16.957 103.692 16.997 ;
      RECT MASK 1 103.844 16.957 104.394 16.997 ;
      RECT MASK 1 104.802 16.957 105.352 16.997 ;
      RECT MASK 1 105.504 16.957 106.054 16.997 ;
      RECT MASK 1 106.462 16.957 107.012 16.997 ;
      RECT MASK 1 107.164 16.957 107.714 16.997 ;
      RECT MASK 1 108.122 16.957 108.672 16.997 ;
      RECT MASK 1 108.824 16.957 109.374 16.997 ;
      RECT MASK 1 109.782 16.957 110.332 16.997 ;
      RECT MASK 1 110.484 16.957 111.034 16.997 ;
      RECT MASK 1 4.251 17.124 111.819 17.164 ;
      RECT MASK 1 116.154 17.28 116.214 18.33 ;
      RECT MASK 1 116.428 17.28 116.488 18.33 ;
      RECT MASK 1 116.702 17.28 116.762 18.33 ;
      RECT MASK 1 116.976 17.28 117.036 18.33 ;
      RECT MASK 1 117.25 17.28 117.31 18.33 ;
      RECT MASK 1 117.524 17.28 117.584 18.33 ;
      RECT MASK 1 117.798 17.28 117.858 18.33 ;
      RECT MASK 1 118.072 17.28 118.132 18.33 ;
      RECT MASK 1 118.346 17.28 118.406 18.33 ;
      RECT MASK 1 118.62 17.28 118.68 18.33 ;
      RECT MASK 1 118.894 17.28 118.954 18.33 ;
      RECT MASK 1 119.168 17.28 119.228 18.33 ;
      RECT MASK 1 119.442 17.28 119.502 18.33 ;
      RECT MASK 1 119.716 17.28 119.776 18.33 ;
      RECT MASK 1 119.99 17.28 120.05 18.33 ;
      RECT MASK 1 120.264 17.28 120.324 18.33 ;
      RECT MASK 1 120.538 17.28 120.598 18.33 ;
      RECT MASK 1 120.812 17.28 120.872 18.33 ;
      RECT MASK 1 121.086 17.28 121.146 18.33 ;
      RECT MASK 1 121.36 17.28 121.42 18.33 ;
      RECT MASK 1 121.634 17.28 121.694 18.33 ;
      RECT MASK 1 121.908 17.28 121.968 18.33 ;
      RECT MASK 1 122.182 17.28 122.242 18.33 ;
      RECT MASK 1 122.456 17.28 122.516 18.33 ;
      RECT MASK 1 122.73 17.28 122.79 18.33 ;
      RECT MASK 1 123.004 17.28 123.064 18.33 ;
      RECT MASK 1 123.278 17.28 123.338 18.33 ;
      RECT MASK 1 123.552 17.28 123.612 18.33 ;
      RECT MASK 1 123.826 17.28 123.886 18.33 ;
      RECT MASK 1 124.1 17.28 124.16 18.33 ;
      RECT MASK 1 124.374 17.28 124.434 18.33 ;
      RECT MASK 1 124.648 17.28 124.708 18.33 ;
      RECT MASK 1 124.922 17.28 124.982 18.33 ;
      RECT MASK 1 125.196 17.28 125.256 18.33 ;
      RECT MASK 1 125.47 17.28 125.53 18.33 ;
      RECT MASK 1 125.744 17.28 125.804 18.33 ;
      RECT MASK 1 126.018 17.28 126.078 18.33 ;
      RECT MASK 1 126.292 17.28 126.352 18.33 ;
      RECT MASK 1 126.566 17.28 126.626 18.33 ;
      RECT MASK 1 126.84 17.28 126.9 18.33 ;
      RECT MASK 1 127.114 17.28 127.174 18.33 ;
      RECT MASK 1 127.388 17.28 127.448 18.33 ;
      RECT MASK 1 127.662 17.28 127.722 18.33 ;
      RECT MASK 1 127.936 17.28 127.996 18.33 ;
      RECT MASK 1 128.21 17.28 128.27 18.33 ;
      RECT MASK 1 4.251 17.299 111.819 17.339 ;
      RECT MASK 1 4.362 17.62 111.708 17.66 ;
      RECT MASK 1 5.062 18.055 109.834 18.095 ;
      RECT MASK 1 5.062 18.391 109.819 18.431 ;
      RECT MASK 1 5.062 18.575 109.898 18.615 ;
      RECT MASK 1 5.816 18.759 5.999 18.799 ;
      RECT MASK 1 6.221 18.759 6.404 18.799 ;
      RECT MASK 1 6.978 18.759 7.161 18.799 ;
      RECT MASK 1 7.383 18.759 7.566 18.799 ;
      RECT MASK 1 8.14 18.759 8.323 18.799 ;
      RECT MASK 1 8.545 18.759 8.728 18.799 ;
      RECT MASK 1 9.302 18.759 9.485 18.799 ;
      RECT MASK 1 9.707 18.759 9.89 18.799 ;
      RECT MASK 1 12.434 18.759 12.617 18.799 ;
      RECT MASK 1 12.839 18.759 13.022 18.799 ;
      RECT MASK 1 13.596 18.759 13.779 18.799 ;
      RECT MASK 1 14.001 18.759 14.184 18.799 ;
      RECT MASK 1 14.758 18.759 14.941 18.799 ;
      RECT MASK 1 15.163 18.759 15.346 18.799 ;
      RECT MASK 1 15.92 18.759 16.103 18.799 ;
      RECT MASK 1 16.325 18.759 16.508 18.799 ;
      RECT MASK 1 19.052 18.759 19.235 18.799 ;
      RECT MASK 1 19.457 18.759 19.64 18.799 ;
      RECT MASK 1 20.214 18.759 20.397 18.799 ;
      RECT MASK 1 20.619 18.759 20.802 18.799 ;
      RECT MASK 1 21.376 18.759 21.559 18.799 ;
      RECT MASK 1 21.781 18.759 21.964 18.799 ;
      RECT MASK 1 22.538 18.759 22.721 18.799 ;
      RECT MASK 1 22.943 18.759 23.126 18.799 ;
      RECT MASK 1 25.67 18.759 25.853 18.799 ;
      RECT MASK 1 26.075 18.759 26.258 18.799 ;
      RECT MASK 1 26.832 18.759 27.015 18.799 ;
      RECT MASK 1 27.237 18.759 27.42 18.799 ;
      RECT MASK 1 27.994 18.759 28.177 18.799 ;
      RECT MASK 1 28.399 18.759 28.582 18.799 ;
      RECT MASK 1 29.156 18.759 29.339 18.799 ;
      RECT MASK 1 29.561 18.759 29.744 18.799 ;
      RECT MASK 1 32.288 18.759 32.471 18.799 ;
      RECT MASK 1 32.693 18.759 32.876 18.799 ;
      RECT MASK 1 33.45 18.759 33.633 18.799 ;
      RECT MASK 1 33.855 18.759 34.038 18.799 ;
      RECT MASK 1 34.612 18.759 34.795 18.799 ;
      RECT MASK 1 35.017 18.759 35.2 18.799 ;
      RECT MASK 1 35.774 18.759 35.957 18.799 ;
      RECT MASK 1 36.179 18.759 36.362 18.799 ;
      RECT MASK 1 38.906 18.759 39.089 18.799 ;
      RECT MASK 1 39.311 18.759 39.494 18.799 ;
      RECT MASK 1 40.068 18.759 40.251 18.799 ;
      RECT MASK 1 40.473 18.759 40.656 18.799 ;
      RECT MASK 1 41.23 18.759 41.413 18.799 ;
      RECT MASK 1 41.635 18.759 41.818 18.799 ;
      RECT MASK 1 42.392 18.759 42.575 18.799 ;
      RECT MASK 1 42.797 18.759 42.98 18.799 ;
      RECT MASK 1 45.524 18.759 45.707 18.799 ;
      RECT MASK 1 45.929 18.759 46.112 18.799 ;
      RECT MASK 1 46.686 18.759 46.869 18.799 ;
      RECT MASK 1 47.091 18.759 47.274 18.799 ;
      RECT MASK 1 47.848 18.759 48.031 18.799 ;
      RECT MASK 1 48.253 18.759 48.436 18.799 ;
      RECT MASK 1 49.01 18.759 49.193 18.799 ;
      RECT MASK 1 49.415 18.759 49.598 18.799 ;
      RECT MASK 1 52.142 18.759 52.325 18.799 ;
      RECT MASK 1 52.547 18.759 52.73 18.799 ;
      RECT MASK 1 53.304 18.759 53.487 18.799 ;
      RECT MASK 1 53.709 18.759 53.892 18.799 ;
      RECT MASK 1 54.466 18.759 54.649 18.799 ;
      RECT MASK 1 54.871 18.759 55.054 18.799 ;
      RECT MASK 1 55.628 18.759 55.811 18.799 ;
      RECT MASK 1 56.033 18.759 56.216 18.799 ;
      RECT MASK 1 58.76 18.759 58.943 18.799 ;
      RECT MASK 1 59.165 18.759 59.348 18.799 ;
      RECT MASK 1 59.922 18.759 60.105 18.799 ;
      RECT MASK 1 60.327 18.759 60.51 18.799 ;
      RECT MASK 1 61.084 18.759 61.267 18.799 ;
      RECT MASK 1 61.489 18.759 61.672 18.799 ;
      RECT MASK 1 62.246 18.759 62.429 18.799 ;
      RECT MASK 1 62.651 18.759 62.834 18.799 ;
      RECT MASK 1 65.378 18.759 65.561 18.799 ;
      RECT MASK 1 65.783 18.759 65.966 18.799 ;
      RECT MASK 1 66.54 18.759 66.723 18.799 ;
      RECT MASK 1 66.945 18.759 67.128 18.799 ;
      RECT MASK 1 67.702 18.759 67.885 18.799 ;
      RECT MASK 1 68.107 18.759 68.29 18.799 ;
      RECT MASK 1 68.864 18.759 69.047 18.799 ;
      RECT MASK 1 69.269 18.759 69.452 18.799 ;
      RECT MASK 1 71.996 18.759 72.179 18.799 ;
      RECT MASK 1 72.401 18.759 72.584 18.799 ;
      RECT MASK 1 73.158 18.759 73.341 18.799 ;
      RECT MASK 1 73.563 18.759 73.746 18.799 ;
      RECT MASK 1 74.32 18.759 74.503 18.799 ;
      RECT MASK 1 74.725 18.759 74.908 18.799 ;
      RECT MASK 1 75.482 18.759 75.665 18.799 ;
      RECT MASK 1 75.887 18.759 76.07 18.799 ;
      RECT MASK 1 78.614 18.759 78.797 18.799 ;
      RECT MASK 1 79.019 18.759 79.202 18.799 ;
      RECT MASK 1 79.776 18.759 79.959 18.799 ;
      RECT MASK 1 80.181 18.759 80.364 18.799 ;
      RECT MASK 1 80.938 18.759 81.121 18.799 ;
      RECT MASK 1 81.343 18.759 81.526 18.799 ;
      RECT MASK 1 82.1 18.759 82.283 18.799 ;
      RECT MASK 1 82.505 18.759 82.688 18.799 ;
      RECT MASK 1 85.232 18.759 85.415 18.799 ;
      RECT MASK 1 85.637 18.759 85.82 18.799 ;
      RECT MASK 1 86.394 18.759 86.577 18.799 ;
      RECT MASK 1 86.799 18.759 86.982 18.799 ;
      RECT MASK 1 87.556 18.759 87.739 18.799 ;
      RECT MASK 1 87.961 18.759 88.144 18.799 ;
      RECT MASK 1 88.718 18.759 88.901 18.799 ;
      RECT MASK 1 89.123 18.759 89.306 18.799 ;
      RECT MASK 1 91.85 18.759 92.033 18.799 ;
      RECT MASK 1 92.255 18.759 92.438 18.799 ;
      RECT MASK 1 93.012 18.759 93.195 18.799 ;
      RECT MASK 1 93.417 18.759 93.6 18.799 ;
      RECT MASK 1 94.174 18.759 94.357 18.799 ;
      RECT MASK 1 94.579 18.759 94.762 18.799 ;
      RECT MASK 1 95.336 18.759 95.519 18.799 ;
      RECT MASK 1 95.741 18.759 95.924 18.799 ;
      RECT MASK 1 98.468 18.759 98.651 18.799 ;
      RECT MASK 1 98.873 18.759 99.056 18.799 ;
      RECT MASK 1 99.63 18.759 99.813 18.799 ;
      RECT MASK 1 100.035 18.759 100.218 18.799 ;
      RECT MASK 1 100.792 18.759 100.975 18.799 ;
      RECT MASK 1 101.197 18.759 101.38 18.799 ;
      RECT MASK 1 101.954 18.759 102.137 18.799 ;
      RECT MASK 1 102.359 18.759 102.542 18.799 ;
      RECT MASK 1 105.086 18.759 105.269 18.799 ;
      RECT MASK 1 105.491 18.759 105.674 18.799 ;
      RECT MASK 1 106.248 18.759 106.431 18.799 ;
      RECT MASK 1 106.653 18.759 106.836 18.799 ;
      RECT MASK 1 107.41 18.759 107.593 18.799 ;
      RECT MASK 1 107.815 18.759 107.998 18.799 ;
      RECT MASK 1 108.572 18.759 108.755 18.799 ;
      RECT MASK 1 108.977 18.759 109.16 18.799 ;
      RECT MASK 1 5.816 18.927 5.999 18.967 ;
      RECT MASK 1 6.221 18.927 6.404 18.967 ;
      RECT MASK 1 6.978 18.927 7.161 18.967 ;
      RECT MASK 1 7.383 18.927 7.566 18.967 ;
      RECT MASK 1 8.14 18.927 8.323 18.967 ;
      RECT MASK 1 8.545 18.927 8.728 18.967 ;
      RECT MASK 1 9.302 18.927 9.485 18.967 ;
      RECT MASK 1 9.707 18.927 9.89 18.967 ;
      RECT MASK 1 12.434 18.927 12.617 18.967 ;
      RECT MASK 1 12.839 18.927 13.022 18.967 ;
      RECT MASK 1 13.596 18.927 13.779 18.967 ;
      RECT MASK 1 14.001 18.927 14.184 18.967 ;
      RECT MASK 1 14.758 18.927 14.941 18.967 ;
      RECT MASK 1 15.163 18.927 15.346 18.967 ;
      RECT MASK 1 15.92 18.927 16.103 18.967 ;
      RECT MASK 1 16.325 18.927 16.508 18.967 ;
      RECT MASK 1 19.052 18.927 19.235 18.967 ;
      RECT MASK 1 19.457 18.927 19.64 18.967 ;
      RECT MASK 1 20.214 18.927 20.397 18.967 ;
      RECT MASK 1 20.619 18.927 20.802 18.967 ;
      RECT MASK 1 21.376 18.927 21.559 18.967 ;
      RECT MASK 1 21.781 18.927 21.964 18.967 ;
      RECT MASK 1 22.538 18.927 22.721 18.967 ;
      RECT MASK 1 22.943 18.927 23.126 18.967 ;
      RECT MASK 1 25.67 18.927 25.853 18.967 ;
      RECT MASK 1 26.075 18.927 26.258 18.967 ;
      RECT MASK 1 26.832 18.927 27.015 18.967 ;
      RECT MASK 1 27.237 18.927 27.42 18.967 ;
      RECT MASK 1 27.994 18.927 28.177 18.967 ;
      RECT MASK 1 28.399 18.927 28.582 18.967 ;
      RECT MASK 1 29.156 18.927 29.339 18.967 ;
      RECT MASK 1 29.561 18.927 29.744 18.967 ;
      RECT MASK 1 32.288 18.927 32.471 18.967 ;
      RECT MASK 1 32.693 18.927 32.876 18.967 ;
      RECT MASK 1 33.45 18.927 33.633 18.967 ;
      RECT MASK 1 33.855 18.927 34.038 18.967 ;
      RECT MASK 1 34.612 18.927 34.795 18.967 ;
      RECT MASK 1 35.017 18.927 35.2 18.967 ;
      RECT MASK 1 35.774 18.927 35.957 18.967 ;
      RECT MASK 1 36.179 18.927 36.362 18.967 ;
      RECT MASK 1 38.906 18.927 39.089 18.967 ;
      RECT MASK 1 39.311 18.927 39.494 18.967 ;
      RECT MASK 1 40.068 18.927 40.251 18.967 ;
      RECT MASK 1 40.473 18.927 40.656 18.967 ;
      RECT MASK 1 41.23 18.927 41.413 18.967 ;
      RECT MASK 1 41.635 18.927 41.818 18.967 ;
      RECT MASK 1 42.392 18.927 42.575 18.967 ;
      RECT MASK 1 42.797 18.927 42.98 18.967 ;
      RECT MASK 1 45.524 18.927 45.707 18.967 ;
      RECT MASK 1 45.929 18.927 46.112 18.967 ;
      RECT MASK 1 46.686 18.927 46.869 18.967 ;
      RECT MASK 1 47.091 18.927 47.274 18.967 ;
      RECT MASK 1 47.848 18.927 48.031 18.967 ;
      RECT MASK 1 48.253 18.927 48.436 18.967 ;
      RECT MASK 1 49.01 18.927 49.193 18.967 ;
      RECT MASK 1 49.415 18.927 49.598 18.967 ;
      RECT MASK 1 52.142 18.927 52.325 18.967 ;
      RECT MASK 1 52.547 18.927 52.73 18.967 ;
      RECT MASK 1 53.304 18.927 53.487 18.967 ;
      RECT MASK 1 53.709 18.927 53.892 18.967 ;
      RECT MASK 1 54.466 18.927 54.649 18.967 ;
      RECT MASK 1 54.871 18.927 55.054 18.967 ;
      RECT MASK 1 55.628 18.927 55.811 18.967 ;
      RECT MASK 1 56.033 18.927 56.216 18.967 ;
      RECT MASK 1 58.76 18.927 58.943 18.967 ;
      RECT MASK 1 59.165 18.927 59.348 18.967 ;
      RECT MASK 1 59.922 18.927 60.105 18.967 ;
      RECT MASK 1 60.327 18.927 60.51 18.967 ;
      RECT MASK 1 61.084 18.927 61.267 18.967 ;
      RECT MASK 1 61.489 18.927 61.672 18.967 ;
      RECT MASK 1 62.246 18.927 62.429 18.967 ;
      RECT MASK 1 62.651 18.927 62.834 18.967 ;
      RECT MASK 1 65.378 18.927 65.561 18.967 ;
      RECT MASK 1 65.783 18.927 65.966 18.967 ;
      RECT MASK 1 66.54 18.927 66.723 18.967 ;
      RECT MASK 1 66.945 18.927 67.128 18.967 ;
      RECT MASK 1 67.702 18.927 67.885 18.967 ;
      RECT MASK 1 68.107 18.927 68.29 18.967 ;
      RECT MASK 1 68.864 18.927 69.047 18.967 ;
      RECT MASK 1 69.269 18.927 69.452 18.967 ;
      RECT MASK 1 71.996 18.927 72.179 18.967 ;
      RECT MASK 1 72.401 18.927 72.584 18.967 ;
      RECT MASK 1 73.158 18.927 73.341 18.967 ;
      RECT MASK 1 73.563 18.927 73.746 18.967 ;
      RECT MASK 1 74.32 18.927 74.503 18.967 ;
      RECT MASK 1 74.725 18.927 74.908 18.967 ;
      RECT MASK 1 75.482 18.927 75.665 18.967 ;
      RECT MASK 1 75.887 18.927 76.07 18.967 ;
      RECT MASK 1 78.614 18.927 78.797 18.967 ;
      RECT MASK 1 79.019 18.927 79.202 18.967 ;
      RECT MASK 1 79.776 18.927 79.959 18.967 ;
      RECT MASK 1 80.181 18.927 80.364 18.967 ;
      RECT MASK 1 80.938 18.927 81.121 18.967 ;
      RECT MASK 1 81.343 18.927 81.526 18.967 ;
      RECT MASK 1 82.1 18.927 82.283 18.967 ;
      RECT MASK 1 82.505 18.927 82.688 18.967 ;
      RECT MASK 1 85.232 18.927 85.415 18.967 ;
      RECT MASK 1 85.637 18.927 85.82 18.967 ;
      RECT MASK 1 86.394 18.927 86.577 18.967 ;
      RECT MASK 1 86.799 18.927 86.982 18.967 ;
      RECT MASK 1 87.556 18.927 87.739 18.967 ;
      RECT MASK 1 87.961 18.927 88.144 18.967 ;
      RECT MASK 1 88.718 18.927 88.901 18.967 ;
      RECT MASK 1 89.123 18.927 89.306 18.967 ;
      RECT MASK 1 91.85 18.927 92.033 18.967 ;
      RECT MASK 1 92.255 18.927 92.438 18.967 ;
      RECT MASK 1 93.012 18.927 93.195 18.967 ;
      RECT MASK 1 93.417 18.927 93.6 18.967 ;
      RECT MASK 1 94.174 18.927 94.357 18.967 ;
      RECT MASK 1 94.579 18.927 94.762 18.967 ;
      RECT MASK 1 95.336 18.927 95.519 18.967 ;
      RECT MASK 1 95.741 18.927 95.924 18.967 ;
      RECT MASK 1 98.468 18.927 98.651 18.967 ;
      RECT MASK 1 98.873 18.927 99.056 18.967 ;
      RECT MASK 1 99.63 18.927 99.813 18.967 ;
      RECT MASK 1 100.035 18.927 100.218 18.967 ;
      RECT MASK 1 100.792 18.927 100.975 18.967 ;
      RECT MASK 1 101.197 18.927 101.38 18.967 ;
      RECT MASK 1 101.954 18.927 102.137 18.967 ;
      RECT MASK 1 102.359 18.927 102.542 18.967 ;
      RECT MASK 1 105.086 18.927 105.269 18.967 ;
      RECT MASK 1 105.491 18.927 105.674 18.967 ;
      RECT MASK 1 106.248 18.927 106.431 18.967 ;
      RECT MASK 1 106.653 18.927 106.836 18.967 ;
      RECT MASK 1 107.41 18.927 107.593 18.967 ;
      RECT MASK 1 107.815 18.927 107.998 18.967 ;
      RECT MASK 1 108.572 18.927 108.755 18.967 ;
      RECT MASK 1 108.977 18.927 109.16 18.967 ;
      RECT MASK 1 5.107 18.981 5.287 19.021 ;
      RECT MASK 1 10.419 18.981 10.599 19.021 ;
      RECT MASK 1 11.725 18.981 11.905 19.021 ;
      RECT MASK 1 17.037 18.981 17.217 19.021 ;
      RECT MASK 1 18.343 18.981 18.523 19.021 ;
      RECT MASK 1 23.655 18.981 23.835 19.021 ;
      RECT MASK 1 24.961 18.981 25.141 19.021 ;
      RECT MASK 1 30.273 18.981 30.453 19.021 ;
      RECT MASK 1 31.579 18.981 31.759 19.021 ;
      RECT MASK 1 36.891 18.981 37.071 19.021 ;
      RECT MASK 1 38.197 18.981 38.377 19.021 ;
      RECT MASK 1 43.509 18.981 43.689 19.021 ;
      RECT MASK 1 44.815 18.981 44.995 19.021 ;
      RECT MASK 1 50.127 18.981 50.307 19.021 ;
      RECT MASK 1 51.433 18.981 51.613 19.021 ;
      RECT MASK 1 56.745 18.981 56.925 19.021 ;
      RECT MASK 1 58.051 18.981 58.231 19.021 ;
      RECT MASK 1 63.363 18.981 63.543 19.021 ;
      RECT MASK 1 64.669 18.981 64.849 19.021 ;
      RECT MASK 1 69.981 18.981 70.161 19.021 ;
      RECT MASK 1 71.287 18.981 71.467 19.021 ;
      RECT MASK 1 76.599 18.981 76.779 19.021 ;
      RECT MASK 1 77.905 18.981 78.085 19.021 ;
      RECT MASK 1 83.217 18.981 83.397 19.021 ;
      RECT MASK 1 84.523 18.981 84.703 19.021 ;
      RECT MASK 1 89.835 18.981 90.015 19.021 ;
      RECT MASK 1 91.141 18.981 91.321 19.021 ;
      RECT MASK 1 96.453 18.981 96.633 19.021 ;
      RECT MASK 1 97.759 18.981 97.939 19.021 ;
      RECT MASK 1 103.071 18.981 103.251 19.021 ;
      RECT MASK 1 104.377 18.981 104.557 19.021 ;
      RECT MASK 1 109.689 18.981 109.869 19.021 ;
      RECT MASK 1 116.154 18.99 116.214 20.04 ;
      RECT MASK 1 116.428 18.99 116.488 20.04 ;
      RECT MASK 1 116.702 18.99 116.762 20.04 ;
      RECT MASK 1 116.976 18.99 117.036 20.04 ;
      RECT MASK 1 117.25 18.99 117.31 20.04 ;
      RECT MASK 1 117.524 18.99 117.584 20.04 ;
      RECT MASK 1 117.798 18.99 117.858 20.04 ;
      RECT MASK 1 118.072 18.99 118.132 20.04 ;
      RECT MASK 1 118.346 18.99 118.406 20.04 ;
      RECT MASK 1 118.62 18.99 118.68 20.04 ;
      RECT MASK 1 118.894 18.99 118.954 20.04 ;
      RECT MASK 1 119.168 18.99 119.228 20.04 ;
      RECT MASK 1 119.442 18.99 119.502 20.04 ;
      RECT MASK 1 119.716 18.99 119.776 20.04 ;
      RECT MASK 1 119.99 18.99 120.05 20.04 ;
      RECT MASK 1 120.264 18.99 120.324 20.04 ;
      RECT MASK 1 120.538 18.99 120.598 20.04 ;
      RECT MASK 1 120.812 18.99 120.872 20.04 ;
      RECT MASK 1 121.086 18.99 121.146 20.04 ;
      RECT MASK 1 121.36 18.99 121.42 20.04 ;
      RECT MASK 1 121.634 18.99 121.694 20.04 ;
      RECT MASK 1 121.908 18.99 121.968 20.04 ;
      RECT MASK 1 122.182 18.99 122.242 20.04 ;
      RECT MASK 1 122.456 18.99 122.516 20.04 ;
      RECT MASK 1 122.73 18.99 122.79 20.04 ;
      RECT MASK 1 123.004 18.99 123.064 20.04 ;
      RECT MASK 1 123.278 18.99 123.338 20.04 ;
      RECT MASK 1 123.552 18.99 123.612 20.04 ;
      RECT MASK 1 123.826 18.99 123.886 20.04 ;
      RECT MASK 1 124.1 18.99 124.16 20.04 ;
      RECT MASK 1 124.374 18.99 124.434 20.04 ;
      RECT MASK 1 124.648 18.99 124.708 20.04 ;
      RECT MASK 1 124.922 18.99 124.982 20.04 ;
      RECT MASK 1 125.196 18.99 125.256 20.04 ;
      RECT MASK 1 125.47 18.99 125.53 20.04 ;
      RECT MASK 1 125.744 18.99 125.804 20.04 ;
      RECT MASK 1 126.018 18.99 126.078 20.04 ;
      RECT MASK 1 126.292 18.99 126.352 20.04 ;
      RECT MASK 1 126.566 18.99 126.626 20.04 ;
      RECT MASK 1 126.84 18.99 126.9 20.04 ;
      RECT MASK 1 127.114 18.99 127.174 20.04 ;
      RECT MASK 1 127.388 18.99 127.448 20.04 ;
      RECT MASK 1 127.662 18.99 127.722 20.04 ;
      RECT MASK 1 127.936 18.99 127.996 20.04 ;
      RECT MASK 1 128.21 18.99 128.27 20.04 ;
      RECT MASK 1 5.107 19.149 5.287 19.189 ;
      RECT MASK 1 5.688 19.149 5.868 19.189 ;
      RECT MASK 1 6.352 19.149 6.532 19.189 ;
      RECT MASK 1 6.85 19.149 7.03 19.189 ;
      RECT MASK 1 7.514 19.149 7.694 19.189 ;
      RECT MASK 1 8.012 19.149 8.192 19.189 ;
      RECT MASK 1 8.676 19.149 8.856 19.189 ;
      RECT MASK 1 9.174 19.149 9.354 19.189 ;
      RECT MASK 1 9.838 19.149 10.018 19.189 ;
      RECT MASK 1 10.419 19.149 10.599 19.189 ;
      RECT MASK 1 11.725 19.149 11.905 19.189 ;
      RECT MASK 1 12.306 19.149 12.486 19.189 ;
      RECT MASK 1 12.97 19.149 13.15 19.189 ;
      RECT MASK 1 13.468 19.149 13.648 19.189 ;
      RECT MASK 1 14.132 19.149 14.312 19.189 ;
      RECT MASK 1 14.63 19.149 14.81 19.189 ;
      RECT MASK 1 15.294 19.149 15.474 19.189 ;
      RECT MASK 1 15.792 19.149 15.972 19.189 ;
      RECT MASK 1 16.456 19.149 16.636 19.189 ;
      RECT MASK 1 17.037 19.149 17.217 19.189 ;
      RECT MASK 1 18.343 19.149 18.523 19.189 ;
      RECT MASK 1 18.924 19.149 19.104 19.189 ;
      RECT MASK 1 19.588 19.149 19.768 19.189 ;
      RECT MASK 1 20.086 19.149 20.266 19.189 ;
      RECT MASK 1 20.75 19.149 20.93 19.189 ;
      RECT MASK 1 21.248 19.149 21.428 19.189 ;
      RECT MASK 1 21.912 19.149 22.092 19.189 ;
      RECT MASK 1 22.41 19.149 22.59 19.189 ;
      RECT MASK 1 23.074 19.149 23.254 19.189 ;
      RECT MASK 1 23.655 19.149 23.835 19.189 ;
      RECT MASK 1 24.961 19.149 25.141 19.189 ;
      RECT MASK 1 25.542 19.149 25.722 19.189 ;
      RECT MASK 1 26.206 19.149 26.386 19.189 ;
      RECT MASK 1 26.704 19.149 26.884 19.189 ;
      RECT MASK 1 27.368 19.149 27.548 19.189 ;
      RECT MASK 1 27.866 19.149 28.046 19.189 ;
      RECT MASK 1 28.53 19.149 28.71 19.189 ;
      RECT MASK 1 29.028 19.149 29.208 19.189 ;
      RECT MASK 1 29.692 19.149 29.872 19.189 ;
      RECT MASK 1 30.273 19.149 30.453 19.189 ;
      RECT MASK 1 31.579 19.149 31.759 19.189 ;
      RECT MASK 1 32.16 19.149 32.34 19.189 ;
      RECT MASK 1 32.824 19.149 33.004 19.189 ;
      RECT MASK 1 33.322 19.149 33.502 19.189 ;
      RECT MASK 1 33.986 19.149 34.166 19.189 ;
      RECT MASK 1 34.484 19.149 34.664 19.189 ;
      RECT MASK 1 35.148 19.149 35.328 19.189 ;
      RECT MASK 1 35.646 19.149 35.826 19.189 ;
      RECT MASK 1 36.31 19.149 36.49 19.189 ;
      RECT MASK 1 36.891 19.149 37.071 19.189 ;
      RECT MASK 1 38.197 19.149 38.377 19.189 ;
      RECT MASK 1 38.778 19.149 38.958 19.189 ;
      RECT MASK 1 39.442 19.149 39.622 19.189 ;
      RECT MASK 1 39.94 19.149 40.12 19.189 ;
      RECT MASK 1 40.604 19.149 40.784 19.189 ;
      RECT MASK 1 41.102 19.149 41.282 19.189 ;
      RECT MASK 1 41.766 19.149 41.946 19.189 ;
      RECT MASK 1 42.264 19.149 42.444 19.189 ;
      RECT MASK 1 42.928 19.149 43.108 19.189 ;
      RECT MASK 1 43.509 19.149 43.689 19.189 ;
      RECT MASK 1 44.815 19.149 44.995 19.189 ;
      RECT MASK 1 45.396 19.149 45.576 19.189 ;
      RECT MASK 1 46.06 19.149 46.24 19.189 ;
      RECT MASK 1 46.558 19.149 46.738 19.189 ;
      RECT MASK 1 47.222 19.149 47.402 19.189 ;
      RECT MASK 1 47.72 19.149 47.9 19.189 ;
      RECT MASK 1 48.384 19.149 48.564 19.189 ;
      RECT MASK 1 48.882 19.149 49.062 19.189 ;
      RECT MASK 1 49.546 19.149 49.726 19.189 ;
      RECT MASK 1 50.127 19.149 50.307 19.189 ;
      RECT MASK 1 51.433 19.149 51.613 19.189 ;
      RECT MASK 1 52.014 19.149 52.194 19.189 ;
      RECT MASK 1 52.678 19.149 52.858 19.189 ;
      RECT MASK 1 53.176 19.149 53.356 19.189 ;
      RECT MASK 1 53.84 19.149 54.02 19.189 ;
      RECT MASK 1 54.338 19.149 54.518 19.189 ;
      RECT MASK 1 55.002 19.149 55.182 19.189 ;
      RECT MASK 1 55.5 19.149 55.68 19.189 ;
      RECT MASK 1 56.164 19.149 56.344 19.189 ;
      RECT MASK 1 56.745 19.149 56.925 19.189 ;
      RECT MASK 1 58.051 19.149 58.231 19.189 ;
      RECT MASK 1 58.632 19.149 58.812 19.189 ;
      RECT MASK 1 59.296 19.149 59.476 19.189 ;
      RECT MASK 1 59.794 19.149 59.974 19.189 ;
      RECT MASK 1 60.458 19.149 60.638 19.189 ;
      RECT MASK 1 60.956 19.149 61.136 19.189 ;
      RECT MASK 1 61.62 19.149 61.8 19.189 ;
      RECT MASK 1 62.118 19.149 62.298 19.189 ;
      RECT MASK 1 62.782 19.149 62.962 19.189 ;
      RECT MASK 1 63.363 19.149 63.543 19.189 ;
      RECT MASK 1 64.669 19.149 64.849 19.189 ;
      RECT MASK 1 65.25 19.149 65.43 19.189 ;
      RECT MASK 1 65.914 19.149 66.094 19.189 ;
      RECT MASK 1 66.412 19.149 66.592 19.189 ;
      RECT MASK 1 67.076 19.149 67.256 19.189 ;
      RECT MASK 1 67.574 19.149 67.754 19.189 ;
      RECT MASK 1 68.238 19.149 68.418 19.189 ;
      RECT MASK 1 68.736 19.149 68.916 19.189 ;
      RECT MASK 1 69.4 19.149 69.58 19.189 ;
      RECT MASK 1 69.981 19.149 70.161 19.189 ;
      RECT MASK 1 71.287 19.149 71.467 19.189 ;
      RECT MASK 1 71.868 19.149 72.048 19.189 ;
      RECT MASK 1 72.532 19.149 72.712 19.189 ;
      RECT MASK 1 73.03 19.149 73.21 19.189 ;
      RECT MASK 1 73.694 19.149 73.874 19.189 ;
      RECT MASK 1 74.192 19.149 74.372 19.189 ;
      RECT MASK 1 74.856 19.149 75.036 19.189 ;
      RECT MASK 1 75.354 19.149 75.534 19.189 ;
      RECT MASK 1 76.018 19.149 76.198 19.189 ;
      RECT MASK 1 76.599 19.149 76.779 19.189 ;
      RECT MASK 1 77.905 19.149 78.085 19.189 ;
      RECT MASK 1 78.486 19.149 78.666 19.189 ;
      RECT MASK 1 79.15 19.149 79.33 19.189 ;
      RECT MASK 1 79.648 19.149 79.828 19.189 ;
      RECT MASK 1 80.312 19.149 80.492 19.189 ;
      RECT MASK 1 80.81 19.149 80.99 19.189 ;
      RECT MASK 1 81.474 19.149 81.654 19.189 ;
      RECT MASK 1 81.972 19.149 82.152 19.189 ;
      RECT MASK 1 82.636 19.149 82.816 19.189 ;
      RECT MASK 1 83.217 19.149 83.397 19.189 ;
      RECT MASK 1 84.523 19.149 84.703 19.189 ;
      RECT MASK 1 85.104 19.149 85.284 19.189 ;
      RECT MASK 1 85.768 19.149 85.948 19.189 ;
      RECT MASK 1 86.266 19.149 86.446 19.189 ;
      RECT MASK 1 86.93 19.149 87.11 19.189 ;
      RECT MASK 1 87.428 19.149 87.608 19.189 ;
      RECT MASK 1 88.092 19.149 88.272 19.189 ;
      RECT MASK 1 88.59 19.149 88.77 19.189 ;
      RECT MASK 1 89.254 19.149 89.434 19.189 ;
      RECT MASK 1 89.835 19.149 90.015 19.189 ;
      RECT MASK 1 91.141 19.149 91.321 19.189 ;
      RECT MASK 1 91.722 19.149 91.902 19.189 ;
      RECT MASK 1 92.386 19.149 92.566 19.189 ;
      RECT MASK 1 92.884 19.149 93.064 19.189 ;
      RECT MASK 1 93.548 19.149 93.728 19.189 ;
      RECT MASK 1 94.046 19.149 94.226 19.189 ;
      RECT MASK 1 94.71 19.149 94.89 19.189 ;
      RECT MASK 1 95.208 19.149 95.388 19.189 ;
      RECT MASK 1 95.872 19.149 96.052 19.189 ;
      RECT MASK 1 96.453 19.149 96.633 19.189 ;
      RECT MASK 1 97.759 19.149 97.939 19.189 ;
      RECT MASK 1 98.34 19.149 98.52 19.189 ;
      RECT MASK 1 99.004 19.149 99.184 19.189 ;
      RECT MASK 1 99.502 19.149 99.682 19.189 ;
      RECT MASK 1 100.166 19.149 100.346 19.189 ;
      RECT MASK 1 100.664 19.149 100.844 19.189 ;
      RECT MASK 1 101.328 19.149 101.508 19.189 ;
      RECT MASK 1 101.826 19.149 102.006 19.189 ;
      RECT MASK 1 102.49 19.149 102.67 19.189 ;
      RECT MASK 1 103.071 19.149 103.251 19.189 ;
      RECT MASK 1 104.377 19.149 104.557 19.189 ;
      RECT MASK 1 104.958 19.149 105.138 19.189 ;
      RECT MASK 1 105.622 19.149 105.802 19.189 ;
      RECT MASK 1 106.12 19.149 106.3 19.189 ;
      RECT MASK 1 106.784 19.149 106.964 19.189 ;
      RECT MASK 1 107.282 19.149 107.462 19.189 ;
      RECT MASK 1 107.946 19.149 108.126 19.189 ;
      RECT MASK 1 108.444 19.149 108.624 19.189 ;
      RECT MASK 1 109.108 19.149 109.288 19.189 ;
      RECT MASK 1 109.689 19.149 109.869 19.189 ;
      RECT MASK 1 1.406 19.165 4.69 19.205 ;
      RECT MASK 1 5.069 19.371 109.907 19.411 ;
      RECT MASK 1 1.431 19.4735 1.511 24.5065 ;
      RECT MASK 1 4.585 19.4735 4.665 24.5065 ;
      RECT MASK 1 5.889 19.75 6.498 19.79 ;
      RECT MASK 1 7.051 19.75 7.66 19.79 ;
      RECT MASK 1 8.213 19.75 8.822 19.79 ;
      RECT MASK 1 9.375 19.75 9.984 19.79 ;
      RECT MASK 1 12.507 19.75 13.116 19.79 ;
      RECT MASK 1 13.669 19.75 14.278 19.79 ;
      RECT MASK 1 14.831 19.75 15.44 19.79 ;
      RECT MASK 1 15.993 19.75 16.602 19.79 ;
      RECT MASK 1 19.125 19.75 19.734 19.79 ;
      RECT MASK 1 20.287 19.75 20.896 19.79 ;
      RECT MASK 1 21.449 19.75 22.058 19.79 ;
      RECT MASK 1 22.611 19.75 23.22 19.79 ;
      RECT MASK 1 25.743 19.75 26.352 19.79 ;
      RECT MASK 1 26.905 19.75 27.514 19.79 ;
      RECT MASK 1 28.067 19.75 28.676 19.79 ;
      RECT MASK 1 29.229 19.75 29.838 19.79 ;
      RECT MASK 1 32.361 19.75 32.97 19.79 ;
      RECT MASK 1 33.523 19.75 34.132 19.79 ;
      RECT MASK 1 34.685 19.75 35.294 19.79 ;
      RECT MASK 1 35.847 19.75 36.456 19.79 ;
      RECT MASK 1 38.979 19.75 39.588 19.79 ;
      RECT MASK 1 40.141 19.75 40.75 19.79 ;
      RECT MASK 1 41.303 19.75 41.912 19.79 ;
      RECT MASK 1 42.465 19.75 43.074 19.79 ;
      RECT MASK 1 45.597 19.75 46.206 19.79 ;
      RECT MASK 1 46.759 19.75 47.368 19.79 ;
      RECT MASK 1 47.921 19.75 48.53 19.79 ;
      RECT MASK 1 49.083 19.75 49.692 19.79 ;
      RECT MASK 1 52.215 19.75 52.824 19.79 ;
      RECT MASK 1 53.377 19.75 53.986 19.79 ;
      RECT MASK 1 54.539 19.75 55.148 19.79 ;
      RECT MASK 1 55.701 19.75 56.31 19.79 ;
      RECT MASK 1 58.833 19.75 59.442 19.79 ;
      RECT MASK 1 59.995 19.75 60.604 19.79 ;
      RECT MASK 1 61.157 19.75 61.766 19.79 ;
      RECT MASK 1 62.319 19.75 62.928 19.79 ;
      RECT MASK 1 65.451 19.75 66.06 19.79 ;
      RECT MASK 1 66.613 19.75 67.222 19.79 ;
      RECT MASK 1 67.775 19.75 68.384 19.79 ;
      RECT MASK 1 68.937 19.75 69.546 19.79 ;
      RECT MASK 1 72.069 19.75 72.678 19.79 ;
      RECT MASK 1 73.231 19.75 73.84 19.79 ;
      RECT MASK 1 74.393 19.75 75.002 19.79 ;
      RECT MASK 1 75.555 19.75 76.164 19.79 ;
      RECT MASK 1 78.687 19.75 79.296 19.79 ;
      RECT MASK 1 79.849 19.75 80.458 19.79 ;
      RECT MASK 1 81.011 19.75 81.62 19.79 ;
      RECT MASK 1 82.173 19.75 82.782 19.79 ;
      RECT MASK 1 85.305 19.75 85.914 19.79 ;
      RECT MASK 1 86.467 19.75 87.076 19.79 ;
      RECT MASK 1 87.629 19.75 88.238 19.79 ;
      RECT MASK 1 88.791 19.75 89.4 19.79 ;
      RECT MASK 1 91.923 19.75 92.532 19.79 ;
      RECT MASK 1 93.085 19.75 93.694 19.79 ;
      RECT MASK 1 94.247 19.75 94.856 19.79 ;
      RECT MASK 1 95.409 19.75 96.018 19.79 ;
      RECT MASK 1 98.541 19.75 99.15 19.79 ;
      RECT MASK 1 99.703 19.75 100.312 19.79 ;
      RECT MASK 1 100.865 19.75 101.474 19.79 ;
      RECT MASK 1 102.027 19.75 102.636 19.79 ;
      RECT MASK 1 105.159 19.75 105.768 19.79 ;
      RECT MASK 1 106.321 19.75 106.93 19.79 ;
      RECT MASK 1 107.483 19.75 108.092 19.79 ;
      RECT MASK 1 108.645 19.75 109.254 19.79 ;
      RECT MASK 1 2.225 19.77 2.285 20.82 ;
      RECT MASK 1 2.499 19.77 2.559 20.82 ;
      RECT MASK 1 2.773 19.77 2.833 20.82 ;
      RECT MASK 1 3.047 19.77 3.107 20.82 ;
      RECT MASK 1 3.321 19.77 3.381 20.82 ;
      RECT MASK 1 3.595 19.77 3.655 20.82 ;
      RECT MASK 1 3.869 19.77 3.929 20.82 ;
      RECT MASK 1 5.031 19.831 5.695 19.871 ;
      RECT MASK 1 10.177 19.831 10.675 19.871 ;
      RECT MASK 1 11.649 19.831 12.313 19.871 ;
      RECT MASK 1 16.795 19.831 17.293 19.871 ;
      RECT MASK 1 18.267 19.831 18.931 19.871 ;
      RECT MASK 1 23.413 19.831 23.911 19.871 ;
      RECT MASK 1 24.885 19.831 25.549 19.871 ;
      RECT MASK 1 30.031 19.831 30.529 19.871 ;
      RECT MASK 1 31.503 19.831 32.167 19.871 ;
      RECT MASK 1 36.649 19.831 37.147 19.871 ;
      RECT MASK 1 38.121 19.831 38.785 19.871 ;
      RECT MASK 1 43.267 19.831 43.765 19.871 ;
      RECT MASK 1 44.739 19.831 45.403 19.871 ;
      RECT MASK 1 49.885 19.831 50.383 19.871 ;
      RECT MASK 1 51.357 19.831 52.021 19.871 ;
      RECT MASK 1 56.503 19.831 57.001 19.871 ;
      RECT MASK 1 57.975 19.831 58.639 19.871 ;
      RECT MASK 1 63.121 19.831 63.619 19.871 ;
      RECT MASK 1 64.593 19.831 65.257 19.871 ;
      RECT MASK 1 69.739 19.831 70.237 19.871 ;
      RECT MASK 1 71.211 19.831 71.875 19.871 ;
      RECT MASK 1 76.357 19.831 76.855 19.871 ;
      RECT MASK 1 77.829 19.831 78.493 19.871 ;
      RECT MASK 1 82.975 19.831 83.473 19.871 ;
      RECT MASK 1 84.447 19.831 85.111 19.871 ;
      RECT MASK 1 89.593 19.831 90.091 19.871 ;
      RECT MASK 1 91.065 19.831 91.729 19.871 ;
      RECT MASK 1 96.211 19.831 96.709 19.871 ;
      RECT MASK 1 97.683 19.831 98.347 19.871 ;
      RECT MASK 1 102.829 19.831 103.327 19.871 ;
      RECT MASK 1 104.301 19.831 104.965 19.871 ;
      RECT MASK 1 109.447 19.831 109.945 19.871 ;
      RECT MASK 1 5.031 20.099 109.945 20.139 ;
      RECT MASK 1 5.688 20.321 5.868 20.361 ;
      RECT MASK 1 6.352 20.321 6.532 20.361 ;
      RECT MASK 1 6.85 20.321 7.03 20.361 ;
      RECT MASK 1 7.514 20.321 7.694 20.361 ;
      RECT MASK 1 8.012 20.321 8.192 20.361 ;
      RECT MASK 1 8.676 20.321 8.856 20.361 ;
      RECT MASK 1 9.174 20.321 9.354 20.361 ;
      RECT MASK 1 9.838 20.321 10.018 20.361 ;
      RECT MASK 1 12.306 20.321 12.486 20.361 ;
      RECT MASK 1 12.97 20.321 13.15 20.361 ;
      RECT MASK 1 13.468 20.321 13.648 20.361 ;
      RECT MASK 1 14.132 20.321 14.312 20.361 ;
      RECT MASK 1 14.63 20.321 14.81 20.361 ;
      RECT MASK 1 15.294 20.321 15.474 20.361 ;
      RECT MASK 1 15.792 20.321 15.972 20.361 ;
      RECT MASK 1 16.456 20.321 16.636 20.361 ;
      RECT MASK 1 18.924 20.321 19.104 20.361 ;
      RECT MASK 1 19.588 20.321 19.768 20.361 ;
      RECT MASK 1 20.086 20.321 20.266 20.361 ;
      RECT MASK 1 20.75 20.321 20.93 20.361 ;
      RECT MASK 1 21.248 20.321 21.428 20.361 ;
      RECT MASK 1 21.912 20.321 22.092 20.361 ;
      RECT MASK 1 22.41 20.321 22.59 20.361 ;
      RECT MASK 1 23.074 20.321 23.254 20.361 ;
      RECT MASK 1 25.542 20.321 25.722 20.361 ;
      RECT MASK 1 26.206 20.321 26.386 20.361 ;
      RECT MASK 1 26.704 20.321 26.884 20.361 ;
      RECT MASK 1 27.368 20.321 27.548 20.361 ;
      RECT MASK 1 27.866 20.321 28.046 20.361 ;
      RECT MASK 1 28.53 20.321 28.71 20.361 ;
      RECT MASK 1 29.028 20.321 29.208 20.361 ;
      RECT MASK 1 29.692 20.321 29.872 20.361 ;
      RECT MASK 1 32.16 20.321 32.34 20.361 ;
      RECT MASK 1 32.824 20.321 33.004 20.361 ;
      RECT MASK 1 33.322 20.321 33.502 20.361 ;
      RECT MASK 1 33.986 20.321 34.166 20.361 ;
      RECT MASK 1 34.484 20.321 34.664 20.361 ;
      RECT MASK 1 35.148 20.321 35.328 20.361 ;
      RECT MASK 1 35.646 20.321 35.826 20.361 ;
      RECT MASK 1 36.31 20.321 36.49 20.361 ;
      RECT MASK 1 38.778 20.321 38.958 20.361 ;
      RECT MASK 1 39.442 20.321 39.622 20.361 ;
      RECT MASK 1 39.94 20.321 40.12 20.361 ;
      RECT MASK 1 40.604 20.321 40.784 20.361 ;
      RECT MASK 1 41.102 20.321 41.282 20.361 ;
      RECT MASK 1 41.766 20.321 41.946 20.361 ;
      RECT MASK 1 42.264 20.321 42.444 20.361 ;
      RECT MASK 1 42.928 20.321 43.108 20.361 ;
      RECT MASK 1 45.396 20.321 45.576 20.361 ;
      RECT MASK 1 46.06 20.321 46.24 20.361 ;
      RECT MASK 1 46.558 20.321 46.738 20.361 ;
      RECT MASK 1 47.222 20.321 47.402 20.361 ;
      RECT MASK 1 47.72 20.321 47.9 20.361 ;
      RECT MASK 1 48.384 20.321 48.564 20.361 ;
      RECT MASK 1 48.882 20.321 49.062 20.361 ;
      RECT MASK 1 49.546 20.321 49.726 20.361 ;
      RECT MASK 1 52.014 20.321 52.194 20.361 ;
      RECT MASK 1 52.678 20.321 52.858 20.361 ;
      RECT MASK 1 53.176 20.321 53.356 20.361 ;
      RECT MASK 1 53.84 20.321 54.02 20.361 ;
      RECT MASK 1 54.338 20.321 54.518 20.361 ;
      RECT MASK 1 55.002 20.321 55.182 20.361 ;
      RECT MASK 1 55.5 20.321 55.68 20.361 ;
      RECT MASK 1 56.164 20.321 56.344 20.361 ;
      RECT MASK 1 58.632 20.321 58.812 20.361 ;
      RECT MASK 1 59.296 20.321 59.476 20.361 ;
      RECT MASK 1 59.794 20.321 59.974 20.361 ;
      RECT MASK 1 60.458 20.321 60.638 20.361 ;
      RECT MASK 1 60.956 20.321 61.136 20.361 ;
      RECT MASK 1 61.62 20.321 61.8 20.361 ;
      RECT MASK 1 62.118 20.321 62.298 20.361 ;
      RECT MASK 1 62.782 20.321 62.962 20.361 ;
      RECT MASK 1 65.25 20.321 65.43 20.361 ;
      RECT MASK 1 65.914 20.321 66.094 20.361 ;
      RECT MASK 1 66.412 20.321 66.592 20.361 ;
      RECT MASK 1 67.076 20.321 67.256 20.361 ;
      RECT MASK 1 67.574 20.321 67.754 20.361 ;
      RECT MASK 1 68.238 20.321 68.418 20.361 ;
      RECT MASK 1 68.736 20.321 68.916 20.361 ;
      RECT MASK 1 69.4 20.321 69.58 20.361 ;
      RECT MASK 1 71.868 20.321 72.048 20.361 ;
      RECT MASK 1 72.532 20.321 72.712 20.361 ;
      RECT MASK 1 73.03 20.321 73.21 20.361 ;
      RECT MASK 1 73.694 20.321 73.874 20.361 ;
      RECT MASK 1 74.192 20.321 74.372 20.361 ;
      RECT MASK 1 74.856 20.321 75.036 20.361 ;
      RECT MASK 1 75.354 20.321 75.534 20.361 ;
      RECT MASK 1 76.018 20.321 76.198 20.361 ;
      RECT MASK 1 78.486 20.321 78.666 20.361 ;
      RECT MASK 1 79.15 20.321 79.33 20.361 ;
      RECT MASK 1 79.648 20.321 79.828 20.361 ;
      RECT MASK 1 80.312 20.321 80.492 20.361 ;
      RECT MASK 1 80.81 20.321 80.99 20.361 ;
      RECT MASK 1 81.474 20.321 81.654 20.361 ;
      RECT MASK 1 81.972 20.321 82.152 20.361 ;
      RECT MASK 1 82.636 20.321 82.816 20.361 ;
      RECT MASK 1 85.104 20.321 85.284 20.361 ;
      RECT MASK 1 85.768 20.321 85.948 20.361 ;
      RECT MASK 1 86.266 20.321 86.446 20.361 ;
      RECT MASK 1 86.93 20.321 87.11 20.361 ;
      RECT MASK 1 87.428 20.321 87.608 20.361 ;
      RECT MASK 1 88.092 20.321 88.272 20.361 ;
      RECT MASK 1 88.59 20.321 88.77 20.361 ;
      RECT MASK 1 89.254 20.321 89.434 20.361 ;
      RECT MASK 1 91.722 20.321 91.902 20.361 ;
      RECT MASK 1 92.386 20.321 92.566 20.361 ;
      RECT MASK 1 92.884 20.321 93.064 20.361 ;
      RECT MASK 1 93.548 20.321 93.728 20.361 ;
      RECT MASK 1 94.046 20.321 94.226 20.361 ;
      RECT MASK 1 94.71 20.321 94.89 20.361 ;
      RECT MASK 1 95.208 20.321 95.388 20.361 ;
      RECT MASK 1 95.872 20.321 96.052 20.361 ;
      RECT MASK 1 98.34 20.321 98.52 20.361 ;
      RECT MASK 1 99.004 20.321 99.184 20.361 ;
      RECT MASK 1 99.502 20.321 99.682 20.361 ;
      RECT MASK 1 100.166 20.321 100.346 20.361 ;
      RECT MASK 1 100.664 20.321 100.844 20.361 ;
      RECT MASK 1 101.328 20.321 101.508 20.361 ;
      RECT MASK 1 101.826 20.321 102.006 20.361 ;
      RECT MASK 1 102.49 20.321 102.67 20.361 ;
      RECT MASK 1 104.958 20.321 105.138 20.361 ;
      RECT MASK 1 105.622 20.321 105.802 20.361 ;
      RECT MASK 1 106.12 20.321 106.3 20.361 ;
      RECT MASK 1 106.784 20.321 106.964 20.361 ;
      RECT MASK 1 107.282 20.321 107.462 20.361 ;
      RECT MASK 1 107.946 20.321 108.126 20.361 ;
      RECT MASK 1 108.444 20.321 108.624 20.361 ;
      RECT MASK 1 109.108 20.321 109.288 20.361 ;
      RECT MASK 1 5.107 20.357 5.287 20.397 ;
      RECT MASK 1 10.419 20.357 10.599 20.397 ;
      RECT MASK 1 11.725 20.357 11.905 20.397 ;
      RECT MASK 1 17.037 20.357 17.217 20.397 ;
      RECT MASK 1 18.343 20.357 18.523 20.397 ;
      RECT MASK 1 23.655 20.357 23.835 20.397 ;
      RECT MASK 1 24.961 20.357 25.141 20.397 ;
      RECT MASK 1 30.273 20.357 30.453 20.397 ;
      RECT MASK 1 31.579 20.357 31.759 20.397 ;
      RECT MASK 1 36.891 20.357 37.071 20.397 ;
      RECT MASK 1 38.197 20.357 38.377 20.397 ;
      RECT MASK 1 43.509 20.357 43.689 20.397 ;
      RECT MASK 1 44.815 20.357 44.995 20.397 ;
      RECT MASK 1 50.127 20.357 50.307 20.397 ;
      RECT MASK 1 51.433 20.357 51.613 20.397 ;
      RECT MASK 1 56.745 20.357 56.925 20.397 ;
      RECT MASK 1 58.051 20.357 58.231 20.397 ;
      RECT MASK 1 63.363 20.357 63.543 20.397 ;
      RECT MASK 1 64.669 20.357 64.849 20.397 ;
      RECT MASK 1 69.981 20.357 70.161 20.397 ;
      RECT MASK 1 71.287 20.357 71.467 20.397 ;
      RECT MASK 1 76.599 20.357 76.779 20.397 ;
      RECT MASK 1 77.905 20.357 78.085 20.397 ;
      RECT MASK 1 83.217 20.357 83.397 20.397 ;
      RECT MASK 1 84.523 20.357 84.703 20.397 ;
      RECT MASK 1 89.835 20.357 90.015 20.397 ;
      RECT MASK 1 91.141 20.357 91.321 20.397 ;
      RECT MASK 1 96.453 20.357 96.633 20.397 ;
      RECT MASK 1 97.759 20.357 97.939 20.397 ;
      RECT MASK 1 103.071 20.357 103.251 20.397 ;
      RECT MASK 1 104.377 20.357 104.557 20.397 ;
      RECT MASK 1 109.689 20.357 109.869 20.397 ;
      RECT MASK 1 5.107 20.525 5.287 20.565 ;
      RECT MASK 1 10.419 20.525 10.599 20.565 ;
      RECT MASK 1 11.725 20.525 11.905 20.565 ;
      RECT MASK 1 17.037 20.525 17.217 20.565 ;
      RECT MASK 1 18.343 20.525 18.523 20.565 ;
      RECT MASK 1 23.655 20.525 23.835 20.565 ;
      RECT MASK 1 24.961 20.525 25.141 20.565 ;
      RECT MASK 1 30.273 20.525 30.453 20.565 ;
      RECT MASK 1 31.579 20.525 31.759 20.565 ;
      RECT MASK 1 36.891 20.525 37.071 20.565 ;
      RECT MASK 1 38.197 20.525 38.377 20.565 ;
      RECT MASK 1 43.509 20.525 43.689 20.565 ;
      RECT MASK 1 44.815 20.525 44.995 20.565 ;
      RECT MASK 1 50.127 20.525 50.307 20.565 ;
      RECT MASK 1 51.433 20.525 51.613 20.565 ;
      RECT MASK 1 56.745 20.525 56.925 20.565 ;
      RECT MASK 1 58.051 20.525 58.231 20.565 ;
      RECT MASK 1 63.363 20.525 63.543 20.565 ;
      RECT MASK 1 64.669 20.525 64.849 20.565 ;
      RECT MASK 1 69.981 20.525 70.161 20.565 ;
      RECT MASK 1 71.287 20.525 71.467 20.565 ;
      RECT MASK 1 76.599 20.525 76.779 20.565 ;
      RECT MASK 1 77.905 20.525 78.085 20.565 ;
      RECT MASK 1 83.217 20.525 83.397 20.565 ;
      RECT MASK 1 84.523 20.525 84.703 20.565 ;
      RECT MASK 1 89.835 20.525 90.015 20.565 ;
      RECT MASK 1 91.141 20.525 91.321 20.565 ;
      RECT MASK 1 96.453 20.525 96.633 20.565 ;
      RECT MASK 1 97.759 20.525 97.939 20.565 ;
      RECT MASK 1 103.071 20.525 103.251 20.565 ;
      RECT MASK 1 104.377 20.525 104.557 20.565 ;
      RECT MASK 1 109.689 20.525 109.869 20.565 ;
      RECT MASK 1 5.816 20.543 5.999 20.583 ;
      RECT MASK 1 6.221 20.543 6.404 20.583 ;
      RECT MASK 1 6.978 20.543 7.161 20.583 ;
      RECT MASK 1 7.383 20.543 7.566 20.583 ;
      RECT MASK 1 8.14 20.543 8.323 20.583 ;
      RECT MASK 1 8.545 20.543 8.728 20.583 ;
      RECT MASK 1 9.302 20.543 9.485 20.583 ;
      RECT MASK 1 9.707 20.543 9.89 20.583 ;
      RECT MASK 1 12.434 20.543 12.617 20.583 ;
      RECT MASK 1 12.839 20.543 13.022 20.583 ;
      RECT MASK 1 13.596 20.543 13.779 20.583 ;
      RECT MASK 1 14.001 20.543 14.184 20.583 ;
      RECT MASK 1 14.758 20.543 14.941 20.583 ;
      RECT MASK 1 15.163 20.543 15.346 20.583 ;
      RECT MASK 1 15.92 20.543 16.103 20.583 ;
      RECT MASK 1 16.325 20.543 16.508 20.583 ;
      RECT MASK 1 19.052 20.543 19.235 20.583 ;
      RECT MASK 1 19.457 20.543 19.64 20.583 ;
      RECT MASK 1 20.214 20.543 20.397 20.583 ;
      RECT MASK 1 20.619 20.543 20.802 20.583 ;
      RECT MASK 1 21.376 20.543 21.559 20.583 ;
      RECT MASK 1 21.781 20.543 21.964 20.583 ;
      RECT MASK 1 22.538 20.543 22.721 20.583 ;
      RECT MASK 1 22.943 20.543 23.126 20.583 ;
      RECT MASK 1 25.67 20.543 25.853 20.583 ;
      RECT MASK 1 26.075 20.543 26.258 20.583 ;
      RECT MASK 1 26.832 20.543 27.015 20.583 ;
      RECT MASK 1 27.237 20.543 27.42 20.583 ;
      RECT MASK 1 27.994 20.543 28.177 20.583 ;
      RECT MASK 1 28.399 20.543 28.582 20.583 ;
      RECT MASK 1 29.156 20.543 29.339 20.583 ;
      RECT MASK 1 29.561 20.543 29.744 20.583 ;
      RECT MASK 1 32.288 20.543 32.471 20.583 ;
      RECT MASK 1 32.693 20.543 32.876 20.583 ;
      RECT MASK 1 33.45 20.543 33.633 20.583 ;
      RECT MASK 1 33.855 20.543 34.038 20.583 ;
      RECT MASK 1 34.612 20.543 34.795 20.583 ;
      RECT MASK 1 35.017 20.543 35.2 20.583 ;
      RECT MASK 1 35.774 20.543 35.957 20.583 ;
      RECT MASK 1 36.179 20.543 36.362 20.583 ;
      RECT MASK 1 38.906 20.543 39.089 20.583 ;
      RECT MASK 1 39.311 20.543 39.494 20.583 ;
      RECT MASK 1 40.068 20.543 40.251 20.583 ;
      RECT MASK 1 40.473 20.543 40.656 20.583 ;
      RECT MASK 1 41.23 20.543 41.413 20.583 ;
      RECT MASK 1 41.635 20.543 41.818 20.583 ;
      RECT MASK 1 42.392 20.543 42.575 20.583 ;
      RECT MASK 1 42.797 20.543 42.98 20.583 ;
      RECT MASK 1 45.524 20.543 45.707 20.583 ;
      RECT MASK 1 45.929 20.543 46.112 20.583 ;
      RECT MASK 1 46.686 20.543 46.869 20.583 ;
      RECT MASK 1 47.091 20.543 47.274 20.583 ;
      RECT MASK 1 47.848 20.543 48.031 20.583 ;
      RECT MASK 1 48.253 20.543 48.436 20.583 ;
      RECT MASK 1 49.01 20.543 49.193 20.583 ;
      RECT MASK 1 49.415 20.543 49.598 20.583 ;
      RECT MASK 1 52.142 20.543 52.325 20.583 ;
      RECT MASK 1 52.547 20.543 52.73 20.583 ;
      RECT MASK 1 53.304 20.543 53.487 20.583 ;
      RECT MASK 1 53.709 20.543 53.892 20.583 ;
      RECT MASK 1 54.466 20.543 54.649 20.583 ;
      RECT MASK 1 54.871 20.543 55.054 20.583 ;
      RECT MASK 1 55.628 20.543 55.811 20.583 ;
      RECT MASK 1 56.033 20.543 56.216 20.583 ;
      RECT MASK 1 58.76 20.543 58.943 20.583 ;
      RECT MASK 1 59.165 20.543 59.348 20.583 ;
      RECT MASK 1 59.922 20.543 60.105 20.583 ;
      RECT MASK 1 60.327 20.543 60.51 20.583 ;
      RECT MASK 1 61.084 20.543 61.267 20.583 ;
      RECT MASK 1 61.489 20.543 61.672 20.583 ;
      RECT MASK 1 62.246 20.543 62.429 20.583 ;
      RECT MASK 1 62.651 20.543 62.834 20.583 ;
      RECT MASK 1 65.378 20.543 65.561 20.583 ;
      RECT MASK 1 65.783 20.543 65.966 20.583 ;
      RECT MASK 1 66.54 20.543 66.723 20.583 ;
      RECT MASK 1 66.945 20.543 67.128 20.583 ;
      RECT MASK 1 67.702 20.543 67.885 20.583 ;
      RECT MASK 1 68.107 20.543 68.29 20.583 ;
      RECT MASK 1 68.864 20.543 69.047 20.583 ;
      RECT MASK 1 69.269 20.543 69.452 20.583 ;
      RECT MASK 1 71.996 20.543 72.179 20.583 ;
      RECT MASK 1 72.401 20.543 72.584 20.583 ;
      RECT MASK 1 73.158 20.543 73.341 20.583 ;
      RECT MASK 1 73.563 20.543 73.746 20.583 ;
      RECT MASK 1 74.32 20.543 74.503 20.583 ;
      RECT MASK 1 74.725 20.543 74.908 20.583 ;
      RECT MASK 1 75.482 20.543 75.665 20.583 ;
      RECT MASK 1 75.887 20.543 76.07 20.583 ;
      RECT MASK 1 78.614 20.543 78.797 20.583 ;
      RECT MASK 1 79.019 20.543 79.202 20.583 ;
      RECT MASK 1 79.776 20.543 79.959 20.583 ;
      RECT MASK 1 80.181 20.543 80.364 20.583 ;
      RECT MASK 1 80.938 20.543 81.121 20.583 ;
      RECT MASK 1 81.343 20.543 81.526 20.583 ;
      RECT MASK 1 82.1 20.543 82.283 20.583 ;
      RECT MASK 1 82.505 20.543 82.688 20.583 ;
      RECT MASK 1 85.232 20.543 85.415 20.583 ;
      RECT MASK 1 85.637 20.543 85.82 20.583 ;
      RECT MASK 1 86.394 20.543 86.577 20.583 ;
      RECT MASK 1 86.799 20.543 86.982 20.583 ;
      RECT MASK 1 87.556 20.543 87.739 20.583 ;
      RECT MASK 1 87.961 20.543 88.144 20.583 ;
      RECT MASK 1 88.718 20.543 88.901 20.583 ;
      RECT MASK 1 89.123 20.543 89.306 20.583 ;
      RECT MASK 1 91.85 20.543 92.033 20.583 ;
      RECT MASK 1 92.255 20.543 92.438 20.583 ;
      RECT MASK 1 93.012 20.543 93.195 20.583 ;
      RECT MASK 1 93.417 20.543 93.6 20.583 ;
      RECT MASK 1 94.174 20.543 94.357 20.583 ;
      RECT MASK 1 94.579 20.543 94.762 20.583 ;
      RECT MASK 1 95.336 20.543 95.519 20.583 ;
      RECT MASK 1 95.741 20.543 95.924 20.583 ;
      RECT MASK 1 98.468 20.543 98.651 20.583 ;
      RECT MASK 1 98.873 20.543 99.056 20.583 ;
      RECT MASK 1 99.63 20.543 99.813 20.583 ;
      RECT MASK 1 100.035 20.543 100.218 20.583 ;
      RECT MASK 1 100.792 20.543 100.975 20.583 ;
      RECT MASK 1 101.197 20.543 101.38 20.583 ;
      RECT MASK 1 101.954 20.543 102.137 20.583 ;
      RECT MASK 1 102.359 20.543 102.542 20.583 ;
      RECT MASK 1 105.086 20.543 105.269 20.583 ;
      RECT MASK 1 105.491 20.543 105.674 20.583 ;
      RECT MASK 1 106.248 20.543 106.431 20.583 ;
      RECT MASK 1 106.653 20.543 106.836 20.583 ;
      RECT MASK 1 107.41 20.543 107.593 20.583 ;
      RECT MASK 1 107.815 20.543 107.998 20.583 ;
      RECT MASK 1 108.572 20.543 108.755 20.583 ;
      RECT MASK 1 108.977 20.543 109.16 20.583 ;
      RECT MASK 1 116.154 20.7 116.214 21.75 ;
      RECT MASK 1 116.428 20.7 116.488 21.75 ;
      RECT MASK 1 116.702 20.7 116.762 21.75 ;
      RECT MASK 1 116.976 20.7 117.036 21.75 ;
      RECT MASK 1 117.25 20.7 117.31 21.75 ;
      RECT MASK 1 117.524 20.7 117.584 21.75 ;
      RECT MASK 1 117.798 20.7 117.858 21.75 ;
      RECT MASK 1 118.072 20.7 118.132 21.75 ;
      RECT MASK 1 118.346 20.7 118.406 21.75 ;
      RECT MASK 1 118.62 20.7 118.68 21.75 ;
      RECT MASK 1 118.894 20.7 118.954 21.75 ;
      RECT MASK 1 119.168 20.7 119.228 21.75 ;
      RECT MASK 1 119.442 20.7 119.502 21.75 ;
      RECT MASK 1 119.716 20.7 119.776 21.75 ;
      RECT MASK 1 119.99 20.7 120.05 21.75 ;
      RECT MASK 1 120.264 20.7 120.324 21.75 ;
      RECT MASK 1 120.538 20.7 120.598 21.75 ;
      RECT MASK 1 120.812 20.7 120.872 21.75 ;
      RECT MASK 1 121.086 20.7 121.146 21.75 ;
      RECT MASK 1 121.36 20.7 121.42 21.75 ;
      RECT MASK 1 121.634 20.7 121.694 21.75 ;
      RECT MASK 1 121.908 20.7 121.968 21.75 ;
      RECT MASK 1 122.182 20.7 122.242 21.75 ;
      RECT MASK 1 122.456 20.7 122.516 21.75 ;
      RECT MASK 1 122.73 20.7 122.79 21.75 ;
      RECT MASK 1 123.004 20.7 123.064 21.75 ;
      RECT MASK 1 123.278 20.7 123.338 21.75 ;
      RECT MASK 1 123.552 20.7 123.612 21.75 ;
      RECT MASK 1 123.826 20.7 123.886 21.75 ;
      RECT MASK 1 124.1 20.7 124.16 21.75 ;
      RECT MASK 1 124.374 20.7 124.434 21.75 ;
      RECT MASK 1 124.648 20.7 124.708 21.75 ;
      RECT MASK 1 124.922 20.7 124.982 21.75 ;
      RECT MASK 1 125.196 20.7 125.256 21.75 ;
      RECT MASK 1 125.47 20.7 125.53 21.75 ;
      RECT MASK 1 125.744 20.7 125.804 21.75 ;
      RECT MASK 1 126.018 20.7 126.078 21.75 ;
      RECT MASK 1 126.292 20.7 126.352 21.75 ;
      RECT MASK 1 126.566 20.7 126.626 21.75 ;
      RECT MASK 1 126.84 20.7 126.9 21.75 ;
      RECT MASK 1 127.114 20.7 127.174 21.75 ;
      RECT MASK 1 127.388 20.7 127.448 21.75 ;
      RECT MASK 1 127.662 20.7 127.722 21.75 ;
      RECT MASK 1 127.936 20.7 127.996 21.75 ;
      RECT MASK 1 128.21 20.7 128.27 21.75 ;
      RECT MASK 1 5.816 20.711 5.999 20.751 ;
      RECT MASK 1 6.221 20.711 6.404 20.751 ;
      RECT MASK 1 6.978 20.711 7.161 20.751 ;
      RECT MASK 1 7.383 20.711 7.566 20.751 ;
      RECT MASK 1 8.14 20.711 8.323 20.751 ;
      RECT MASK 1 8.545 20.711 8.728 20.751 ;
      RECT MASK 1 9.302 20.711 9.485 20.751 ;
      RECT MASK 1 9.707 20.711 9.89 20.751 ;
      RECT MASK 1 12.434 20.711 12.617 20.751 ;
      RECT MASK 1 12.839 20.711 13.022 20.751 ;
      RECT MASK 1 13.596 20.711 13.779 20.751 ;
      RECT MASK 1 14.001 20.711 14.184 20.751 ;
      RECT MASK 1 14.758 20.711 14.941 20.751 ;
      RECT MASK 1 15.163 20.711 15.346 20.751 ;
      RECT MASK 1 15.92 20.711 16.103 20.751 ;
      RECT MASK 1 16.325 20.711 16.508 20.751 ;
      RECT MASK 1 19.052 20.711 19.235 20.751 ;
      RECT MASK 1 19.457 20.711 19.64 20.751 ;
      RECT MASK 1 20.214 20.711 20.397 20.751 ;
      RECT MASK 1 20.619 20.711 20.802 20.751 ;
      RECT MASK 1 21.376 20.711 21.559 20.751 ;
      RECT MASK 1 21.781 20.711 21.964 20.751 ;
      RECT MASK 1 22.538 20.711 22.721 20.751 ;
      RECT MASK 1 22.943 20.711 23.126 20.751 ;
      RECT MASK 1 25.67 20.711 25.853 20.751 ;
      RECT MASK 1 26.075 20.711 26.258 20.751 ;
      RECT MASK 1 26.832 20.711 27.015 20.751 ;
      RECT MASK 1 27.237 20.711 27.42 20.751 ;
      RECT MASK 1 27.994 20.711 28.177 20.751 ;
      RECT MASK 1 28.399 20.711 28.582 20.751 ;
      RECT MASK 1 29.156 20.711 29.339 20.751 ;
      RECT MASK 1 29.561 20.711 29.744 20.751 ;
      RECT MASK 1 32.288 20.711 32.471 20.751 ;
      RECT MASK 1 32.693 20.711 32.876 20.751 ;
      RECT MASK 1 33.45 20.711 33.633 20.751 ;
      RECT MASK 1 33.855 20.711 34.038 20.751 ;
      RECT MASK 1 34.612 20.711 34.795 20.751 ;
      RECT MASK 1 35.017 20.711 35.2 20.751 ;
      RECT MASK 1 35.774 20.711 35.957 20.751 ;
      RECT MASK 1 36.179 20.711 36.362 20.751 ;
      RECT MASK 1 38.906 20.711 39.089 20.751 ;
      RECT MASK 1 39.311 20.711 39.494 20.751 ;
      RECT MASK 1 40.068 20.711 40.251 20.751 ;
      RECT MASK 1 40.473 20.711 40.656 20.751 ;
      RECT MASK 1 41.23 20.711 41.413 20.751 ;
      RECT MASK 1 41.635 20.711 41.818 20.751 ;
      RECT MASK 1 42.392 20.711 42.575 20.751 ;
      RECT MASK 1 42.797 20.711 42.98 20.751 ;
      RECT MASK 1 45.524 20.711 45.707 20.751 ;
      RECT MASK 1 45.929 20.711 46.112 20.751 ;
      RECT MASK 1 46.686 20.711 46.869 20.751 ;
      RECT MASK 1 47.091 20.711 47.274 20.751 ;
      RECT MASK 1 47.848 20.711 48.031 20.751 ;
      RECT MASK 1 48.253 20.711 48.436 20.751 ;
      RECT MASK 1 49.01 20.711 49.193 20.751 ;
      RECT MASK 1 49.415 20.711 49.598 20.751 ;
      RECT MASK 1 52.142 20.711 52.325 20.751 ;
      RECT MASK 1 52.547 20.711 52.73 20.751 ;
      RECT MASK 1 53.304 20.711 53.487 20.751 ;
      RECT MASK 1 53.709 20.711 53.892 20.751 ;
      RECT MASK 1 54.466 20.711 54.649 20.751 ;
      RECT MASK 1 54.871 20.711 55.054 20.751 ;
      RECT MASK 1 55.628 20.711 55.811 20.751 ;
      RECT MASK 1 56.033 20.711 56.216 20.751 ;
      RECT MASK 1 58.76 20.711 58.943 20.751 ;
      RECT MASK 1 59.165 20.711 59.348 20.751 ;
      RECT MASK 1 59.922 20.711 60.105 20.751 ;
      RECT MASK 1 60.327 20.711 60.51 20.751 ;
      RECT MASK 1 61.084 20.711 61.267 20.751 ;
      RECT MASK 1 61.489 20.711 61.672 20.751 ;
      RECT MASK 1 62.246 20.711 62.429 20.751 ;
      RECT MASK 1 62.651 20.711 62.834 20.751 ;
      RECT MASK 1 65.378 20.711 65.561 20.751 ;
      RECT MASK 1 65.783 20.711 65.966 20.751 ;
      RECT MASK 1 66.54 20.711 66.723 20.751 ;
      RECT MASK 1 66.945 20.711 67.128 20.751 ;
      RECT MASK 1 67.702 20.711 67.885 20.751 ;
      RECT MASK 1 68.107 20.711 68.29 20.751 ;
      RECT MASK 1 68.864 20.711 69.047 20.751 ;
      RECT MASK 1 69.269 20.711 69.452 20.751 ;
      RECT MASK 1 71.996 20.711 72.179 20.751 ;
      RECT MASK 1 72.401 20.711 72.584 20.751 ;
      RECT MASK 1 73.158 20.711 73.341 20.751 ;
      RECT MASK 1 73.563 20.711 73.746 20.751 ;
      RECT MASK 1 74.32 20.711 74.503 20.751 ;
      RECT MASK 1 74.725 20.711 74.908 20.751 ;
      RECT MASK 1 75.482 20.711 75.665 20.751 ;
      RECT MASK 1 75.887 20.711 76.07 20.751 ;
      RECT MASK 1 78.614 20.711 78.797 20.751 ;
      RECT MASK 1 79.019 20.711 79.202 20.751 ;
      RECT MASK 1 79.776 20.711 79.959 20.751 ;
      RECT MASK 1 80.181 20.711 80.364 20.751 ;
      RECT MASK 1 80.938 20.711 81.121 20.751 ;
      RECT MASK 1 81.343 20.711 81.526 20.751 ;
      RECT MASK 1 82.1 20.711 82.283 20.751 ;
      RECT MASK 1 82.505 20.711 82.688 20.751 ;
      RECT MASK 1 85.232 20.711 85.415 20.751 ;
      RECT MASK 1 85.637 20.711 85.82 20.751 ;
      RECT MASK 1 86.394 20.711 86.577 20.751 ;
      RECT MASK 1 86.799 20.711 86.982 20.751 ;
      RECT MASK 1 87.556 20.711 87.739 20.751 ;
      RECT MASK 1 87.961 20.711 88.144 20.751 ;
      RECT MASK 1 88.718 20.711 88.901 20.751 ;
      RECT MASK 1 89.123 20.711 89.306 20.751 ;
      RECT MASK 1 91.85 20.711 92.033 20.751 ;
      RECT MASK 1 92.255 20.711 92.438 20.751 ;
      RECT MASK 1 93.012 20.711 93.195 20.751 ;
      RECT MASK 1 93.417 20.711 93.6 20.751 ;
      RECT MASK 1 94.174 20.711 94.357 20.751 ;
      RECT MASK 1 94.579 20.711 94.762 20.751 ;
      RECT MASK 1 95.336 20.711 95.519 20.751 ;
      RECT MASK 1 95.741 20.711 95.924 20.751 ;
      RECT MASK 1 98.468 20.711 98.651 20.751 ;
      RECT MASK 1 98.873 20.711 99.056 20.751 ;
      RECT MASK 1 99.63 20.711 99.813 20.751 ;
      RECT MASK 1 100.035 20.711 100.218 20.751 ;
      RECT MASK 1 100.792 20.711 100.975 20.751 ;
      RECT MASK 1 101.197 20.711 101.38 20.751 ;
      RECT MASK 1 101.954 20.711 102.137 20.751 ;
      RECT MASK 1 102.359 20.711 102.542 20.751 ;
      RECT MASK 1 105.086 20.711 105.269 20.751 ;
      RECT MASK 1 105.491 20.711 105.674 20.751 ;
      RECT MASK 1 106.248 20.711 106.431 20.751 ;
      RECT MASK 1 106.653 20.711 106.836 20.751 ;
      RECT MASK 1 107.41 20.711 107.593 20.751 ;
      RECT MASK 1 107.815 20.711 107.998 20.751 ;
      RECT MASK 1 108.572 20.711 108.755 20.751 ;
      RECT MASK 1 108.977 20.711 109.16 20.751 ;
      RECT MASK 1 5.107 20.895 109.869 20.935 ;
      RECT MASK 1 5.1135 21.079 109.836 21.119 ;
      RECT MASK 1 5.1135 21.445 109.836 21.485 ;
      RECT MASK 1 2.225 21.48 2.285 22.53 ;
      RECT MASK 1 2.499 21.48 2.559 22.53 ;
      RECT MASK 1 2.773 21.48 2.833 22.53 ;
      RECT MASK 1 3.047 21.48 3.107 22.53 ;
      RECT MASK 1 3.321 21.48 3.381 22.53 ;
      RECT MASK 1 3.595 21.48 3.655 22.53 ;
      RECT MASK 1 3.869 21.48 3.929 22.53 ;
      RECT MASK 1 5.157 21.742 5.237 23.16 ;
      RECT MASK 1 10.469 21.742 10.549 23.16 ;
      RECT MASK 1 11.775 21.742 11.855 23.16 ;
      RECT MASK 1 17.087 21.742 17.167 23.16 ;
      RECT MASK 1 18.393 21.742 18.473 23.16 ;
      RECT MASK 1 23.705 21.742 23.785 23.16 ;
      RECT MASK 1 25.011 21.742 25.091 23.16 ;
      RECT MASK 1 30.323 21.742 30.403 23.16 ;
      RECT MASK 1 31.629 21.742 31.709 23.16 ;
      RECT MASK 1 36.941 21.742 37.021 23.16 ;
      RECT MASK 1 38.247 21.742 38.327 23.16 ;
      RECT MASK 1 43.559 21.742 43.639 23.16 ;
      RECT MASK 1 44.865 21.742 44.945 23.16 ;
      RECT MASK 1 50.177 21.742 50.257 23.16 ;
      RECT MASK 1 51.483 21.742 51.563 23.16 ;
      RECT MASK 1 56.795 21.742 56.875 23.16 ;
      RECT MASK 1 58.101 21.742 58.181 23.16 ;
      RECT MASK 1 63.413 21.742 63.493 23.16 ;
      RECT MASK 1 64.719 21.742 64.799 23.16 ;
      RECT MASK 1 70.031 21.742 70.111 23.16 ;
      RECT MASK 1 71.337 21.742 71.417 23.16 ;
      RECT MASK 1 76.649 21.742 76.729 23.16 ;
      RECT MASK 1 77.955 21.742 78.035 23.16 ;
      RECT MASK 1 83.267 21.742 83.347 23.16 ;
      RECT MASK 1 84.573 21.742 84.653 23.16 ;
      RECT MASK 1 89.885 21.742 89.965 23.16 ;
      RECT MASK 1 91.191 21.742 91.271 23.16 ;
      RECT MASK 1 96.503 21.742 96.583 23.16 ;
      RECT MASK 1 97.809 21.742 97.889 23.16 ;
      RECT MASK 1 103.121 21.742 103.201 23.16 ;
      RECT MASK 1 104.427 21.742 104.507 23.16 ;
      RECT MASK 1 109.739 21.742 109.819 23.16 ;
      RECT MASK 1 5.8885 21.874 6.165 21.914 ;
      RECT MASK 1 7.0505 21.874 7.327 21.914 ;
      RECT MASK 1 8.2125 21.874 8.489 21.914 ;
      RECT MASK 1 9.3745 21.874 9.651 21.914 ;
      RECT MASK 1 12.5065 21.874 12.783 21.914 ;
      RECT MASK 1 13.6685 21.874 13.945 21.914 ;
      RECT MASK 1 14.8305 21.874 15.107 21.914 ;
      RECT MASK 1 15.9925 21.874 16.269 21.914 ;
      RECT MASK 1 19.1245 21.874 19.401 21.914 ;
      RECT MASK 1 20.2865 21.874 20.563 21.914 ;
      RECT MASK 1 21.4485 21.874 21.725 21.914 ;
      RECT MASK 1 22.6105 21.874 22.887 21.914 ;
      RECT MASK 1 25.7425 21.874 26.019 21.914 ;
      RECT MASK 1 26.9045 21.874 27.181 21.914 ;
      RECT MASK 1 28.0665 21.874 28.343 21.914 ;
      RECT MASK 1 29.2285 21.874 29.505 21.914 ;
      RECT MASK 1 32.3605 21.874 32.637 21.914 ;
      RECT MASK 1 33.5225 21.874 33.799 21.914 ;
      RECT MASK 1 34.6845 21.874 34.961 21.914 ;
      RECT MASK 1 35.8465 21.874 36.123 21.914 ;
      RECT MASK 1 38.9785 21.874 39.255 21.914 ;
      RECT MASK 1 40.1405 21.874 40.417 21.914 ;
      RECT MASK 1 41.3025 21.874 41.579 21.914 ;
      RECT MASK 1 42.4645 21.874 42.741 21.914 ;
      RECT MASK 1 45.5965 21.874 45.873 21.914 ;
      RECT MASK 1 46.7585 21.874 47.035 21.914 ;
      RECT MASK 1 47.9205 21.874 48.197 21.914 ;
      RECT MASK 1 49.0825 21.874 49.359 21.914 ;
      RECT MASK 1 52.2145 21.874 52.491 21.914 ;
      RECT MASK 1 53.3765 21.874 53.653 21.914 ;
      RECT MASK 1 54.5385 21.874 54.815 21.914 ;
      RECT MASK 1 55.7005 21.874 55.977 21.914 ;
      RECT MASK 1 58.8325 21.874 59.109 21.914 ;
      RECT MASK 1 59.9945 21.874 60.271 21.914 ;
      RECT MASK 1 61.1565 21.874 61.433 21.914 ;
      RECT MASK 1 62.3185 21.874 62.595 21.914 ;
      RECT MASK 1 65.4505 21.874 65.727 21.914 ;
      RECT MASK 1 66.6125 21.874 66.889 21.914 ;
      RECT MASK 1 67.7745 21.874 68.051 21.914 ;
      RECT MASK 1 68.9365 21.874 69.213 21.914 ;
      RECT MASK 1 72.0685 21.874 72.345 21.914 ;
      RECT MASK 1 73.2305 21.874 73.507 21.914 ;
      RECT MASK 1 74.3925 21.874 74.669 21.914 ;
      RECT MASK 1 75.5545 21.874 75.831 21.914 ;
      RECT MASK 1 78.6865 21.874 78.963 21.914 ;
      RECT MASK 1 79.8485 21.874 80.125 21.914 ;
      RECT MASK 1 81.0105 21.874 81.287 21.914 ;
      RECT MASK 1 82.1725 21.874 82.449 21.914 ;
      RECT MASK 1 85.3045 21.874 85.581 21.914 ;
      RECT MASK 1 86.4665 21.874 86.743 21.914 ;
      RECT MASK 1 87.6285 21.874 87.905 21.914 ;
      RECT MASK 1 88.7905 21.874 89.067 21.914 ;
      RECT MASK 1 91.9225 21.874 92.199 21.914 ;
      RECT MASK 1 93.0845 21.874 93.361 21.914 ;
      RECT MASK 1 94.2465 21.874 94.523 21.914 ;
      RECT MASK 1 95.4085 21.874 95.685 21.914 ;
      RECT MASK 1 98.5405 21.874 98.817 21.914 ;
      RECT MASK 1 99.7025 21.874 99.979 21.914 ;
      RECT MASK 1 100.8645 21.874 101.141 21.914 ;
      RECT MASK 1 102.0265 21.874 102.303 21.914 ;
      RECT MASK 1 105.1585 21.874 105.435 21.914 ;
      RECT MASK 1 106.3205 21.874 106.597 21.914 ;
      RECT MASK 1 107.4825 21.874 107.759 21.914 ;
      RECT MASK 1 108.6445 21.874 108.921 21.914 ;
      RECT MASK 1 5.821 22.098 5.901 22.3285 ;
      RECT MASK 1 6.153 22.098 6.233 22.3285 ;
      RECT MASK 1 6.983 22.098 7.063 22.3285 ;
      RECT MASK 1 7.315 22.098 7.395 22.3285 ;
      RECT MASK 1 8.145 22.098 8.225 22.3285 ;
      RECT MASK 1 8.477 22.098 8.557 22.3285 ;
      RECT MASK 1 9.307 22.098 9.387 22.3285 ;
      RECT MASK 1 9.639 22.098 9.719 22.3285 ;
      RECT MASK 1 12.439 22.098 12.519 22.3285 ;
      RECT MASK 1 12.771 22.098 12.851 22.3285 ;
      RECT MASK 1 13.601 22.098 13.681 22.3285 ;
      RECT MASK 1 13.933 22.098 14.013 22.3285 ;
      RECT MASK 1 14.763 22.098 14.843 22.3285 ;
      RECT MASK 1 15.095 22.098 15.175 22.3285 ;
      RECT MASK 1 15.925 22.098 16.005 22.3285 ;
      RECT MASK 1 16.257 22.098 16.337 22.3285 ;
      RECT MASK 1 19.057 22.098 19.137 22.3285 ;
      RECT MASK 1 19.389 22.098 19.469 22.3285 ;
      RECT MASK 1 20.219 22.098 20.299 22.3285 ;
      RECT MASK 1 20.551 22.098 20.631 22.3285 ;
      RECT MASK 1 21.381 22.098 21.461 22.3285 ;
      RECT MASK 1 21.713 22.098 21.793 22.3285 ;
      RECT MASK 1 22.543 22.098 22.623 22.3285 ;
      RECT MASK 1 22.875 22.098 22.955 22.3285 ;
      RECT MASK 1 25.675 22.098 25.755 22.3285 ;
      RECT MASK 1 26.007 22.098 26.087 22.3285 ;
      RECT MASK 1 26.837 22.098 26.917 22.3285 ;
      RECT MASK 1 27.169 22.098 27.249 22.3285 ;
      RECT MASK 1 27.999 22.098 28.079 22.3285 ;
      RECT MASK 1 28.331 22.098 28.411 22.3285 ;
      RECT MASK 1 29.161 22.098 29.241 22.3285 ;
      RECT MASK 1 29.493 22.098 29.573 22.3285 ;
      RECT MASK 1 32.293 22.098 32.373 22.3285 ;
      RECT MASK 1 32.625 22.098 32.705 22.3285 ;
      RECT MASK 1 33.455 22.098 33.535 22.3285 ;
      RECT MASK 1 33.787 22.098 33.867 22.3285 ;
      RECT MASK 1 34.617 22.098 34.697 22.3285 ;
      RECT MASK 1 34.949 22.098 35.029 22.3285 ;
      RECT MASK 1 35.779 22.098 35.859 22.3285 ;
      RECT MASK 1 36.111 22.098 36.191 22.3285 ;
      RECT MASK 1 38.911 22.098 38.991 22.3285 ;
      RECT MASK 1 39.243 22.098 39.323 22.3285 ;
      RECT MASK 1 40.073 22.098 40.153 22.3285 ;
      RECT MASK 1 40.405 22.098 40.485 22.3285 ;
      RECT MASK 1 41.235 22.098 41.315 22.3285 ;
      RECT MASK 1 41.567 22.098 41.647 22.3285 ;
      RECT MASK 1 42.397 22.098 42.477 22.3285 ;
      RECT MASK 1 42.729 22.098 42.809 22.3285 ;
      RECT MASK 1 45.529 22.098 45.609 22.3285 ;
      RECT MASK 1 45.861 22.098 45.941 22.3285 ;
      RECT MASK 1 46.691 22.098 46.771 22.3285 ;
      RECT MASK 1 47.023 22.098 47.103 22.3285 ;
      RECT MASK 1 47.853 22.098 47.933 22.3285 ;
      RECT MASK 1 48.185 22.098 48.265 22.3285 ;
      RECT MASK 1 49.015 22.098 49.095 22.3285 ;
      RECT MASK 1 49.347 22.098 49.427 22.3285 ;
      RECT MASK 1 52.147 22.098 52.227 22.3285 ;
      RECT MASK 1 52.479 22.098 52.559 22.3285 ;
      RECT MASK 1 53.309 22.098 53.389 22.3285 ;
      RECT MASK 1 53.641 22.098 53.721 22.3285 ;
      RECT MASK 1 54.471 22.098 54.551 22.3285 ;
      RECT MASK 1 54.803 22.098 54.883 22.3285 ;
      RECT MASK 1 55.633 22.098 55.713 22.3285 ;
      RECT MASK 1 55.965 22.098 56.045 22.3285 ;
      RECT MASK 1 58.765 22.098 58.845 22.3285 ;
      RECT MASK 1 59.097 22.098 59.177 22.3285 ;
      RECT MASK 1 59.927 22.098 60.007 22.3285 ;
      RECT MASK 1 60.259 22.098 60.339 22.3285 ;
      RECT MASK 1 61.089 22.098 61.169 22.3285 ;
      RECT MASK 1 61.421 22.098 61.501 22.3285 ;
      RECT MASK 1 62.251 22.098 62.331 22.3285 ;
      RECT MASK 1 62.583 22.098 62.663 22.3285 ;
      RECT MASK 1 65.383 22.098 65.463 22.3285 ;
      RECT MASK 1 65.715 22.098 65.795 22.3285 ;
      RECT MASK 1 66.545 22.098 66.625 22.3285 ;
      RECT MASK 1 66.877 22.098 66.957 22.3285 ;
      RECT MASK 1 67.707 22.098 67.787 22.3285 ;
      RECT MASK 1 68.039 22.098 68.119 22.3285 ;
      RECT MASK 1 68.869 22.098 68.949 22.3285 ;
      RECT MASK 1 69.201 22.098 69.281 22.3285 ;
      RECT MASK 1 72.001 22.098 72.081 22.3285 ;
      RECT MASK 1 72.333 22.098 72.413 22.3285 ;
      RECT MASK 1 73.163 22.098 73.243 22.3285 ;
      RECT MASK 1 73.495 22.098 73.575 22.3285 ;
      RECT MASK 1 74.325 22.098 74.405 22.3285 ;
      RECT MASK 1 74.657 22.098 74.737 22.3285 ;
      RECT MASK 1 75.487 22.098 75.567 22.3285 ;
      RECT MASK 1 75.819 22.098 75.899 22.3285 ;
      RECT MASK 1 78.619 22.098 78.699 22.3285 ;
      RECT MASK 1 78.951 22.098 79.031 22.3285 ;
      RECT MASK 1 79.781 22.098 79.861 22.3285 ;
      RECT MASK 1 80.113 22.098 80.193 22.3285 ;
      RECT MASK 1 80.943 22.098 81.023 22.3285 ;
      RECT MASK 1 81.275 22.098 81.355 22.3285 ;
      RECT MASK 1 82.105 22.098 82.185 22.3285 ;
      RECT MASK 1 82.437 22.098 82.517 22.3285 ;
      RECT MASK 1 85.237 22.098 85.317 22.3285 ;
      RECT MASK 1 85.569 22.098 85.649 22.3285 ;
      RECT MASK 1 86.399 22.098 86.479 22.3285 ;
      RECT MASK 1 86.731 22.098 86.811 22.3285 ;
      RECT MASK 1 87.561 22.098 87.641 22.3285 ;
      RECT MASK 1 87.893 22.098 87.973 22.3285 ;
      RECT MASK 1 88.723 22.098 88.803 22.3285 ;
      RECT MASK 1 89.055 22.098 89.135 22.3285 ;
      RECT MASK 1 91.855 22.098 91.935 22.3285 ;
      RECT MASK 1 92.187 22.098 92.267 22.3285 ;
      RECT MASK 1 93.017 22.098 93.097 22.3285 ;
      RECT MASK 1 93.349 22.098 93.429 22.3285 ;
      RECT MASK 1 94.179 22.098 94.259 22.3285 ;
      RECT MASK 1 94.511 22.098 94.591 22.3285 ;
      RECT MASK 1 95.341 22.098 95.421 22.3285 ;
      RECT MASK 1 95.673 22.098 95.753 22.3285 ;
      RECT MASK 1 98.473 22.098 98.553 22.3285 ;
      RECT MASK 1 98.805 22.098 98.885 22.3285 ;
      RECT MASK 1 99.635 22.098 99.715 22.3285 ;
      RECT MASK 1 99.967 22.098 100.047 22.3285 ;
      RECT MASK 1 100.797 22.098 100.877 22.3285 ;
      RECT MASK 1 101.129 22.098 101.209 22.3285 ;
      RECT MASK 1 101.959 22.098 102.039 22.3285 ;
      RECT MASK 1 102.291 22.098 102.371 22.3285 ;
      RECT MASK 1 105.091 22.098 105.171 22.3285 ;
      RECT MASK 1 105.423 22.098 105.503 22.3285 ;
      RECT MASK 1 106.253 22.098 106.333 22.3285 ;
      RECT MASK 1 106.585 22.098 106.665 22.3285 ;
      RECT MASK 1 107.415 22.098 107.495 22.3285 ;
      RECT MASK 1 107.747 22.098 107.827 22.3285 ;
      RECT MASK 1 108.577 22.098 108.657 22.3285 ;
      RECT MASK 1 108.909 22.098 108.989 22.3285 ;
      RECT MASK 1 116.154 22.41 116.214 23.46 ;
      RECT MASK 1 116.428 22.41 116.488 23.46 ;
      RECT MASK 1 116.702 22.41 116.762 23.46 ;
      RECT MASK 1 116.976 22.41 117.036 23.46 ;
      RECT MASK 1 117.25 22.41 117.31 23.46 ;
      RECT MASK 1 117.524 22.41 117.584 23.46 ;
      RECT MASK 1 117.798 22.41 117.858 23.46 ;
      RECT MASK 1 118.072 22.41 118.132 23.46 ;
      RECT MASK 1 118.346 22.41 118.406 23.46 ;
      RECT MASK 1 118.62 22.41 118.68 23.46 ;
      RECT MASK 1 118.894 22.41 118.954 23.46 ;
      RECT MASK 1 119.168 22.41 119.228 23.46 ;
      RECT MASK 1 119.442 22.41 119.502 23.46 ;
      RECT MASK 1 119.716 22.41 119.776 23.46 ;
      RECT MASK 1 119.99 22.41 120.05 23.46 ;
      RECT MASK 1 120.264 22.41 120.324 23.46 ;
      RECT MASK 1 120.538 22.41 120.598 23.46 ;
      RECT MASK 1 120.812 22.41 120.872 23.46 ;
      RECT MASK 1 121.086 22.41 121.146 23.46 ;
      RECT MASK 1 121.36 22.41 121.42 23.46 ;
      RECT MASK 1 121.634 22.41 121.694 23.46 ;
      RECT MASK 1 121.908 22.41 121.968 23.46 ;
      RECT MASK 1 122.182 22.41 122.242 23.46 ;
      RECT MASK 1 122.456 22.41 122.516 23.46 ;
      RECT MASK 1 122.73 22.41 122.79 23.46 ;
      RECT MASK 1 123.004 22.41 123.064 23.46 ;
      RECT MASK 1 123.278 22.41 123.338 23.46 ;
      RECT MASK 1 123.552 22.41 123.612 23.46 ;
      RECT MASK 1 123.826 22.41 123.886 23.46 ;
      RECT MASK 1 124.1 22.41 124.16 23.46 ;
      RECT MASK 1 124.374 22.41 124.434 23.46 ;
      RECT MASK 1 124.648 22.41 124.708 23.46 ;
      RECT MASK 1 124.922 22.41 124.982 23.46 ;
      RECT MASK 1 125.196 22.41 125.256 23.46 ;
      RECT MASK 1 125.47 22.41 125.53 23.46 ;
      RECT MASK 1 125.744 22.41 125.804 23.46 ;
      RECT MASK 1 126.018 22.41 126.078 23.46 ;
      RECT MASK 1 126.292 22.41 126.352 23.46 ;
      RECT MASK 1 126.566 22.41 126.626 23.46 ;
      RECT MASK 1 126.84 22.41 126.9 23.46 ;
      RECT MASK 1 127.114 22.41 127.174 23.46 ;
      RECT MASK 1 127.388 22.41 127.448 23.46 ;
      RECT MASK 1 127.662 22.41 127.722 23.46 ;
      RECT MASK 1 127.936 22.41 127.996 23.46 ;
      RECT MASK 1 128.21 22.41 128.27 23.46 ;
      RECT MASK 1 5.529 22.54 10.315 22.58 ;
      RECT MASK 1 12.009 22.54 16.933 22.58 ;
      RECT MASK 1 18.627 22.54 23.551 22.58 ;
      RECT MASK 1 25.245 22.54 30.169 22.58 ;
      RECT MASK 1 31.863 22.54 36.787 22.58 ;
      RECT MASK 1 38.481 22.54 43.405 22.58 ;
      RECT MASK 1 45.099 22.54 50.023 22.58 ;
      RECT MASK 1 51.717 22.54 56.641 22.58 ;
      RECT MASK 1 58.335 22.54 63.259 22.58 ;
      RECT MASK 1 64.953 22.54 69.877 22.58 ;
      RECT MASK 1 71.571 22.54 76.495 22.58 ;
      RECT MASK 1 78.189 22.54 83.113 22.58 ;
      RECT MASK 1 84.807 22.54 89.731 22.58 ;
      RECT MASK 1 91.425 22.54 96.349 22.58 ;
      RECT MASK 1 98.043 22.54 102.967 22.58 ;
      RECT MASK 1 104.661 22.54 109.585 22.58 ;
      RECT MASK 1 5.821 22.769 5.901 22.994 ;
      RECT MASK 1 6.153 22.769 6.233 22.994 ;
      RECT MASK 1 6.983 22.769 7.063 22.994 ;
      RECT MASK 1 7.315 22.769 7.395 22.994 ;
      RECT MASK 1 8.145 22.769 8.225 22.994 ;
      RECT MASK 1 8.477 22.769 8.557 22.994 ;
      RECT MASK 1 9.307 22.769 9.387 22.994 ;
      RECT MASK 1 9.639 22.769 9.719 22.994 ;
      RECT MASK 1 12.439 22.769 12.519 22.994 ;
      RECT MASK 1 12.771 22.769 12.851 22.994 ;
      RECT MASK 1 13.601 22.769 13.681 22.994 ;
      RECT MASK 1 13.933 22.769 14.013 22.994 ;
      RECT MASK 1 14.763 22.769 14.843 22.994 ;
      RECT MASK 1 15.095 22.769 15.175 22.994 ;
      RECT MASK 1 15.925 22.769 16.005 22.994 ;
      RECT MASK 1 16.257 22.769 16.337 22.994 ;
      RECT MASK 1 19.057 22.769 19.137 22.994 ;
      RECT MASK 1 19.389 22.769 19.469 22.994 ;
      RECT MASK 1 20.219 22.769 20.299 22.994 ;
      RECT MASK 1 20.551 22.769 20.631 22.994 ;
      RECT MASK 1 21.381 22.769 21.461 22.994 ;
      RECT MASK 1 21.713 22.769 21.793 22.994 ;
      RECT MASK 1 22.543 22.769 22.623 22.994 ;
      RECT MASK 1 22.875 22.769 22.955 22.994 ;
      RECT MASK 1 25.675 22.769 25.755 22.994 ;
      RECT MASK 1 26.007 22.769 26.087 22.994 ;
      RECT MASK 1 26.837 22.769 26.917 22.994 ;
      RECT MASK 1 27.169 22.769 27.249 22.994 ;
      RECT MASK 1 27.999 22.769 28.079 22.994 ;
      RECT MASK 1 28.331 22.769 28.411 22.994 ;
      RECT MASK 1 29.161 22.769 29.241 22.994 ;
      RECT MASK 1 29.493 22.769 29.573 22.994 ;
      RECT MASK 1 32.293 22.769 32.373 22.994 ;
      RECT MASK 1 32.625 22.769 32.705 22.994 ;
      RECT MASK 1 33.455 22.769 33.535 22.994 ;
      RECT MASK 1 33.787 22.769 33.867 22.994 ;
      RECT MASK 1 34.617 22.769 34.697 22.994 ;
      RECT MASK 1 34.949 22.769 35.029 22.994 ;
      RECT MASK 1 35.779 22.769 35.859 22.994 ;
      RECT MASK 1 36.111 22.769 36.191 22.994 ;
      RECT MASK 1 38.911 22.769 38.991 22.994 ;
      RECT MASK 1 39.243 22.769 39.323 22.994 ;
      RECT MASK 1 40.073 22.769 40.153 22.994 ;
      RECT MASK 1 40.405 22.769 40.485 22.994 ;
      RECT MASK 1 41.235 22.769 41.315 22.994 ;
      RECT MASK 1 41.567 22.769 41.647 22.994 ;
      RECT MASK 1 42.397 22.769 42.477 22.994 ;
      RECT MASK 1 42.729 22.769 42.809 22.994 ;
      RECT MASK 1 45.529 22.769 45.609 22.994 ;
      RECT MASK 1 45.861 22.769 45.941 22.994 ;
      RECT MASK 1 46.691 22.769 46.771 22.994 ;
      RECT MASK 1 47.023 22.769 47.103 22.994 ;
      RECT MASK 1 47.853 22.769 47.933 22.994 ;
      RECT MASK 1 48.185 22.769 48.265 22.994 ;
      RECT MASK 1 49.015 22.769 49.095 22.994 ;
      RECT MASK 1 49.347 22.769 49.427 22.994 ;
      RECT MASK 1 52.147 22.769 52.227 22.994 ;
      RECT MASK 1 52.479 22.769 52.559 22.994 ;
      RECT MASK 1 53.309 22.769 53.389 22.994 ;
      RECT MASK 1 53.641 22.769 53.721 22.994 ;
      RECT MASK 1 54.471 22.769 54.551 22.994 ;
      RECT MASK 1 54.803 22.769 54.883 22.994 ;
      RECT MASK 1 55.633 22.769 55.713 22.994 ;
      RECT MASK 1 55.965 22.769 56.045 22.994 ;
      RECT MASK 1 58.765 22.769 58.845 22.994 ;
      RECT MASK 1 59.097 22.769 59.177 22.994 ;
      RECT MASK 1 59.927 22.769 60.007 22.994 ;
      RECT MASK 1 60.259 22.769 60.339 22.994 ;
      RECT MASK 1 61.089 22.769 61.169 22.994 ;
      RECT MASK 1 61.421 22.769 61.501 22.994 ;
      RECT MASK 1 62.251 22.769 62.331 22.994 ;
      RECT MASK 1 62.583 22.769 62.663 22.994 ;
      RECT MASK 1 65.383 22.769 65.463 22.994 ;
      RECT MASK 1 65.715 22.769 65.795 22.994 ;
      RECT MASK 1 66.545 22.769 66.625 22.994 ;
      RECT MASK 1 66.877 22.769 66.957 22.994 ;
      RECT MASK 1 67.707 22.769 67.787 22.994 ;
      RECT MASK 1 68.039 22.769 68.119 22.994 ;
      RECT MASK 1 68.869 22.769 68.949 22.994 ;
      RECT MASK 1 69.201 22.769 69.281 22.994 ;
      RECT MASK 1 72.001 22.769 72.081 22.994 ;
      RECT MASK 1 72.333 22.769 72.413 22.994 ;
      RECT MASK 1 73.163 22.769 73.243 22.994 ;
      RECT MASK 1 73.495 22.769 73.575 22.994 ;
      RECT MASK 1 74.325 22.769 74.405 22.994 ;
      RECT MASK 1 74.657 22.769 74.737 22.994 ;
      RECT MASK 1 75.487 22.769 75.567 22.994 ;
      RECT MASK 1 75.819 22.769 75.899 22.994 ;
      RECT MASK 1 78.619 22.769 78.699 22.994 ;
      RECT MASK 1 78.951 22.769 79.031 22.994 ;
      RECT MASK 1 79.781 22.769 79.861 22.994 ;
      RECT MASK 1 80.113 22.769 80.193 22.994 ;
      RECT MASK 1 80.943 22.769 81.023 22.994 ;
      RECT MASK 1 81.275 22.769 81.355 22.994 ;
      RECT MASK 1 82.105 22.769 82.185 22.994 ;
      RECT MASK 1 82.437 22.769 82.517 22.994 ;
      RECT MASK 1 85.237 22.769 85.317 22.994 ;
      RECT MASK 1 85.569 22.769 85.649 22.994 ;
      RECT MASK 1 86.399 22.769 86.479 22.994 ;
      RECT MASK 1 86.731 22.769 86.811 22.994 ;
      RECT MASK 1 87.561 22.769 87.641 22.994 ;
      RECT MASK 1 87.893 22.769 87.973 22.994 ;
      RECT MASK 1 88.723 22.769 88.803 22.994 ;
      RECT MASK 1 89.055 22.769 89.135 22.994 ;
      RECT MASK 1 91.855 22.769 91.935 22.994 ;
      RECT MASK 1 92.187 22.769 92.267 22.994 ;
      RECT MASK 1 93.017 22.769 93.097 22.994 ;
      RECT MASK 1 93.349 22.769 93.429 22.994 ;
      RECT MASK 1 94.179 22.769 94.259 22.994 ;
      RECT MASK 1 94.511 22.769 94.591 22.994 ;
      RECT MASK 1 95.341 22.769 95.421 22.994 ;
      RECT MASK 1 95.673 22.769 95.753 22.994 ;
      RECT MASK 1 98.473 22.769 98.553 22.994 ;
      RECT MASK 1 98.805 22.769 98.885 22.994 ;
      RECT MASK 1 99.635 22.769 99.715 22.994 ;
      RECT MASK 1 99.967 22.769 100.047 22.994 ;
      RECT MASK 1 100.797 22.769 100.877 22.994 ;
      RECT MASK 1 101.129 22.769 101.209 22.994 ;
      RECT MASK 1 101.959 22.769 102.039 22.994 ;
      RECT MASK 1 102.291 22.769 102.371 22.994 ;
      RECT MASK 1 105.091 22.769 105.171 22.994 ;
      RECT MASK 1 105.423 22.769 105.503 22.994 ;
      RECT MASK 1 106.253 22.769 106.333 22.994 ;
      RECT MASK 1 106.585 22.769 106.665 22.994 ;
      RECT MASK 1 107.415 22.769 107.495 22.994 ;
      RECT MASK 1 107.747 22.769 107.827 22.994 ;
      RECT MASK 1 108.577 22.769 108.657 22.994 ;
      RECT MASK 1 108.909 22.769 108.989 22.994 ;
      RECT MASK 1 2.225 23.19 2.285 24.24 ;
      RECT MASK 1 2.499 23.19 2.559 24.24 ;
      RECT MASK 1 2.773 23.19 2.833 24.24 ;
      RECT MASK 1 3.047 23.19 3.107 24.24 ;
      RECT MASK 1 3.321 23.19 3.381 24.24 ;
      RECT MASK 1 3.595 23.19 3.655 24.24 ;
      RECT MASK 1 3.869 23.19 3.929 24.24 ;
      RECT MASK 1 5.1135 23.395 109.836 23.435 ;
      RECT MASK 1 5.1135 23.845 110.065 23.885 ;
      RECT MASK 1 115.425 23.845 129.001 23.885 ;
      RECT MASK 1 5.157 24.142 5.237 25.56 ;
      RECT MASK 1 10.469 24.142 10.549 25.56 ;
      RECT MASK 1 11.775 24.142 11.855 25.56 ;
      RECT MASK 1 17.087 24.142 17.167 25.56 ;
      RECT MASK 1 18.393 24.142 18.473 25.56 ;
      RECT MASK 1 23.705 24.142 23.785 25.56 ;
      RECT MASK 1 25.011 24.142 25.091 25.56 ;
      RECT MASK 1 30.323 24.142 30.403 25.56 ;
      RECT MASK 1 31.629 24.142 31.709 25.56 ;
      RECT MASK 1 36.941 24.142 37.021 25.56 ;
      RECT MASK 1 38.247 24.142 38.327 25.56 ;
      RECT MASK 1 43.559 24.142 43.639 25.56 ;
      RECT MASK 1 44.865 24.142 44.945 25.56 ;
      RECT MASK 1 50.177 24.142 50.257 25.56 ;
      RECT MASK 1 51.483 24.142 51.563 25.56 ;
      RECT MASK 1 56.795 24.142 56.875 25.56 ;
      RECT MASK 1 58.101 24.142 58.181 25.56 ;
      RECT MASK 1 63.413 24.142 63.493 25.56 ;
      RECT MASK 1 64.719 24.142 64.799 25.56 ;
      RECT MASK 1 70.031 24.142 70.111 25.56 ;
      RECT MASK 1 71.337 24.142 71.417 25.56 ;
      RECT MASK 1 76.649 24.142 76.729 25.56 ;
      RECT MASK 1 77.955 24.142 78.035 25.56 ;
      RECT MASK 1 83.267 24.142 83.347 25.56 ;
      RECT MASK 1 84.573 24.142 84.653 25.56 ;
      RECT MASK 1 89.885 24.142 89.965 25.56 ;
      RECT MASK 1 91.191 24.142 91.271 25.56 ;
      RECT MASK 1 96.503 24.142 96.583 25.56 ;
      RECT MASK 1 97.809 24.142 97.889 25.56 ;
      RECT MASK 1 103.121 24.142 103.201 25.56 ;
      RECT MASK 1 104.427 24.142 104.507 25.56 ;
      RECT MASK 1 109.739 24.142 109.819 25.56 ;
      RECT MASK 1 5.529 24.264 10.315 24.304 ;
      RECT MASK 1 12.009 24.264 16.933 24.304 ;
      RECT MASK 1 18.627 24.264 23.551 24.304 ;
      RECT MASK 1 25.245 24.264 30.169 24.304 ;
      RECT MASK 1 31.863 24.264 36.787 24.304 ;
      RECT MASK 1 38.481 24.264 43.405 24.304 ;
      RECT MASK 1 45.099 24.264 50.023 24.304 ;
      RECT MASK 1 51.717 24.264 56.641 24.304 ;
      RECT MASK 1 58.335 24.264 63.259 24.304 ;
      RECT MASK 1 64.953 24.264 69.877 24.304 ;
      RECT MASK 1 71.571 24.264 76.495 24.304 ;
      RECT MASK 1 78.189 24.264 83.113 24.304 ;
      RECT MASK 1 84.807 24.264 89.731 24.304 ;
      RECT MASK 1 91.425 24.264 96.349 24.304 ;
      RECT MASK 1 98.043 24.264 102.967 24.304 ;
      RECT MASK 1 104.661 24.264 109.585 24.304 ;
      RECT MASK 1 5.821 24.502 5.901 24.7285 ;
      RECT MASK 1 6.153 24.502 6.233 24.7285 ;
      RECT MASK 1 6.983 24.502 7.063 24.7285 ;
      RECT MASK 1 7.315 24.502 7.395 24.7285 ;
      RECT MASK 1 8.145 24.502 8.225 24.7285 ;
      RECT MASK 1 8.477 24.502 8.557 24.7285 ;
      RECT MASK 1 9.307 24.502 9.387 24.7285 ;
      RECT MASK 1 9.639 24.502 9.719 24.7285 ;
      RECT MASK 1 12.439 24.502 12.519 24.7285 ;
      RECT MASK 1 12.771 24.502 12.851 24.7285 ;
      RECT MASK 1 13.601 24.502 13.681 24.7285 ;
      RECT MASK 1 13.933 24.502 14.013 24.7285 ;
      RECT MASK 1 14.763 24.502 14.843 24.7285 ;
      RECT MASK 1 15.095 24.502 15.175 24.7285 ;
      RECT MASK 1 15.925 24.502 16.005 24.7285 ;
      RECT MASK 1 16.257 24.502 16.337 24.7285 ;
      RECT MASK 1 19.057 24.502 19.137 24.7285 ;
      RECT MASK 1 19.389 24.502 19.469 24.7285 ;
      RECT MASK 1 20.219 24.502 20.299 24.7285 ;
      RECT MASK 1 20.551 24.502 20.631 24.7285 ;
      RECT MASK 1 21.381 24.502 21.461 24.7285 ;
      RECT MASK 1 21.713 24.502 21.793 24.7285 ;
      RECT MASK 1 22.543 24.502 22.623 24.7285 ;
      RECT MASK 1 22.875 24.502 22.955 24.7285 ;
      RECT MASK 1 25.675 24.502 25.755 24.7285 ;
      RECT MASK 1 26.007 24.502 26.087 24.7285 ;
      RECT MASK 1 26.837 24.502 26.917 24.7285 ;
      RECT MASK 1 27.169 24.502 27.249 24.7285 ;
      RECT MASK 1 27.999 24.502 28.079 24.7285 ;
      RECT MASK 1 28.331 24.502 28.411 24.7285 ;
      RECT MASK 1 29.161 24.502 29.241 24.7285 ;
      RECT MASK 1 29.493 24.502 29.573 24.7285 ;
      RECT MASK 1 32.293 24.502 32.373 24.7285 ;
      RECT MASK 1 32.625 24.502 32.705 24.7285 ;
      RECT MASK 1 33.455 24.502 33.535 24.7285 ;
      RECT MASK 1 33.787 24.502 33.867 24.7285 ;
      RECT MASK 1 34.617 24.502 34.697 24.7285 ;
      RECT MASK 1 34.949 24.502 35.029 24.7285 ;
      RECT MASK 1 35.779 24.502 35.859 24.7285 ;
      RECT MASK 1 36.111 24.502 36.191 24.7285 ;
      RECT MASK 1 38.911 24.502 38.991 24.7285 ;
      RECT MASK 1 39.243 24.502 39.323 24.7285 ;
      RECT MASK 1 40.073 24.502 40.153 24.7285 ;
      RECT MASK 1 40.405 24.502 40.485 24.7285 ;
      RECT MASK 1 41.235 24.502 41.315 24.7285 ;
      RECT MASK 1 41.567 24.502 41.647 24.7285 ;
      RECT MASK 1 42.397 24.502 42.477 24.7285 ;
      RECT MASK 1 42.729 24.502 42.809 24.7285 ;
      RECT MASK 1 45.529 24.502 45.609 24.7285 ;
      RECT MASK 1 45.861 24.502 45.941 24.7285 ;
      RECT MASK 1 46.691 24.502 46.771 24.7285 ;
      RECT MASK 1 47.023 24.502 47.103 24.7285 ;
      RECT MASK 1 47.853 24.502 47.933 24.7285 ;
      RECT MASK 1 48.185 24.502 48.265 24.7285 ;
      RECT MASK 1 49.015 24.502 49.095 24.7285 ;
      RECT MASK 1 49.347 24.502 49.427 24.7285 ;
      RECT MASK 1 52.147 24.502 52.227 24.7285 ;
      RECT MASK 1 52.479 24.502 52.559 24.7285 ;
      RECT MASK 1 53.309 24.502 53.389 24.7285 ;
      RECT MASK 1 53.641 24.502 53.721 24.7285 ;
      RECT MASK 1 54.471 24.502 54.551 24.7285 ;
      RECT MASK 1 54.803 24.502 54.883 24.7285 ;
      RECT MASK 1 55.633 24.502 55.713 24.7285 ;
      RECT MASK 1 55.965 24.502 56.045 24.7285 ;
      RECT MASK 1 58.765 24.502 58.845 24.7285 ;
      RECT MASK 1 59.097 24.502 59.177 24.7285 ;
      RECT MASK 1 59.927 24.502 60.007 24.7285 ;
      RECT MASK 1 60.259 24.502 60.339 24.7285 ;
      RECT MASK 1 61.089 24.502 61.169 24.7285 ;
      RECT MASK 1 61.421 24.502 61.501 24.7285 ;
      RECT MASK 1 62.251 24.502 62.331 24.7285 ;
      RECT MASK 1 62.583 24.502 62.663 24.7285 ;
      RECT MASK 1 65.383 24.502 65.463 24.7285 ;
      RECT MASK 1 65.715 24.502 65.795 24.7285 ;
      RECT MASK 1 66.545 24.502 66.625 24.7285 ;
      RECT MASK 1 66.877 24.502 66.957 24.7285 ;
      RECT MASK 1 67.707 24.502 67.787 24.7285 ;
      RECT MASK 1 68.039 24.502 68.119 24.7285 ;
      RECT MASK 1 68.869 24.502 68.949 24.7285 ;
      RECT MASK 1 69.201 24.502 69.281 24.7285 ;
      RECT MASK 1 72.001 24.502 72.081 24.7285 ;
      RECT MASK 1 72.333 24.502 72.413 24.7285 ;
      RECT MASK 1 73.163 24.502 73.243 24.7285 ;
      RECT MASK 1 73.495 24.502 73.575 24.7285 ;
      RECT MASK 1 74.325 24.502 74.405 24.7285 ;
      RECT MASK 1 74.657 24.502 74.737 24.7285 ;
      RECT MASK 1 75.487 24.502 75.567 24.7285 ;
      RECT MASK 1 75.819 24.502 75.899 24.7285 ;
      RECT MASK 1 78.619 24.502 78.699 24.7285 ;
      RECT MASK 1 78.951 24.502 79.031 24.7285 ;
      RECT MASK 1 79.781 24.502 79.861 24.7285 ;
      RECT MASK 1 80.113 24.502 80.193 24.7285 ;
      RECT MASK 1 80.943 24.502 81.023 24.7285 ;
      RECT MASK 1 81.275 24.502 81.355 24.7285 ;
      RECT MASK 1 82.105 24.502 82.185 24.7285 ;
      RECT MASK 1 82.437 24.502 82.517 24.7285 ;
      RECT MASK 1 85.237 24.502 85.317 24.7285 ;
      RECT MASK 1 85.569 24.502 85.649 24.7285 ;
      RECT MASK 1 86.399 24.502 86.479 24.7285 ;
      RECT MASK 1 86.731 24.502 86.811 24.7285 ;
      RECT MASK 1 87.561 24.502 87.641 24.7285 ;
      RECT MASK 1 87.893 24.502 87.973 24.7285 ;
      RECT MASK 1 88.723 24.502 88.803 24.7285 ;
      RECT MASK 1 89.055 24.502 89.135 24.7285 ;
      RECT MASK 1 91.855 24.502 91.935 24.7285 ;
      RECT MASK 1 92.187 24.502 92.267 24.7285 ;
      RECT MASK 1 93.017 24.502 93.097 24.7285 ;
      RECT MASK 1 93.349 24.502 93.429 24.7285 ;
      RECT MASK 1 94.179 24.502 94.259 24.7285 ;
      RECT MASK 1 94.511 24.502 94.591 24.7285 ;
      RECT MASK 1 95.341 24.502 95.421 24.7285 ;
      RECT MASK 1 95.673 24.502 95.753 24.7285 ;
      RECT MASK 1 98.473 24.502 98.553 24.7285 ;
      RECT MASK 1 98.805 24.502 98.885 24.7285 ;
      RECT MASK 1 99.635 24.502 99.715 24.7285 ;
      RECT MASK 1 99.967 24.502 100.047 24.7285 ;
      RECT MASK 1 100.797 24.502 100.877 24.7285 ;
      RECT MASK 1 101.129 24.502 101.209 24.7285 ;
      RECT MASK 1 101.959 24.502 102.039 24.7285 ;
      RECT MASK 1 102.291 24.502 102.371 24.7285 ;
      RECT MASK 1 105.091 24.502 105.171 24.7285 ;
      RECT MASK 1 105.423 24.502 105.503 24.7285 ;
      RECT MASK 1 106.253 24.502 106.333 24.7285 ;
      RECT MASK 1 106.585 24.502 106.665 24.7285 ;
      RECT MASK 1 107.415 24.502 107.495 24.7285 ;
      RECT MASK 1 107.747 24.502 107.827 24.7285 ;
      RECT MASK 1 108.577 24.502 108.657 24.7285 ;
      RECT MASK 1 108.909 24.502 108.989 24.7285 ;
      RECT MASK 1 1.406 24.775 4.69 24.815 ;
      RECT MASK 1 5.899 24.939 6.58 24.979 ;
      RECT MASK 1 7.061 24.939 7.742 24.979 ;
      RECT MASK 1 8.223 24.939 8.904 24.979 ;
      RECT MASK 1 9.385 24.939 10.066 24.979 ;
      RECT MASK 1 12.517 24.939 13.198 24.979 ;
      RECT MASK 1 13.679 24.939 14.36 24.979 ;
      RECT MASK 1 14.841 24.939 15.522 24.979 ;
      RECT MASK 1 16.003 24.939 16.684 24.979 ;
      RECT MASK 1 19.135 24.939 19.816 24.979 ;
      RECT MASK 1 20.297 24.939 20.978 24.979 ;
      RECT MASK 1 21.459 24.939 22.14 24.979 ;
      RECT MASK 1 22.621 24.939 23.302 24.979 ;
      RECT MASK 1 25.753 24.939 26.434 24.979 ;
      RECT MASK 1 26.915 24.939 27.596 24.979 ;
      RECT MASK 1 28.077 24.939 28.758 24.979 ;
      RECT MASK 1 29.239 24.939 29.92 24.979 ;
      RECT MASK 1 32.371 24.939 33.052 24.979 ;
      RECT MASK 1 33.533 24.939 34.214 24.979 ;
      RECT MASK 1 34.695 24.939 35.376 24.979 ;
      RECT MASK 1 35.857 24.939 36.538 24.979 ;
      RECT MASK 1 38.989 24.939 39.67 24.979 ;
      RECT MASK 1 40.151 24.939 40.832 24.979 ;
      RECT MASK 1 41.313 24.939 41.994 24.979 ;
      RECT MASK 1 42.475 24.939 43.156 24.979 ;
      RECT MASK 1 45.607 24.939 46.288 24.979 ;
      RECT MASK 1 46.769 24.939 47.45 24.979 ;
      RECT MASK 1 47.931 24.939 48.612 24.979 ;
      RECT MASK 1 49.093 24.939 49.774 24.979 ;
      RECT MASK 1 52.225 24.939 52.906 24.979 ;
      RECT MASK 1 53.387 24.939 54.068 24.979 ;
      RECT MASK 1 54.549 24.939 55.23 24.979 ;
      RECT MASK 1 55.711 24.939 56.392 24.979 ;
      RECT MASK 1 58.843 24.939 59.524 24.979 ;
      RECT MASK 1 60.005 24.939 60.686 24.979 ;
      RECT MASK 1 61.167 24.939 61.848 24.979 ;
      RECT MASK 1 62.329 24.939 63.01 24.979 ;
      RECT MASK 1 65.461 24.939 66.142 24.979 ;
      RECT MASK 1 66.623 24.939 67.304 24.979 ;
      RECT MASK 1 67.785 24.939 68.466 24.979 ;
      RECT MASK 1 68.947 24.939 69.628 24.979 ;
      RECT MASK 1 72.079 24.939 72.76 24.979 ;
      RECT MASK 1 73.241 24.939 73.922 24.979 ;
      RECT MASK 1 74.403 24.939 75.084 24.979 ;
      RECT MASK 1 75.565 24.939 76.246 24.979 ;
      RECT MASK 1 78.697 24.939 79.378 24.979 ;
      RECT MASK 1 79.859 24.939 80.54 24.979 ;
      RECT MASK 1 81.021 24.939 81.702 24.979 ;
      RECT MASK 1 82.183 24.939 82.864 24.979 ;
      RECT MASK 1 85.315 24.939 85.996 24.979 ;
      RECT MASK 1 86.477 24.939 87.158 24.979 ;
      RECT MASK 1 87.639 24.939 88.32 24.979 ;
      RECT MASK 1 88.801 24.939 89.482 24.979 ;
      RECT MASK 1 91.933 24.939 92.614 24.979 ;
      RECT MASK 1 93.095 24.939 93.776 24.979 ;
      RECT MASK 1 94.257 24.939 94.938 24.979 ;
      RECT MASK 1 95.419 24.939 96.1 24.979 ;
      RECT MASK 1 98.551 24.939 99.232 24.979 ;
      RECT MASK 1 99.713 24.939 100.394 24.979 ;
      RECT MASK 1 100.875 24.939 101.556 24.979 ;
      RECT MASK 1 102.037 24.939 102.718 24.979 ;
      RECT MASK 1 105.169 24.939 105.85 24.979 ;
      RECT MASK 1 106.331 24.939 107.012 24.979 ;
      RECT MASK 1 107.493 24.939 108.174 24.979 ;
      RECT MASK 1 108.655 24.939 109.336 24.979 ;
      RECT MASK 1 5.821 25.167 5.901 25.394 ;
      RECT MASK 1 6.153 25.167 6.233 25.394 ;
      RECT MASK 1 6.983 25.167 7.063 25.394 ;
      RECT MASK 1 7.315 25.167 7.395 25.394 ;
      RECT MASK 1 8.145 25.167 8.225 25.394 ;
      RECT MASK 1 8.477 25.167 8.557 25.394 ;
      RECT MASK 1 9.307 25.167 9.387 25.394 ;
      RECT MASK 1 9.639 25.167 9.719 25.394 ;
      RECT MASK 1 12.439 25.167 12.519 25.394 ;
      RECT MASK 1 12.771 25.167 12.851 25.394 ;
      RECT MASK 1 13.601 25.167 13.681 25.394 ;
      RECT MASK 1 13.933 25.167 14.013 25.394 ;
      RECT MASK 1 14.763 25.167 14.843 25.394 ;
      RECT MASK 1 15.095 25.167 15.175 25.394 ;
      RECT MASK 1 15.925 25.167 16.005 25.394 ;
      RECT MASK 1 16.257 25.167 16.337 25.394 ;
      RECT MASK 1 19.057 25.167 19.137 25.394 ;
      RECT MASK 1 19.389 25.167 19.469 25.394 ;
      RECT MASK 1 20.219 25.167 20.299 25.394 ;
      RECT MASK 1 20.551 25.167 20.631 25.394 ;
      RECT MASK 1 21.381 25.167 21.461 25.394 ;
      RECT MASK 1 21.713 25.167 21.793 25.394 ;
      RECT MASK 1 22.543 25.167 22.623 25.394 ;
      RECT MASK 1 22.875 25.167 22.955 25.394 ;
      RECT MASK 1 25.675 25.167 25.755 25.394 ;
      RECT MASK 1 26.007 25.167 26.087 25.394 ;
      RECT MASK 1 26.837 25.167 26.917 25.394 ;
      RECT MASK 1 27.169 25.167 27.249 25.394 ;
      RECT MASK 1 27.999 25.167 28.079 25.394 ;
      RECT MASK 1 28.331 25.167 28.411 25.394 ;
      RECT MASK 1 29.161 25.167 29.241 25.394 ;
      RECT MASK 1 29.493 25.167 29.573 25.394 ;
      RECT MASK 1 32.293 25.167 32.373 25.394 ;
      RECT MASK 1 32.625 25.167 32.705 25.394 ;
      RECT MASK 1 33.455 25.167 33.535 25.394 ;
      RECT MASK 1 33.787 25.167 33.867 25.394 ;
      RECT MASK 1 34.617 25.167 34.697 25.394 ;
      RECT MASK 1 34.949 25.167 35.029 25.394 ;
      RECT MASK 1 35.779 25.167 35.859 25.394 ;
      RECT MASK 1 36.111 25.167 36.191 25.394 ;
      RECT MASK 1 38.911 25.167 38.991 25.394 ;
      RECT MASK 1 39.243 25.167 39.323 25.394 ;
      RECT MASK 1 40.073 25.167 40.153 25.394 ;
      RECT MASK 1 40.405 25.167 40.485 25.394 ;
      RECT MASK 1 41.235 25.167 41.315 25.394 ;
      RECT MASK 1 41.567 25.167 41.647 25.394 ;
      RECT MASK 1 42.397 25.167 42.477 25.394 ;
      RECT MASK 1 42.729 25.167 42.809 25.394 ;
      RECT MASK 1 45.529 25.167 45.609 25.394 ;
      RECT MASK 1 45.861 25.167 45.941 25.394 ;
      RECT MASK 1 46.691 25.167 46.771 25.394 ;
      RECT MASK 1 47.023 25.167 47.103 25.394 ;
      RECT MASK 1 47.853 25.167 47.933 25.394 ;
      RECT MASK 1 48.185 25.167 48.265 25.394 ;
      RECT MASK 1 49.015 25.167 49.095 25.394 ;
      RECT MASK 1 49.347 25.167 49.427 25.394 ;
      RECT MASK 1 52.147 25.167 52.227 25.394 ;
      RECT MASK 1 52.479 25.167 52.559 25.394 ;
      RECT MASK 1 53.309 25.167 53.389 25.394 ;
      RECT MASK 1 53.641 25.167 53.721 25.394 ;
      RECT MASK 1 54.471 25.167 54.551 25.394 ;
      RECT MASK 1 54.803 25.167 54.883 25.394 ;
      RECT MASK 1 55.633 25.167 55.713 25.394 ;
      RECT MASK 1 55.965 25.167 56.045 25.394 ;
      RECT MASK 1 58.765 25.167 58.845 25.394 ;
      RECT MASK 1 59.097 25.167 59.177 25.394 ;
      RECT MASK 1 59.927 25.167 60.007 25.394 ;
      RECT MASK 1 60.259 25.167 60.339 25.394 ;
      RECT MASK 1 61.089 25.167 61.169 25.394 ;
      RECT MASK 1 61.421 25.167 61.501 25.394 ;
      RECT MASK 1 62.251 25.167 62.331 25.394 ;
      RECT MASK 1 62.583 25.167 62.663 25.394 ;
      RECT MASK 1 65.383 25.167 65.463 25.394 ;
      RECT MASK 1 65.715 25.167 65.795 25.394 ;
      RECT MASK 1 66.545 25.167 66.625 25.394 ;
      RECT MASK 1 66.877 25.167 66.957 25.394 ;
      RECT MASK 1 67.707 25.167 67.787 25.394 ;
      RECT MASK 1 68.039 25.167 68.119 25.394 ;
      RECT MASK 1 68.869 25.167 68.949 25.394 ;
      RECT MASK 1 69.201 25.167 69.281 25.394 ;
      RECT MASK 1 72.001 25.167 72.081 25.394 ;
      RECT MASK 1 72.333 25.167 72.413 25.394 ;
      RECT MASK 1 73.163 25.167 73.243 25.394 ;
      RECT MASK 1 73.495 25.167 73.575 25.394 ;
      RECT MASK 1 74.325 25.167 74.405 25.394 ;
      RECT MASK 1 74.657 25.167 74.737 25.394 ;
      RECT MASK 1 75.487 25.167 75.567 25.394 ;
      RECT MASK 1 75.819 25.167 75.899 25.394 ;
      RECT MASK 1 78.619 25.167 78.699 25.394 ;
      RECT MASK 1 78.951 25.167 79.031 25.394 ;
      RECT MASK 1 79.781 25.167 79.861 25.394 ;
      RECT MASK 1 80.113 25.167 80.193 25.394 ;
      RECT MASK 1 80.943 25.167 81.023 25.394 ;
      RECT MASK 1 81.275 25.167 81.355 25.394 ;
      RECT MASK 1 82.105 25.167 82.185 25.394 ;
      RECT MASK 1 82.437 25.167 82.517 25.394 ;
      RECT MASK 1 85.237 25.167 85.317 25.394 ;
      RECT MASK 1 85.569 25.167 85.649 25.394 ;
      RECT MASK 1 86.399 25.167 86.479 25.394 ;
      RECT MASK 1 86.731 25.167 86.811 25.394 ;
      RECT MASK 1 87.561 25.167 87.641 25.394 ;
      RECT MASK 1 87.893 25.167 87.973 25.394 ;
      RECT MASK 1 88.723 25.167 88.803 25.394 ;
      RECT MASK 1 89.055 25.167 89.135 25.394 ;
      RECT MASK 1 91.855 25.167 91.935 25.394 ;
      RECT MASK 1 92.187 25.167 92.267 25.394 ;
      RECT MASK 1 93.017 25.167 93.097 25.394 ;
      RECT MASK 1 93.349 25.167 93.429 25.394 ;
      RECT MASK 1 94.179 25.167 94.259 25.394 ;
      RECT MASK 1 94.511 25.167 94.591 25.394 ;
      RECT MASK 1 95.341 25.167 95.421 25.394 ;
      RECT MASK 1 95.673 25.167 95.753 25.394 ;
      RECT MASK 1 98.473 25.167 98.553 25.394 ;
      RECT MASK 1 98.805 25.167 98.885 25.394 ;
      RECT MASK 1 99.635 25.167 99.715 25.394 ;
      RECT MASK 1 99.967 25.167 100.047 25.394 ;
      RECT MASK 1 100.797 25.167 100.877 25.394 ;
      RECT MASK 1 101.129 25.167 101.209 25.394 ;
      RECT MASK 1 101.959 25.167 102.039 25.394 ;
      RECT MASK 1 102.291 25.167 102.371 25.394 ;
      RECT MASK 1 105.091 25.167 105.171 25.394 ;
      RECT MASK 1 105.423 25.167 105.503 25.394 ;
      RECT MASK 1 106.253 25.167 106.333 25.394 ;
      RECT MASK 1 106.585 25.167 106.665 25.394 ;
      RECT MASK 1 107.415 25.167 107.495 25.394 ;
      RECT MASK 1 107.747 25.167 107.827 25.394 ;
      RECT MASK 1 108.577 25.167 108.657 25.394 ;
      RECT MASK 1 108.909 25.167 108.989 25.394 ;
      RECT MASK 1 5.1135 25.795 110.065 25.835 ;
      RECT MASK 1 0.689 26.1 0.769 77.88 ;
      RECT MASK 1 1.31 26.305 113.989 26.345 ;
      RECT MASK 1 115.539 26.545 126.947 26.585 ;
      RECT MASK 1 1.341 26.5545 1.421 77.3665 ;
      RECT MASK 1 113.889 26.6135 113.969 31.08 ;
      RECT MASK 1 115.559 26.8535 115.639 30.0865 ;
      RECT MASK 1 126.847 26.8535 126.927 30.0865 ;
      RECT MASK 1 116.277 27.028 126.675 27.068 ;
      RECT MASK 1 116.271 27.188 116.331 27.412 ;
      RECT MASK 1 116.603 27.188 116.663 27.412 ;
      RECT MASK 1 116.935 27.188 116.995 27.412 ;
      RECT MASK 1 117.267 27.188 117.327 27.412 ;
      RECT MASK 1 117.599 27.188 117.659 27.412 ;
      RECT MASK 1 117.931 27.188 117.991 27.412 ;
      RECT MASK 1 118.263 27.188 118.323 27.412 ;
      RECT MASK 1 118.595 27.188 118.655 27.412 ;
      RECT MASK 1 118.927 27.188 118.987 27.412 ;
      RECT MASK 1 119.259 27.188 119.319 27.412 ;
      RECT MASK 1 119.591 27.188 119.651 27.412 ;
      RECT MASK 1 119.923 27.188 119.983 27.412 ;
      RECT MASK 1 120.255 27.188 120.315 27.412 ;
      RECT MASK 1 120.587 27.188 120.647 27.412 ;
      RECT MASK 1 120.919 27.188 120.979 27.412 ;
      RECT MASK 1 121.251 27.188 121.311 27.412 ;
      RECT MASK 1 121.583 27.188 121.643 27.412 ;
      RECT MASK 1 121.915 27.188 121.975 27.412 ;
      RECT MASK 1 122.247 27.188 122.307 27.412 ;
      RECT MASK 1 122.579 27.188 122.639 27.412 ;
      RECT MASK 1 122.911 27.188 122.971 27.412 ;
      RECT MASK 1 123.243 27.188 123.303 27.412 ;
      RECT MASK 1 123.575 27.188 123.635 27.412 ;
      RECT MASK 1 123.907 27.188 123.967 27.412 ;
      RECT MASK 1 124.239 27.188 124.299 27.412 ;
      RECT MASK 1 124.571 27.188 124.631 27.412 ;
      RECT MASK 1 124.903 27.188 124.963 27.412 ;
      RECT MASK 1 125.235 27.188 125.295 27.412 ;
      RECT MASK 1 125.567 27.188 125.627 27.412 ;
      RECT MASK 1 125.899 27.188 125.959 27.412 ;
      RECT MASK 1 126.231 27.188 126.291 27.412 ;
      RECT MASK 1 116.277 27.808 126.675 27.848 ;
      RECT MASK 1 116.271 27.968 116.331 28.192 ;
      RECT MASK 1 116.603 27.968 116.663 28.192 ;
      RECT MASK 1 116.935 27.968 116.995 28.192 ;
      RECT MASK 1 117.267 27.968 117.327 28.192 ;
      RECT MASK 1 117.599 27.968 117.659 28.192 ;
      RECT MASK 1 117.931 27.968 117.991 28.192 ;
      RECT MASK 1 118.263 27.968 118.323 28.192 ;
      RECT MASK 1 118.595 27.968 118.655 28.192 ;
      RECT MASK 1 118.927 27.968 118.987 28.192 ;
      RECT MASK 1 119.259 27.968 119.319 28.192 ;
      RECT MASK 1 119.591 27.968 119.651 28.192 ;
      RECT MASK 1 119.923 27.968 119.983 28.192 ;
      RECT MASK 1 120.255 27.968 120.315 28.192 ;
      RECT MASK 1 120.587 27.968 120.647 28.192 ;
      RECT MASK 1 120.919 27.968 120.979 28.192 ;
      RECT MASK 1 121.251 27.968 121.311 28.192 ;
      RECT MASK 1 121.583 27.968 121.643 28.192 ;
      RECT MASK 1 121.915 27.968 121.975 28.192 ;
      RECT MASK 1 122.247 27.968 122.307 28.192 ;
      RECT MASK 1 122.579 27.968 122.639 28.192 ;
      RECT MASK 1 122.911 27.968 122.971 28.192 ;
      RECT MASK 1 123.243 27.968 123.303 28.192 ;
      RECT MASK 1 123.575 27.968 123.635 28.192 ;
      RECT MASK 1 123.907 27.968 123.967 28.192 ;
      RECT MASK 1 124.239 27.968 124.299 28.192 ;
      RECT MASK 1 124.571 27.968 124.631 28.192 ;
      RECT MASK 1 124.903 27.968 124.963 28.192 ;
      RECT MASK 1 125.235 27.968 125.295 28.192 ;
      RECT MASK 1 125.567 27.968 125.627 28.192 ;
      RECT MASK 1 125.899 27.968 125.959 28.192 ;
      RECT MASK 1 126.231 27.968 126.291 28.192 ;
      RECT MASK 1 116.277 28.588 126.675 28.628 ;
      RECT MASK 1 116.271 28.748 116.331 28.972 ;
      RECT MASK 1 116.603 28.748 116.663 28.972 ;
      RECT MASK 1 116.935 28.748 116.995 28.972 ;
      RECT MASK 1 117.267 28.748 117.327 28.972 ;
      RECT MASK 1 117.599 28.748 117.659 28.972 ;
      RECT MASK 1 117.931 28.748 117.991 28.972 ;
      RECT MASK 1 118.263 28.748 118.323 28.972 ;
      RECT MASK 1 118.595 28.748 118.655 28.972 ;
      RECT MASK 1 118.927 28.748 118.987 28.972 ;
      RECT MASK 1 119.259 28.748 119.319 28.972 ;
      RECT MASK 1 119.591 28.748 119.651 28.972 ;
      RECT MASK 1 119.923 28.748 119.983 28.972 ;
      RECT MASK 1 120.255 28.748 120.315 28.972 ;
      RECT MASK 1 120.587 28.748 120.647 28.972 ;
      RECT MASK 1 120.919 28.748 120.979 28.972 ;
      RECT MASK 1 121.251 28.748 121.311 28.972 ;
      RECT MASK 1 121.583 28.748 121.643 28.972 ;
      RECT MASK 1 121.915 28.748 121.975 28.972 ;
      RECT MASK 1 122.247 28.748 122.307 28.972 ;
      RECT MASK 1 122.579 28.748 122.639 28.972 ;
      RECT MASK 1 122.911 28.748 122.971 28.972 ;
      RECT MASK 1 123.243 28.748 123.303 28.972 ;
      RECT MASK 1 123.575 28.748 123.635 28.972 ;
      RECT MASK 1 123.907 28.748 123.967 28.972 ;
      RECT MASK 1 124.239 28.748 124.299 28.972 ;
      RECT MASK 1 124.571 28.748 124.631 28.972 ;
      RECT MASK 1 124.903 28.748 124.963 28.972 ;
      RECT MASK 1 125.235 28.748 125.295 28.972 ;
      RECT MASK 1 125.567 28.748 125.627 28.972 ;
      RECT MASK 1 125.899 28.748 125.959 28.972 ;
      RECT MASK 1 126.231 28.748 126.291 28.972 ;
      RECT MASK 1 116.277 29.368 126.683 29.408 ;
      RECT MASK 1 116.271 29.528 116.331 29.752 ;
      RECT MASK 1 116.603 29.528 116.663 29.752 ;
      RECT MASK 1 116.935 29.528 116.995 29.752 ;
      RECT MASK 1 117.267 29.528 117.327 29.752 ;
      RECT MASK 1 117.599 29.528 117.659 29.752 ;
      RECT MASK 1 117.931 29.528 117.991 29.752 ;
      RECT MASK 1 118.263 29.528 118.323 29.752 ;
      RECT MASK 1 118.595 29.528 118.655 29.752 ;
      RECT MASK 1 118.927 29.528 118.987 29.752 ;
      RECT MASK 1 119.259 29.528 119.319 29.752 ;
      RECT MASK 1 119.591 29.528 119.651 29.752 ;
      RECT MASK 1 119.923 29.528 119.983 29.752 ;
      RECT MASK 1 120.255 29.528 120.315 29.752 ;
      RECT MASK 1 120.587 29.528 120.647 29.752 ;
      RECT MASK 1 120.919 29.528 120.979 29.752 ;
      RECT MASK 1 121.251 29.528 121.311 29.752 ;
      RECT MASK 1 121.583 29.528 121.643 29.752 ;
      RECT MASK 1 121.915 29.528 121.975 29.752 ;
      RECT MASK 1 122.247 29.528 122.307 29.752 ;
      RECT MASK 1 122.579 29.528 122.639 29.752 ;
      RECT MASK 1 122.911 29.528 122.971 29.752 ;
      RECT MASK 1 123.243 29.528 123.303 29.752 ;
      RECT MASK 1 123.575 29.528 123.635 29.752 ;
      RECT MASK 1 123.907 29.528 123.967 29.752 ;
      RECT MASK 1 124.239 29.528 124.299 29.752 ;
      RECT MASK 1 124.571 29.528 124.631 29.752 ;
      RECT MASK 1 124.903 29.528 124.963 29.752 ;
      RECT MASK 1 125.235 29.528 125.295 29.752 ;
      RECT MASK 1 125.567 29.528 125.627 29.752 ;
      RECT MASK 1 125.899 29.528 125.959 29.752 ;
      RECT MASK 1 126.231 29.528 126.291 29.752 ;
      RECT MASK 1 115.539 30.355 126.947 30.395 ;
      RECT MASK 1 113.869 31.285 129.1075 31.325 ;
      RECT MASK 1 128.995 31.5935 129.075 72.1165 ;
      RECT MASK 1 1.9425 33.37 41.8765 33.41 ;
      RECT MASK 1 42.6605 33.37 82.5945 33.41 ;
      RECT MASK 1 83.4005 33.37 128.3145 33.41 ;
      RECT MASK 1 1.9425 33.79 41.8765 33.83 ;
      RECT MASK 1 42.6605 33.79 82.5945 33.83 ;
      RECT MASK 1 83.4005 33.79 128.3145 33.83 ;
      RECT MASK 1 1.9425 39.46 41.8765 39.5 ;
      RECT MASK 1 42.6605 39.46 82.5945 39.5 ;
      RECT MASK 1 83.4005 39.46 128.3145 39.5 ;
      RECT MASK 1 1.9425 39.88 41.8765 39.92 ;
      RECT MASK 1 42.6605 39.88 82.5945 39.92 ;
      RECT MASK 1 83.4005 39.88 128.3145 39.92 ;
      RECT MASK 1 1.9425 45.58 41.8765 45.62 ;
      RECT MASK 1 42.6605 45.58 82.5945 45.62 ;
      RECT MASK 1 83.4005 45.58 128.3145 45.62 ;
      RECT MASK 1 1.9425 46 41.8765 46.04 ;
      RECT MASK 1 42.6605 46 82.5945 46.04 ;
      RECT MASK 1 83.4005 46 128.3145 46.04 ;
      RECT MASK 1 1.9425 51.7 41.8765 51.74 ;
      RECT MASK 1 42.6605 51.7 82.5945 51.74 ;
      RECT MASK 1 83.4005 51.7 128.3145 51.74 ;
      RECT MASK 1 1.9425 52.12 41.8765 52.16 ;
      RECT MASK 1 42.6605 52.12 82.5945 52.16 ;
      RECT MASK 1 83.4005 52.12 128.3145 52.16 ;
      RECT MASK 1 1.9425 57.82 41.8765 57.86 ;
      RECT MASK 1 42.6605 57.82 82.5945 57.86 ;
      RECT MASK 1 83.4005 57.82 128.3145 57.86 ;
      RECT MASK 1 1.9425 58.24 41.8765 58.28 ;
      RECT MASK 1 42.6605 58.24 82.5945 58.28 ;
      RECT MASK 1 83.4005 58.24 128.3145 58.28 ;
      RECT MASK 1 1.9425 63.94 41.8765 63.98 ;
      RECT MASK 1 42.6605 63.94 82.5945 63.98 ;
      RECT MASK 1 83.4005 63.94 128.3145 63.98 ;
      RECT MASK 1 1.9425 64.36 41.8765 64.4 ;
      RECT MASK 1 42.6605 64.36 82.5945 64.4 ;
      RECT MASK 1 83.4005 64.36 128.3145 64.4 ;
      RECT MASK 1 1.9425 70.06 41.8765 70.1 ;
      RECT MASK 1 42.6605 70.06 82.5945 70.1 ;
      RECT MASK 1 83.4005 70.06 128.3145 70.1 ;
      RECT MASK 1 1.9425 70.48 41.8765 70.52 ;
      RECT MASK 1 42.6605 70.48 82.5945 70.52 ;
      RECT MASK 1 83.4005 70.48 128.3145 70.52 ;
      RECT MASK 1 113.869 72.385 129.095 72.425 ;
      RECT MASK 1 113.889 72.63 113.969 77.3665 ;
      RECT MASK 1 114.345 72.865 129.322 72.905 ;
      RECT MASK 1 114.461 73.11 114.541 78.51 ;
      RECT MASK 1 115.539 73.345 126.947 73.385 ;
      RECT MASK 1 115.559 73.6535 115.639 80.0065 ;
      RECT MASK 1 126.847 73.6535 126.927 80.0065 ;
      RECT MASK 1 116.271 73.988 116.331 74.212 ;
      RECT MASK 1 116.603 73.988 116.663 74.212 ;
      RECT MASK 1 116.935 73.988 116.995 74.212 ;
      RECT MASK 1 117.267 73.988 117.327 74.212 ;
      RECT MASK 1 117.599 73.988 117.659 74.212 ;
      RECT MASK 1 117.931 73.988 117.991 74.212 ;
      RECT MASK 1 118.263 73.988 118.323 74.212 ;
      RECT MASK 1 118.595 73.988 118.655 74.212 ;
      RECT MASK 1 118.927 73.988 118.987 74.212 ;
      RECT MASK 1 119.259 73.988 119.319 74.212 ;
      RECT MASK 1 119.591 73.988 119.651 74.212 ;
      RECT MASK 1 119.923 73.988 119.983 74.212 ;
      RECT MASK 1 120.255 73.988 120.315 74.212 ;
      RECT MASK 1 120.587 73.988 120.647 74.212 ;
      RECT MASK 1 120.919 73.988 120.979 74.212 ;
      RECT MASK 1 121.251 73.988 121.311 74.212 ;
      RECT MASK 1 121.583 73.988 121.643 74.212 ;
      RECT MASK 1 121.915 73.988 121.975 74.212 ;
      RECT MASK 1 122.247 73.988 122.307 74.212 ;
      RECT MASK 1 122.579 73.988 122.639 74.212 ;
      RECT MASK 1 122.911 73.988 122.971 74.212 ;
      RECT MASK 1 123.243 73.988 123.303 74.212 ;
      RECT MASK 1 123.575 73.988 123.635 74.212 ;
      RECT MASK 1 123.907 73.988 123.967 74.212 ;
      RECT MASK 1 124.239 73.988 124.299 74.212 ;
      RECT MASK 1 124.571 73.988 124.631 74.212 ;
      RECT MASK 1 124.903 73.988 124.963 74.212 ;
      RECT MASK 1 125.235 73.988 125.295 74.212 ;
      RECT MASK 1 125.567 73.988 125.627 74.212 ;
      RECT MASK 1 125.899 73.988 125.959 74.212 ;
      RECT MASK 1 126.231 73.988 126.291 74.212 ;
      RECT MASK 1 116.339 74.332 126.649 74.372 ;
      RECT MASK 1 116.271 74.768 116.331 74.992 ;
      RECT MASK 1 116.603 74.768 116.663 74.992 ;
      RECT MASK 1 116.935 74.768 116.995 74.992 ;
      RECT MASK 1 117.267 74.768 117.327 74.992 ;
      RECT MASK 1 117.599 74.768 117.659 74.992 ;
      RECT MASK 1 117.931 74.768 117.991 74.992 ;
      RECT MASK 1 118.263 74.768 118.323 74.992 ;
      RECT MASK 1 118.595 74.768 118.655 74.992 ;
      RECT MASK 1 118.927 74.768 118.987 74.992 ;
      RECT MASK 1 119.259 74.768 119.319 74.992 ;
      RECT MASK 1 119.591 74.768 119.651 74.992 ;
      RECT MASK 1 119.923 74.768 119.983 74.992 ;
      RECT MASK 1 120.255 74.768 120.315 74.992 ;
      RECT MASK 1 120.587 74.768 120.647 74.992 ;
      RECT MASK 1 120.919 74.768 120.979 74.992 ;
      RECT MASK 1 121.251 74.768 121.311 74.992 ;
      RECT MASK 1 121.583 74.768 121.643 74.992 ;
      RECT MASK 1 121.915 74.768 121.975 74.992 ;
      RECT MASK 1 122.247 74.768 122.307 74.992 ;
      RECT MASK 1 122.579 74.768 122.639 74.992 ;
      RECT MASK 1 122.911 74.768 122.971 74.992 ;
      RECT MASK 1 123.243 74.768 123.303 74.992 ;
      RECT MASK 1 123.575 74.768 123.635 74.992 ;
      RECT MASK 1 123.907 74.768 123.967 74.992 ;
      RECT MASK 1 124.239 74.768 124.299 74.992 ;
      RECT MASK 1 124.571 74.768 124.631 74.992 ;
      RECT MASK 1 124.903 74.768 124.963 74.992 ;
      RECT MASK 1 125.235 74.768 125.295 74.992 ;
      RECT MASK 1 125.567 74.768 125.627 74.992 ;
      RECT MASK 1 125.899 74.768 125.959 74.992 ;
      RECT MASK 1 126.231 74.768 126.291 74.992 ;
      RECT MASK 1 116.339 75.112 126.649 75.152 ;
      RECT MASK 1 116.271 75.548 116.331 75.772 ;
      RECT MASK 1 116.603 75.548 116.663 75.772 ;
      RECT MASK 1 116.935 75.548 116.995 75.772 ;
      RECT MASK 1 117.267 75.548 117.327 75.772 ;
      RECT MASK 1 117.599 75.548 117.659 75.772 ;
      RECT MASK 1 117.931 75.548 117.991 75.772 ;
      RECT MASK 1 118.263 75.548 118.323 75.772 ;
      RECT MASK 1 118.595 75.548 118.655 75.772 ;
      RECT MASK 1 118.927 75.548 118.987 75.772 ;
      RECT MASK 1 119.259 75.548 119.319 75.772 ;
      RECT MASK 1 119.591 75.548 119.651 75.772 ;
      RECT MASK 1 119.923 75.548 119.983 75.772 ;
      RECT MASK 1 120.255 75.548 120.315 75.772 ;
      RECT MASK 1 120.587 75.548 120.647 75.772 ;
      RECT MASK 1 120.919 75.548 120.979 75.772 ;
      RECT MASK 1 121.251 75.548 121.311 75.772 ;
      RECT MASK 1 121.583 75.548 121.643 75.772 ;
      RECT MASK 1 121.915 75.548 121.975 75.772 ;
      RECT MASK 1 122.247 75.548 122.307 75.772 ;
      RECT MASK 1 122.579 75.548 122.639 75.772 ;
      RECT MASK 1 122.911 75.548 122.971 75.772 ;
      RECT MASK 1 123.243 75.548 123.303 75.772 ;
      RECT MASK 1 123.575 75.548 123.635 75.772 ;
      RECT MASK 1 123.907 75.548 123.967 75.772 ;
      RECT MASK 1 124.239 75.548 124.299 75.772 ;
      RECT MASK 1 124.571 75.548 124.631 75.772 ;
      RECT MASK 1 124.903 75.548 124.963 75.772 ;
      RECT MASK 1 125.235 75.548 125.295 75.772 ;
      RECT MASK 1 125.567 75.548 125.627 75.772 ;
      RECT MASK 1 125.899 75.548 125.959 75.772 ;
      RECT MASK 1 126.231 75.548 126.291 75.772 ;
      RECT MASK 1 116.3385 75.892 126.649 75.932 ;
      RECT MASK 1 116.271 76.328 116.331 76.552 ;
      RECT MASK 1 116.603 76.328 116.663 76.552 ;
      RECT MASK 1 116.935 76.328 116.995 76.552 ;
      RECT MASK 1 117.267 76.328 117.327 76.552 ;
      RECT MASK 1 117.599 76.328 117.659 76.552 ;
      RECT MASK 1 117.931 76.328 117.991 76.552 ;
      RECT MASK 1 118.263 76.328 118.323 76.552 ;
      RECT MASK 1 118.595 76.328 118.655 76.552 ;
      RECT MASK 1 118.927 76.328 118.987 76.552 ;
      RECT MASK 1 119.259 76.328 119.319 76.552 ;
      RECT MASK 1 119.591 76.328 119.651 76.552 ;
      RECT MASK 1 119.923 76.328 119.983 76.552 ;
      RECT MASK 1 120.255 76.328 120.315 76.552 ;
      RECT MASK 1 120.587 76.328 120.647 76.552 ;
      RECT MASK 1 120.919 76.328 120.979 76.552 ;
      RECT MASK 1 121.251 76.328 121.311 76.552 ;
      RECT MASK 1 121.583 76.328 121.643 76.552 ;
      RECT MASK 1 121.915 76.328 121.975 76.552 ;
      RECT MASK 1 122.247 76.328 122.307 76.552 ;
      RECT MASK 1 122.579 76.328 122.639 76.552 ;
      RECT MASK 1 122.911 76.328 122.971 76.552 ;
      RECT MASK 1 123.243 76.328 123.303 76.552 ;
      RECT MASK 1 123.575 76.328 123.635 76.552 ;
      RECT MASK 1 123.907 76.328 123.967 76.552 ;
      RECT MASK 1 124.239 76.328 124.299 76.552 ;
      RECT MASK 1 124.571 76.328 124.631 76.552 ;
      RECT MASK 1 124.903 76.328 124.963 76.552 ;
      RECT MASK 1 125.235 76.328 125.295 76.552 ;
      RECT MASK 1 125.567 76.328 125.627 76.552 ;
      RECT MASK 1 125.899 76.328 125.959 76.552 ;
      RECT MASK 1 126.231 76.328 126.291 76.552 ;
      RECT MASK 1 116.339 76.672 126.649 76.712 ;
      RECT MASK 1 116.271 77.108 116.331 77.332 ;
      RECT MASK 1 116.603 77.108 116.663 77.332 ;
      RECT MASK 1 116.935 77.108 116.995 77.332 ;
      RECT MASK 1 117.267 77.108 117.327 77.332 ;
      RECT MASK 1 117.599 77.108 117.659 77.332 ;
      RECT MASK 1 117.931 77.108 117.991 77.332 ;
      RECT MASK 1 118.263 77.108 118.323 77.332 ;
      RECT MASK 1 118.595 77.108 118.655 77.332 ;
      RECT MASK 1 118.927 77.108 118.987 77.332 ;
      RECT MASK 1 119.259 77.108 119.319 77.332 ;
      RECT MASK 1 119.591 77.108 119.651 77.332 ;
      RECT MASK 1 119.923 77.108 119.983 77.332 ;
      RECT MASK 1 120.255 77.108 120.315 77.332 ;
      RECT MASK 1 120.587 77.108 120.647 77.332 ;
      RECT MASK 1 120.919 77.108 120.979 77.332 ;
      RECT MASK 1 121.251 77.108 121.311 77.332 ;
      RECT MASK 1 121.583 77.108 121.643 77.332 ;
      RECT MASK 1 121.915 77.108 121.975 77.332 ;
      RECT MASK 1 122.247 77.108 122.307 77.332 ;
      RECT MASK 1 122.579 77.108 122.639 77.332 ;
      RECT MASK 1 122.911 77.108 122.971 77.332 ;
      RECT MASK 1 123.243 77.108 123.303 77.332 ;
      RECT MASK 1 123.575 77.108 123.635 77.332 ;
      RECT MASK 1 123.907 77.108 123.967 77.332 ;
      RECT MASK 1 124.239 77.108 124.299 77.332 ;
      RECT MASK 1 124.571 77.108 124.631 77.332 ;
      RECT MASK 1 124.903 77.108 124.963 77.332 ;
      RECT MASK 1 125.235 77.108 125.295 77.332 ;
      RECT MASK 1 125.567 77.108 125.627 77.332 ;
      RECT MASK 1 125.899 77.108 125.959 77.332 ;
      RECT MASK 1 126.231 77.108 126.291 77.332 ;
      RECT MASK 1 116.339 77.452 126.651 77.492 ;
      RECT MASK 1 1.31 77.635 113.984 77.675 ;
      RECT MASK 1 116.271 77.888 116.331 78.112 ;
      RECT MASK 1 116.603 77.888 116.663 78.112 ;
      RECT MASK 1 116.935 77.888 116.995 78.112 ;
      RECT MASK 1 117.267 77.888 117.327 78.112 ;
      RECT MASK 1 117.599 77.888 117.659 78.112 ;
      RECT MASK 1 117.931 77.888 117.991 78.112 ;
      RECT MASK 1 118.263 77.888 118.323 78.112 ;
      RECT MASK 1 118.595 77.888 118.655 78.112 ;
      RECT MASK 1 118.927 77.888 118.987 78.112 ;
      RECT MASK 1 119.259 77.888 119.319 78.112 ;
      RECT MASK 1 119.591 77.888 119.651 78.112 ;
      RECT MASK 1 119.923 77.888 119.983 78.112 ;
      RECT MASK 1 120.255 77.888 120.315 78.112 ;
      RECT MASK 1 120.587 77.888 120.647 78.112 ;
      RECT MASK 1 120.919 77.888 120.979 78.112 ;
      RECT MASK 1 121.251 77.888 121.311 78.112 ;
      RECT MASK 1 121.583 77.888 121.643 78.112 ;
      RECT MASK 1 121.915 77.888 121.975 78.112 ;
      RECT MASK 1 122.247 77.888 122.307 78.112 ;
      RECT MASK 1 122.579 77.888 122.639 78.112 ;
      RECT MASK 1 122.911 77.888 122.971 78.112 ;
      RECT MASK 1 123.243 77.888 123.303 78.112 ;
      RECT MASK 1 123.575 77.888 123.635 78.112 ;
      RECT MASK 1 123.907 77.888 123.967 78.112 ;
      RECT MASK 1 124.239 77.888 124.299 78.112 ;
      RECT MASK 1 124.571 77.888 124.631 78.112 ;
      RECT MASK 1 124.903 77.888 124.963 78.112 ;
      RECT MASK 1 125.235 77.888 125.295 78.112 ;
      RECT MASK 1 125.567 77.888 125.627 78.112 ;
      RECT MASK 1 125.899 77.888 125.959 78.112 ;
      RECT MASK 1 126.231 77.888 126.291 78.112 ;
      RECT MASK 1 6.224 78.145 110.065 78.185 ;
      RECT MASK 1 116.339 78.232 126.65 78.272 ;
      RECT MASK 1 6.319 78.42 6.399 79.838 ;
      RECT MASK 1 10.469 78.42 10.549 79.838 ;
      RECT MASK 1 11.775 78.42 11.855 79.838 ;
      RECT MASK 1 17.087 78.42 17.167 79.838 ;
      RECT MASK 1 18.393 78.42 18.473 79.838 ;
      RECT MASK 1 23.705 78.42 23.785 79.838 ;
      RECT MASK 1 25.011 78.42 25.091 79.838 ;
      RECT MASK 1 30.323 78.42 30.403 79.838 ;
      RECT MASK 1 31.629 78.42 31.709 79.838 ;
      RECT MASK 1 36.941 78.42 37.021 79.838 ;
      RECT MASK 1 38.247 78.42 38.327 79.838 ;
      RECT MASK 1 43.559 78.42 43.639 79.838 ;
      RECT MASK 1 44.865 78.42 44.945 79.838 ;
      RECT MASK 1 50.177 78.42 50.257 79.838 ;
      RECT MASK 1 51.483 78.42 51.563 79.838 ;
      RECT MASK 1 56.795 78.42 56.875 79.838 ;
      RECT MASK 1 58.101 78.42 58.181 79.838 ;
      RECT MASK 1 63.413 78.42 63.493 79.838 ;
      RECT MASK 1 64.719 78.42 64.799 79.838 ;
      RECT MASK 1 70.031 78.42 70.111 79.838 ;
      RECT MASK 1 71.337 78.42 71.417 79.838 ;
      RECT MASK 1 76.649 78.42 76.729 79.838 ;
      RECT MASK 1 77.955 78.42 78.035 79.838 ;
      RECT MASK 1 83.267 78.42 83.347 79.838 ;
      RECT MASK 1 84.573 78.42 84.653 79.838 ;
      RECT MASK 1 89.885 78.42 89.965 79.838 ;
      RECT MASK 1 91.191 78.42 91.271 79.838 ;
      RECT MASK 1 96.503 78.42 96.583 79.838 ;
      RECT MASK 1 97.809 78.42 97.889 79.838 ;
      RECT MASK 1 103.121 78.42 103.201 79.838 ;
      RECT MASK 1 104.427 78.42 104.507 79.838 ;
      RECT MASK 1 109.739 78.42 109.819 79.838 ;
      RECT MASK 1 16.755 78.4895 16.835 78.77 ;
      RECT MASK 1 23.373 78.4895 23.453 78.77 ;
      RECT MASK 1 29.991 78.4895 30.071 78.77 ;
      RECT MASK 1 36.609 78.4895 36.689 78.77 ;
      RECT MASK 1 43.227 78.4895 43.307 78.77 ;
      RECT MASK 1 49.845 78.4895 49.925 78.77 ;
      RECT MASK 1 56.463 78.4895 56.543 78.77 ;
      RECT MASK 1 63.081 78.4895 63.161 78.77 ;
      RECT MASK 1 69.699 78.4895 69.779 78.77 ;
      RECT MASK 1 76.317 78.4895 76.397 78.77 ;
      RECT MASK 1 82.935 78.4895 83.015 78.77 ;
      RECT MASK 1 89.553 78.4895 89.633 78.77 ;
      RECT MASK 1 96.171 78.4895 96.251 78.77 ;
      RECT MASK 1 102.789 78.4895 102.869 78.77 ;
      RECT MASK 1 109.407 78.4895 109.487 78.77 ;
      RECT MASK 1 6.983 78.586 7.063 78.813 ;
      RECT MASK 1 7.315 78.586 7.395 78.813 ;
      RECT MASK 1 8.145 78.586 8.225 78.813 ;
      RECT MASK 1 8.477 78.586 8.557 78.813 ;
      RECT MASK 1 9.307 78.586 9.387 78.813 ;
      RECT MASK 1 9.639 78.586 9.719 78.813 ;
      RECT MASK 1 12.439 78.586 12.519 78.813 ;
      RECT MASK 1 12.771 78.586 12.851 78.813 ;
      RECT MASK 1 13.601 78.586 13.681 78.813 ;
      RECT MASK 1 13.933 78.586 14.013 78.813 ;
      RECT MASK 1 14.763 78.586 14.843 78.813 ;
      RECT MASK 1 15.095 78.586 15.175 78.813 ;
      RECT MASK 1 15.925 78.586 16.005 78.813 ;
      RECT MASK 1 16.257 78.586 16.337 78.813 ;
      RECT MASK 1 19.057 78.586 19.137 78.813 ;
      RECT MASK 1 19.389 78.586 19.469 78.813 ;
      RECT MASK 1 20.219 78.586 20.299 78.813 ;
      RECT MASK 1 20.551 78.586 20.631 78.813 ;
      RECT MASK 1 21.381 78.586 21.461 78.813 ;
      RECT MASK 1 21.713 78.586 21.793 78.813 ;
      RECT MASK 1 22.543 78.586 22.623 78.813 ;
      RECT MASK 1 22.875 78.586 22.955 78.813 ;
      RECT MASK 1 25.675 78.586 25.755 78.813 ;
      RECT MASK 1 26.007 78.586 26.087 78.813 ;
      RECT MASK 1 26.837 78.586 26.917 78.813 ;
      RECT MASK 1 27.169 78.586 27.249 78.813 ;
      RECT MASK 1 27.999 78.586 28.079 78.813 ;
      RECT MASK 1 28.331 78.586 28.411 78.813 ;
      RECT MASK 1 29.161 78.586 29.241 78.813 ;
      RECT MASK 1 29.493 78.586 29.573 78.813 ;
      RECT MASK 1 32.293 78.586 32.373 78.813 ;
      RECT MASK 1 32.625 78.586 32.705 78.813 ;
      RECT MASK 1 33.455 78.586 33.535 78.813 ;
      RECT MASK 1 33.787 78.586 33.867 78.813 ;
      RECT MASK 1 34.617 78.586 34.697 78.813 ;
      RECT MASK 1 34.949 78.586 35.029 78.813 ;
      RECT MASK 1 35.779 78.586 35.859 78.813 ;
      RECT MASK 1 36.111 78.586 36.191 78.813 ;
      RECT MASK 1 38.911 78.586 38.991 78.813 ;
      RECT MASK 1 39.243 78.586 39.323 78.813 ;
      RECT MASK 1 40.073 78.586 40.153 78.813 ;
      RECT MASK 1 40.405 78.586 40.485 78.813 ;
      RECT MASK 1 41.235 78.586 41.315 78.813 ;
      RECT MASK 1 41.567 78.586 41.647 78.813 ;
      RECT MASK 1 42.397 78.586 42.477 78.813 ;
      RECT MASK 1 42.729 78.586 42.809 78.813 ;
      RECT MASK 1 45.529 78.586 45.609 78.813 ;
      RECT MASK 1 45.861 78.586 45.941 78.813 ;
      RECT MASK 1 46.691 78.586 46.771 78.813 ;
      RECT MASK 1 47.023 78.586 47.103 78.813 ;
      RECT MASK 1 47.853 78.586 47.933 78.813 ;
      RECT MASK 1 48.185 78.586 48.265 78.813 ;
      RECT MASK 1 49.015 78.586 49.095 78.813 ;
      RECT MASK 1 49.347 78.586 49.427 78.813 ;
      RECT MASK 1 52.147 78.586 52.227 78.813 ;
      RECT MASK 1 52.479 78.586 52.559 78.813 ;
      RECT MASK 1 53.309 78.586 53.389 78.813 ;
      RECT MASK 1 53.641 78.586 53.721 78.813 ;
      RECT MASK 1 54.471 78.586 54.551 78.813 ;
      RECT MASK 1 54.803 78.586 54.883 78.813 ;
      RECT MASK 1 55.633 78.586 55.713 78.813 ;
      RECT MASK 1 55.965 78.586 56.045 78.813 ;
      RECT MASK 1 58.765 78.586 58.845 78.813 ;
      RECT MASK 1 59.097 78.586 59.177 78.813 ;
      RECT MASK 1 59.927 78.586 60.007 78.813 ;
      RECT MASK 1 60.259 78.586 60.339 78.813 ;
      RECT MASK 1 61.089 78.586 61.169 78.813 ;
      RECT MASK 1 61.421 78.586 61.501 78.813 ;
      RECT MASK 1 62.251 78.586 62.331 78.813 ;
      RECT MASK 1 62.583 78.586 62.663 78.813 ;
      RECT MASK 1 65.383 78.586 65.463 78.813 ;
      RECT MASK 1 65.715 78.586 65.795 78.813 ;
      RECT MASK 1 66.545 78.586 66.625 78.813 ;
      RECT MASK 1 66.877 78.586 66.957 78.813 ;
      RECT MASK 1 67.707 78.586 67.787 78.813 ;
      RECT MASK 1 68.039 78.586 68.119 78.813 ;
      RECT MASK 1 68.869 78.586 68.949 78.813 ;
      RECT MASK 1 69.201 78.586 69.281 78.813 ;
      RECT MASK 1 72.001 78.586 72.081 78.813 ;
      RECT MASK 1 72.333 78.586 72.413 78.813 ;
      RECT MASK 1 73.163 78.586 73.243 78.813 ;
      RECT MASK 1 73.495 78.586 73.575 78.813 ;
      RECT MASK 1 74.325 78.586 74.405 78.813 ;
      RECT MASK 1 74.657 78.586 74.737 78.813 ;
      RECT MASK 1 75.487 78.586 75.567 78.813 ;
      RECT MASK 1 75.819 78.586 75.899 78.813 ;
      RECT MASK 1 78.619 78.586 78.699 78.813 ;
      RECT MASK 1 78.951 78.586 79.031 78.813 ;
      RECT MASK 1 79.781 78.586 79.861 78.813 ;
      RECT MASK 1 80.113 78.586 80.193 78.813 ;
      RECT MASK 1 80.943 78.586 81.023 78.813 ;
      RECT MASK 1 81.275 78.586 81.355 78.813 ;
      RECT MASK 1 82.105 78.586 82.185 78.813 ;
      RECT MASK 1 82.437 78.586 82.517 78.813 ;
      RECT MASK 1 85.237 78.586 85.317 78.813 ;
      RECT MASK 1 85.569 78.586 85.649 78.813 ;
      RECT MASK 1 86.399 78.586 86.479 78.813 ;
      RECT MASK 1 86.731 78.586 86.811 78.813 ;
      RECT MASK 1 87.561 78.586 87.641 78.813 ;
      RECT MASK 1 87.893 78.586 87.973 78.813 ;
      RECT MASK 1 88.723 78.586 88.803 78.813 ;
      RECT MASK 1 89.055 78.586 89.135 78.813 ;
      RECT MASK 1 91.855 78.586 91.935 78.813 ;
      RECT MASK 1 92.187 78.586 92.267 78.813 ;
      RECT MASK 1 93.017 78.586 93.097 78.813 ;
      RECT MASK 1 93.349 78.586 93.429 78.813 ;
      RECT MASK 1 94.179 78.586 94.259 78.813 ;
      RECT MASK 1 94.511 78.586 94.591 78.813 ;
      RECT MASK 1 95.341 78.586 95.421 78.813 ;
      RECT MASK 1 95.673 78.586 95.753 78.813 ;
      RECT MASK 1 98.473 78.586 98.553 78.813 ;
      RECT MASK 1 98.805 78.586 98.885 78.813 ;
      RECT MASK 1 99.635 78.586 99.715 78.813 ;
      RECT MASK 1 99.967 78.586 100.047 78.813 ;
      RECT MASK 1 100.797 78.586 100.877 78.813 ;
      RECT MASK 1 101.129 78.586 101.209 78.813 ;
      RECT MASK 1 101.959 78.586 102.039 78.813 ;
      RECT MASK 1 102.291 78.586 102.371 78.813 ;
      RECT MASK 1 105.091 78.586 105.171 78.813 ;
      RECT MASK 1 105.423 78.586 105.503 78.813 ;
      RECT MASK 1 106.253 78.586 106.333 78.813 ;
      RECT MASK 1 106.585 78.586 106.665 78.813 ;
      RECT MASK 1 107.415 78.586 107.495 78.813 ;
      RECT MASK 1 107.747 78.586 107.827 78.813 ;
      RECT MASK 1 108.577 78.586 108.657 78.813 ;
      RECT MASK 1 108.909 78.586 108.989 78.813 ;
      RECT MASK 1 1.248 78.655 5.362 78.695 ;
      RECT MASK 1 116.271 78.668 116.331 78.892 ;
      RECT MASK 1 116.603 78.668 116.663 78.892 ;
      RECT MASK 1 116.935 78.668 116.995 78.892 ;
      RECT MASK 1 117.267 78.668 117.327 78.892 ;
      RECT MASK 1 117.599 78.668 117.659 78.892 ;
      RECT MASK 1 117.931 78.668 117.991 78.892 ;
      RECT MASK 1 118.263 78.668 118.323 78.892 ;
      RECT MASK 1 118.595 78.668 118.655 78.892 ;
      RECT MASK 1 118.927 78.668 118.987 78.892 ;
      RECT MASK 1 119.259 78.668 119.319 78.892 ;
      RECT MASK 1 119.591 78.668 119.651 78.892 ;
      RECT MASK 1 119.923 78.668 119.983 78.892 ;
      RECT MASK 1 120.255 78.668 120.315 78.892 ;
      RECT MASK 1 120.587 78.668 120.647 78.892 ;
      RECT MASK 1 120.919 78.668 120.979 78.892 ;
      RECT MASK 1 121.251 78.668 121.311 78.892 ;
      RECT MASK 1 121.583 78.668 121.643 78.892 ;
      RECT MASK 1 121.915 78.668 121.975 78.892 ;
      RECT MASK 1 122.247 78.668 122.307 78.892 ;
      RECT MASK 1 122.579 78.668 122.639 78.892 ;
      RECT MASK 1 122.911 78.668 122.971 78.892 ;
      RECT MASK 1 123.243 78.668 123.303 78.892 ;
      RECT MASK 1 123.575 78.668 123.635 78.892 ;
      RECT MASK 1 123.907 78.668 123.967 78.892 ;
      RECT MASK 1 124.239 78.668 124.299 78.892 ;
      RECT MASK 1 124.571 78.668 124.631 78.892 ;
      RECT MASK 1 124.903 78.668 124.963 78.892 ;
      RECT MASK 1 125.235 78.668 125.295 78.892 ;
      RECT MASK 1 125.567 78.668 125.627 78.892 ;
      RECT MASK 1 125.899 78.668 125.959 78.892 ;
      RECT MASK 1 126.231 78.668 126.291 78.892 ;
      RECT MASK 1 111.186 78.895 113.288 78.935 ;
      RECT MASK 1 11.039 78.9455 11.119 79.217 ;
      RECT MASK 1 11.371 78.9455 11.451 79.217 ;
      RECT MASK 1 17.657 78.9455 17.737 79.217 ;
      RECT MASK 1 17.989 78.9455 18.069 79.217 ;
      RECT MASK 1 24.275 78.9455 24.355 79.217 ;
      RECT MASK 1 24.607 78.9455 24.687 79.217 ;
      RECT MASK 1 30.893 78.9455 30.973 79.217 ;
      RECT MASK 1 31.225 78.9455 31.305 79.217 ;
      RECT MASK 1 37.511 78.9455 37.591 79.217 ;
      RECT MASK 1 37.843 78.9455 37.923 79.217 ;
      RECT MASK 1 44.129 78.9455 44.209 79.217 ;
      RECT MASK 1 44.461 78.9455 44.541 79.217 ;
      RECT MASK 1 50.747 78.9455 50.827 79.217 ;
      RECT MASK 1 51.079 78.9455 51.159 79.217 ;
      RECT MASK 1 57.365 78.9455 57.445 79.217 ;
      RECT MASK 1 57.697 78.9455 57.777 79.217 ;
      RECT MASK 1 63.983 78.9455 64.063 79.217 ;
      RECT MASK 1 64.315 78.9455 64.395 79.217 ;
      RECT MASK 1 70.601 78.9455 70.681 79.217 ;
      RECT MASK 1 70.933 78.9455 71.013 79.217 ;
      RECT MASK 1 77.219 78.9455 77.299 79.217 ;
      RECT MASK 1 77.551 78.9455 77.631 79.217 ;
      RECT MASK 1 83.837 78.9455 83.917 79.217 ;
      RECT MASK 1 84.169 78.9455 84.249 79.217 ;
      RECT MASK 1 90.455 78.9455 90.535 79.217 ;
      RECT MASK 1 90.787 78.9455 90.867 79.217 ;
      RECT MASK 1 97.073 78.9455 97.153 79.217 ;
      RECT MASK 1 97.405 78.9455 97.485 79.217 ;
      RECT MASK 1 103.691 78.9455 103.771 79.217 ;
      RECT MASK 1 104.023 78.9455 104.103 79.217 ;
      RECT MASK 1 1.273 78.9635 1.353 95.9665 ;
      RECT MASK 1 5.257 78.9635 5.337 95.9665 ;
      RECT MASK 1 7.061 79.001 7.742 79.041 ;
      RECT MASK 1 8.223 79.001 8.904 79.041 ;
      RECT MASK 1 9.385 79.001 10.066 79.041 ;
      RECT MASK 1 12.517 79.001 13.198 79.041 ;
      RECT MASK 1 13.679 79.001 14.36 79.041 ;
      RECT MASK 1 14.841 79.001 15.522 79.041 ;
      RECT MASK 1 16.003 79.001 16.684 79.041 ;
      RECT MASK 1 19.135 79.001 19.816 79.041 ;
      RECT MASK 1 20.297 79.001 20.978 79.041 ;
      RECT MASK 1 21.459 79.001 22.14 79.041 ;
      RECT MASK 1 22.621 79.001 23.302 79.041 ;
      RECT MASK 1 25.753 79.001 26.434 79.041 ;
      RECT MASK 1 26.915 79.001 27.596 79.041 ;
      RECT MASK 1 28.077 79.001 28.758 79.041 ;
      RECT MASK 1 29.239 79.001 29.92 79.041 ;
      RECT MASK 1 32.371 79.001 33.052 79.041 ;
      RECT MASK 1 33.533 79.001 34.214 79.041 ;
      RECT MASK 1 34.695 79.001 35.376 79.041 ;
      RECT MASK 1 35.857 79.001 36.538 79.041 ;
      RECT MASK 1 38.989 79.001 39.67 79.041 ;
      RECT MASK 1 40.151 79.001 40.832 79.041 ;
      RECT MASK 1 41.313 79.001 41.994 79.041 ;
      RECT MASK 1 42.475 79.001 43.156 79.041 ;
      RECT MASK 1 45.607 79.001 46.288 79.041 ;
      RECT MASK 1 46.769 79.001 47.45 79.041 ;
      RECT MASK 1 47.931 79.001 48.612 79.041 ;
      RECT MASK 1 49.093 79.001 49.774 79.041 ;
      RECT MASK 1 52.225 79.001 52.906 79.041 ;
      RECT MASK 1 53.387 79.001 54.068 79.041 ;
      RECT MASK 1 54.549 79.001 55.23 79.041 ;
      RECT MASK 1 55.711 79.001 56.392 79.041 ;
      RECT MASK 1 58.843 79.001 59.524 79.041 ;
      RECT MASK 1 60.005 79.001 60.686 79.041 ;
      RECT MASK 1 61.167 79.001 61.848 79.041 ;
      RECT MASK 1 62.329 79.001 63.01 79.041 ;
      RECT MASK 1 65.461 79.001 66.142 79.041 ;
      RECT MASK 1 66.623 79.001 67.304 79.041 ;
      RECT MASK 1 67.785 79.001 68.466 79.041 ;
      RECT MASK 1 68.947 79.001 69.628 79.041 ;
      RECT MASK 1 72.079 79.001 72.76 79.041 ;
      RECT MASK 1 73.241 79.001 73.922 79.041 ;
      RECT MASK 1 74.403 79.001 75.084 79.041 ;
      RECT MASK 1 75.565 79.001 76.246 79.041 ;
      RECT MASK 1 78.697 79.001 79.378 79.041 ;
      RECT MASK 1 79.859 79.001 80.54 79.041 ;
      RECT MASK 1 81.021 79.001 81.702 79.041 ;
      RECT MASK 1 82.183 79.001 82.864 79.041 ;
      RECT MASK 1 85.315 79.001 85.996 79.041 ;
      RECT MASK 1 86.477 79.001 87.158 79.041 ;
      RECT MASK 1 87.639 79.001 88.32 79.041 ;
      RECT MASK 1 88.801 79.001 89.482 79.041 ;
      RECT MASK 1 91.933 79.001 92.614 79.041 ;
      RECT MASK 1 93.095 79.001 93.776 79.041 ;
      RECT MASK 1 94.257 79.001 94.938 79.041 ;
      RECT MASK 1 95.419 79.001 96.1 79.041 ;
      RECT MASK 1 98.551 79.001 99.232 79.041 ;
      RECT MASK 1 99.713 79.001 100.394 79.041 ;
      RECT MASK 1 100.875 79.001 101.556 79.041 ;
      RECT MASK 1 102.037 79.001 102.718 79.041 ;
      RECT MASK 1 105.169 79.001 105.85 79.041 ;
      RECT MASK 1 106.331 79.001 107.012 79.041 ;
      RECT MASK 1 107.493 79.001 108.174 79.041 ;
      RECT MASK 1 108.655 79.001 109.336 79.041 ;
      RECT MASK 1 116.339 79.012 126.654 79.052 ;
      RECT MASK 1 16.755 79.194 16.835 79.4645 ;
      RECT MASK 1 23.373 79.194 23.453 79.4645 ;
      RECT MASK 1 29.991 79.194 30.071 79.4645 ;
      RECT MASK 1 36.609 79.194 36.689 79.4645 ;
      RECT MASK 1 43.227 79.194 43.307 79.4645 ;
      RECT MASK 1 49.845 79.194 49.925 79.4645 ;
      RECT MASK 1 56.463 79.194 56.543 79.4645 ;
      RECT MASK 1 63.081 79.194 63.161 79.4645 ;
      RECT MASK 1 69.699 79.194 69.779 79.4645 ;
      RECT MASK 1 76.317 79.194 76.397 79.4645 ;
      RECT MASK 1 82.935 79.194 83.015 79.4645 ;
      RECT MASK 1 89.553 79.194 89.633 79.4645 ;
      RECT MASK 1 96.171 79.194 96.251 79.4645 ;
      RECT MASK 1 102.789 79.194 102.869 79.4645 ;
      RECT MASK 1 109.407 79.194 109.487 79.4645 ;
      RECT MASK 1 111.573 79.231 112.901 79.271 ;
      RECT MASK 1 6.983 79.2515 7.063 79.478 ;
      RECT MASK 1 7.315 79.2515 7.395 79.478 ;
      RECT MASK 1 8.145 79.2515 8.225 79.478 ;
      RECT MASK 1 8.477 79.2515 8.557 79.478 ;
      RECT MASK 1 9.307 79.2515 9.387 79.478 ;
      RECT MASK 1 9.639 79.2515 9.719 79.478 ;
      RECT MASK 1 12.439 79.2515 12.519 79.478 ;
      RECT MASK 1 12.771 79.2515 12.851 79.478 ;
      RECT MASK 1 13.601 79.2515 13.681 79.478 ;
      RECT MASK 1 13.933 79.2515 14.013 79.478 ;
      RECT MASK 1 14.763 79.2515 14.843 79.478 ;
      RECT MASK 1 15.095 79.2515 15.175 79.478 ;
      RECT MASK 1 15.925 79.2515 16.005 79.478 ;
      RECT MASK 1 16.257 79.2515 16.337 79.478 ;
      RECT MASK 1 19.057 79.2515 19.137 79.478 ;
      RECT MASK 1 19.389 79.2515 19.469 79.478 ;
      RECT MASK 1 20.219 79.2515 20.299 79.478 ;
      RECT MASK 1 20.551 79.2515 20.631 79.478 ;
      RECT MASK 1 21.381 79.2515 21.461 79.478 ;
      RECT MASK 1 21.713 79.2515 21.793 79.478 ;
      RECT MASK 1 22.543 79.2515 22.623 79.478 ;
      RECT MASK 1 22.875 79.2515 22.955 79.478 ;
      RECT MASK 1 25.675 79.2515 25.755 79.478 ;
      RECT MASK 1 26.007 79.2515 26.087 79.478 ;
      RECT MASK 1 26.837 79.2515 26.917 79.478 ;
      RECT MASK 1 27.169 79.2515 27.249 79.478 ;
      RECT MASK 1 27.999 79.2515 28.079 79.478 ;
      RECT MASK 1 28.331 79.2515 28.411 79.478 ;
      RECT MASK 1 29.161 79.2515 29.241 79.478 ;
      RECT MASK 1 29.493 79.2515 29.573 79.478 ;
      RECT MASK 1 32.293 79.2515 32.373 79.478 ;
      RECT MASK 1 32.625 79.2515 32.705 79.478 ;
      RECT MASK 1 33.455 79.2515 33.535 79.478 ;
      RECT MASK 1 33.787 79.2515 33.867 79.478 ;
      RECT MASK 1 34.617 79.2515 34.697 79.478 ;
      RECT MASK 1 34.949 79.2515 35.029 79.478 ;
      RECT MASK 1 35.779 79.2515 35.859 79.478 ;
      RECT MASK 1 36.111 79.2515 36.191 79.478 ;
      RECT MASK 1 38.911 79.2515 38.991 79.478 ;
      RECT MASK 1 39.243 79.2515 39.323 79.478 ;
      RECT MASK 1 40.073 79.2515 40.153 79.478 ;
      RECT MASK 1 40.405 79.2515 40.485 79.478 ;
      RECT MASK 1 41.235 79.2515 41.315 79.478 ;
      RECT MASK 1 41.567 79.2515 41.647 79.478 ;
      RECT MASK 1 42.397 79.2515 42.477 79.478 ;
      RECT MASK 1 42.729 79.2515 42.809 79.478 ;
      RECT MASK 1 45.529 79.2515 45.609 79.478 ;
      RECT MASK 1 45.861 79.2515 45.941 79.478 ;
      RECT MASK 1 46.691 79.2515 46.771 79.478 ;
      RECT MASK 1 47.023 79.2515 47.103 79.478 ;
      RECT MASK 1 47.853 79.2515 47.933 79.478 ;
      RECT MASK 1 48.185 79.2515 48.265 79.478 ;
      RECT MASK 1 49.015 79.2515 49.095 79.478 ;
      RECT MASK 1 49.347 79.2515 49.427 79.478 ;
      RECT MASK 1 52.147 79.2515 52.227 79.478 ;
      RECT MASK 1 52.479 79.2515 52.559 79.478 ;
      RECT MASK 1 53.309 79.2515 53.389 79.478 ;
      RECT MASK 1 53.641 79.2515 53.721 79.478 ;
      RECT MASK 1 54.471 79.2515 54.551 79.478 ;
      RECT MASK 1 54.803 79.2515 54.883 79.478 ;
      RECT MASK 1 55.633 79.2515 55.713 79.478 ;
      RECT MASK 1 55.965 79.2515 56.045 79.478 ;
      RECT MASK 1 58.765 79.2515 58.845 79.478 ;
      RECT MASK 1 59.097 79.2515 59.177 79.478 ;
      RECT MASK 1 59.927 79.2515 60.007 79.478 ;
      RECT MASK 1 60.259 79.2515 60.339 79.478 ;
      RECT MASK 1 61.089 79.2515 61.169 79.478 ;
      RECT MASK 1 61.421 79.2515 61.501 79.478 ;
      RECT MASK 1 62.251 79.2515 62.331 79.478 ;
      RECT MASK 1 62.583 79.2515 62.663 79.478 ;
      RECT MASK 1 65.383 79.2515 65.463 79.478 ;
      RECT MASK 1 65.715 79.2515 65.795 79.478 ;
      RECT MASK 1 66.545 79.2515 66.625 79.478 ;
      RECT MASK 1 66.877 79.2515 66.957 79.478 ;
      RECT MASK 1 67.707 79.2515 67.787 79.478 ;
      RECT MASK 1 68.039 79.2515 68.119 79.478 ;
      RECT MASK 1 68.869 79.2515 68.949 79.478 ;
      RECT MASK 1 69.201 79.2515 69.281 79.478 ;
      RECT MASK 1 72.001 79.2515 72.081 79.478 ;
      RECT MASK 1 72.333 79.2515 72.413 79.478 ;
      RECT MASK 1 73.163 79.2515 73.243 79.478 ;
      RECT MASK 1 73.495 79.2515 73.575 79.478 ;
      RECT MASK 1 74.325 79.2515 74.405 79.478 ;
      RECT MASK 1 74.657 79.2515 74.737 79.478 ;
      RECT MASK 1 75.487 79.2515 75.567 79.478 ;
      RECT MASK 1 75.819 79.2515 75.899 79.478 ;
      RECT MASK 1 78.619 79.2515 78.699 79.478 ;
      RECT MASK 1 78.951 79.2515 79.031 79.478 ;
      RECT MASK 1 79.781 79.2515 79.861 79.478 ;
      RECT MASK 1 80.113 79.2515 80.193 79.478 ;
      RECT MASK 1 80.943 79.2515 81.023 79.478 ;
      RECT MASK 1 81.275 79.2515 81.355 79.478 ;
      RECT MASK 1 82.105 79.2515 82.185 79.478 ;
      RECT MASK 1 82.437 79.2515 82.517 79.478 ;
      RECT MASK 1 85.237 79.2515 85.317 79.478 ;
      RECT MASK 1 85.569 79.2515 85.649 79.478 ;
      RECT MASK 1 86.399 79.2515 86.479 79.478 ;
      RECT MASK 1 86.731 79.2515 86.811 79.478 ;
      RECT MASK 1 87.561 79.2515 87.641 79.478 ;
      RECT MASK 1 87.893 79.2515 87.973 79.478 ;
      RECT MASK 1 88.723 79.2515 88.803 79.478 ;
      RECT MASK 1 89.055 79.2515 89.135 79.478 ;
      RECT MASK 1 91.855 79.2515 91.935 79.478 ;
      RECT MASK 1 92.187 79.2515 92.267 79.478 ;
      RECT MASK 1 93.017 79.2515 93.097 79.478 ;
      RECT MASK 1 93.349 79.2515 93.429 79.478 ;
      RECT MASK 1 94.179 79.2515 94.259 79.478 ;
      RECT MASK 1 94.511 79.2515 94.591 79.478 ;
      RECT MASK 1 95.341 79.2515 95.421 79.478 ;
      RECT MASK 1 95.673 79.2515 95.753 79.478 ;
      RECT MASK 1 98.473 79.2515 98.553 79.478 ;
      RECT MASK 1 98.805 79.2515 98.885 79.478 ;
      RECT MASK 1 99.635 79.2515 99.715 79.478 ;
      RECT MASK 1 99.967 79.2515 100.047 79.478 ;
      RECT MASK 1 100.797 79.2515 100.877 79.478 ;
      RECT MASK 1 101.129 79.2515 101.209 79.478 ;
      RECT MASK 1 101.959 79.2515 102.039 79.478 ;
      RECT MASK 1 102.291 79.2515 102.371 79.478 ;
      RECT MASK 1 105.091 79.2515 105.171 79.478 ;
      RECT MASK 1 105.423 79.2515 105.503 79.478 ;
      RECT MASK 1 106.253 79.2515 106.333 79.478 ;
      RECT MASK 1 106.585 79.2515 106.665 79.478 ;
      RECT MASK 1 107.415 79.2515 107.495 79.478 ;
      RECT MASK 1 107.747 79.2515 107.827 79.478 ;
      RECT MASK 1 108.577 79.2515 108.657 79.478 ;
      RECT MASK 1 108.909 79.2515 108.989 79.478 ;
      RECT MASK 1 2.067 79.26 2.127 80.31 ;
      RECT MASK 1 2.341 79.26 2.401 80.31 ;
      RECT MASK 1 2.615 79.26 2.675 80.31 ;
      RECT MASK 1 2.889 79.26 2.949 80.31 ;
      RECT MASK 1 3.163 79.26 3.223 80.31 ;
      RECT MASK 1 3.437 79.26 3.497 80.31 ;
      RECT MASK 1 3.711 79.26 3.771 80.31 ;
      RECT MASK 1 3.985 79.26 4.045 80.31 ;
      RECT MASK 1 4.259 79.26 4.319 80.31 ;
      RECT MASK 1 4.533 79.26 4.593 80.31 ;
      RECT MASK 1 111.122 79.415 113.352 79.455 ;
      RECT MASK 1 116.271 79.448 116.331 79.672 ;
      RECT MASK 1 116.603 79.448 116.663 79.672 ;
      RECT MASK 1 116.935 79.448 116.995 79.672 ;
      RECT MASK 1 117.267 79.448 117.327 79.672 ;
      RECT MASK 1 117.599 79.448 117.659 79.672 ;
      RECT MASK 1 117.931 79.448 117.991 79.672 ;
      RECT MASK 1 118.263 79.448 118.323 79.672 ;
      RECT MASK 1 118.595 79.448 118.655 79.672 ;
      RECT MASK 1 118.927 79.448 118.987 79.672 ;
      RECT MASK 1 119.259 79.448 119.319 79.672 ;
      RECT MASK 1 119.591 79.448 119.651 79.672 ;
      RECT MASK 1 119.923 79.448 119.983 79.672 ;
      RECT MASK 1 120.255 79.448 120.315 79.672 ;
      RECT MASK 1 120.587 79.448 120.647 79.672 ;
      RECT MASK 1 120.919 79.448 120.979 79.672 ;
      RECT MASK 1 121.251 79.448 121.311 79.672 ;
      RECT MASK 1 121.583 79.448 121.643 79.672 ;
      RECT MASK 1 121.915 79.448 121.975 79.672 ;
      RECT MASK 1 122.247 79.448 122.307 79.672 ;
      RECT MASK 1 122.579 79.448 122.639 79.672 ;
      RECT MASK 1 122.911 79.448 122.971 79.672 ;
      RECT MASK 1 123.243 79.448 123.303 79.672 ;
      RECT MASK 1 123.575 79.448 123.635 79.672 ;
      RECT MASK 1 123.907 79.448 123.967 79.672 ;
      RECT MASK 1 124.239 79.448 124.299 79.672 ;
      RECT MASK 1 124.571 79.448 124.631 79.672 ;
      RECT MASK 1 124.903 79.448 124.963 79.672 ;
      RECT MASK 1 125.235 79.448 125.295 79.672 ;
      RECT MASK 1 125.567 79.448 125.627 79.672 ;
      RECT MASK 1 125.899 79.448 125.959 79.672 ;
      RECT MASK 1 126.231 79.448 126.291 79.672 ;
      RECT MASK 1 111.767 79.599 111.95 79.639 ;
      RECT MASK 1 112.431 79.599 112.614 79.639 ;
      RECT MASK 1 6.691 79.676 10.315 79.716 ;
      RECT MASK 1 12.009 79.676 16.933 79.716 ;
      RECT MASK 1 18.627 79.676 23.551 79.716 ;
      RECT MASK 1 25.245 79.676 30.169 79.716 ;
      RECT MASK 1 31.863 79.676 36.787 79.716 ;
      RECT MASK 1 38.481 79.676 43.405 79.716 ;
      RECT MASK 1 45.099 79.676 50.023 79.716 ;
      RECT MASK 1 51.717 79.676 56.641 79.716 ;
      RECT MASK 1 58.335 79.676 63.259 79.716 ;
      RECT MASK 1 64.953 79.676 69.877 79.716 ;
      RECT MASK 1 71.571 79.676 76.495 79.716 ;
      RECT MASK 1 78.189 79.676 83.113 79.716 ;
      RECT MASK 1 84.807 79.676 89.731 79.716 ;
      RECT MASK 1 91.425 79.676 96.349 79.716 ;
      RECT MASK 1 98.043 79.676 102.967 79.716 ;
      RECT MASK 1 104.661 79.676 109.585 79.716 ;
      RECT MASK 1 111.767 79.767 111.95 79.807 ;
      RECT MASK 1 112.431 79.767 112.614 79.807 ;
      RECT MASK 1 116.339 79.792 126.649 79.832 ;
      RECT MASK 1 111.151 79.821 111.331 79.861 ;
      RECT MASK 1 113.143 79.821 113.323 79.861 ;
      RECT MASK 1 111.151 79.989 111.331 80.029 ;
      RECT MASK 1 111.732 79.989 112.078 80.029 ;
      RECT MASK 1 112.396 79.989 112.742 80.029 ;
      RECT MASK 1 113.143 79.989 113.323 80.029 ;
      RECT MASK 1 6.2775 80.095 110.065 80.135 ;
      RECT MASK 1 111.113 80.211 113.361 80.251 ;
      RECT MASK 1 115.539 80.275 126.947 80.315 ;
      RECT MASK 1 6.2775 80.545 109.836 80.585 ;
      RECT MASK 1 6.319 80.82 6.399 82.238 ;
      RECT MASK 1 10.469 80.82 10.549 82.238 ;
      RECT MASK 1 11.775 80.82 11.855 82.238 ;
      RECT MASK 1 17.087 80.82 17.167 82.238 ;
      RECT MASK 1 18.393 80.82 18.473 82.238 ;
      RECT MASK 1 23.705 80.82 23.785 82.238 ;
      RECT MASK 1 25.011 80.82 25.091 82.238 ;
      RECT MASK 1 30.323 80.82 30.403 82.238 ;
      RECT MASK 1 31.629 80.82 31.709 82.238 ;
      RECT MASK 1 36.941 80.82 37.021 82.238 ;
      RECT MASK 1 38.247 80.82 38.327 82.238 ;
      RECT MASK 1 43.559 80.82 43.639 82.238 ;
      RECT MASK 1 44.865 80.82 44.945 82.238 ;
      RECT MASK 1 50.177 80.82 50.257 82.238 ;
      RECT MASK 1 51.483 80.82 51.563 82.238 ;
      RECT MASK 1 56.795 80.82 56.875 82.238 ;
      RECT MASK 1 58.101 80.82 58.181 82.238 ;
      RECT MASK 1 63.413 80.82 63.493 82.238 ;
      RECT MASK 1 64.719 80.82 64.799 82.238 ;
      RECT MASK 1 70.031 80.82 70.111 82.238 ;
      RECT MASK 1 71.337 80.82 71.417 82.238 ;
      RECT MASK 1 76.649 80.82 76.729 82.238 ;
      RECT MASK 1 77.955 80.82 78.035 82.238 ;
      RECT MASK 1 83.267 80.82 83.347 82.238 ;
      RECT MASK 1 84.573 80.82 84.653 82.238 ;
      RECT MASK 1 89.885 80.82 89.965 82.238 ;
      RECT MASK 1 91.191 80.82 91.271 82.238 ;
      RECT MASK 1 96.503 80.82 96.583 82.238 ;
      RECT MASK 1 97.809 80.82 97.889 82.238 ;
      RECT MASK 1 103.121 80.82 103.201 82.238 ;
      RECT MASK 1 104.427 80.82 104.507 82.238 ;
      RECT MASK 1 109.739 80.82 109.819 82.238 ;
      RECT MASK 1 111.075 80.939 113.399 80.979 ;
      RECT MASK 1 2.067 80.97 2.127 82.02 ;
      RECT MASK 1 2.341 80.97 2.401 82.02 ;
      RECT MASK 1 2.615 80.97 2.675 82.02 ;
      RECT MASK 1 2.889 80.97 2.949 82.02 ;
      RECT MASK 1 3.163 80.97 3.223 82.02 ;
      RECT MASK 1 3.437 80.97 3.497 82.02 ;
      RECT MASK 1 3.711 80.97 3.771 82.02 ;
      RECT MASK 1 3.985 80.97 4.045 82.02 ;
      RECT MASK 1 4.259 80.97 4.319 82.02 ;
      RECT MASK 1 4.533 80.97 4.593 82.02 ;
      RECT MASK 1 6.983 80.986 7.063 81.211 ;
      RECT MASK 1 7.315 80.986 7.395 81.211 ;
      RECT MASK 1 8.145 80.986 8.225 81.211 ;
      RECT MASK 1 8.477 80.986 8.557 81.211 ;
      RECT MASK 1 9.307 80.986 9.387 81.211 ;
      RECT MASK 1 9.639 80.986 9.719 81.211 ;
      RECT MASK 1 12.439 80.986 12.519 81.211 ;
      RECT MASK 1 12.771 80.986 12.851 81.211 ;
      RECT MASK 1 13.601 80.986 13.681 81.211 ;
      RECT MASK 1 13.933 80.986 14.013 81.211 ;
      RECT MASK 1 14.763 80.986 14.843 81.211 ;
      RECT MASK 1 15.095 80.986 15.175 81.211 ;
      RECT MASK 1 15.925 80.986 16.005 81.211 ;
      RECT MASK 1 16.257 80.986 16.337 81.211 ;
      RECT MASK 1 19.057 80.986 19.137 81.211 ;
      RECT MASK 1 19.389 80.986 19.469 81.211 ;
      RECT MASK 1 20.219 80.986 20.299 81.211 ;
      RECT MASK 1 20.551 80.986 20.631 81.211 ;
      RECT MASK 1 21.381 80.986 21.461 81.211 ;
      RECT MASK 1 21.713 80.986 21.793 81.211 ;
      RECT MASK 1 22.543 80.986 22.623 81.211 ;
      RECT MASK 1 22.875 80.986 22.955 81.211 ;
      RECT MASK 1 25.675 80.986 25.755 81.211 ;
      RECT MASK 1 26.007 80.986 26.087 81.211 ;
      RECT MASK 1 26.837 80.986 26.917 81.211 ;
      RECT MASK 1 27.169 80.986 27.249 81.211 ;
      RECT MASK 1 27.999 80.986 28.079 81.211 ;
      RECT MASK 1 28.331 80.986 28.411 81.211 ;
      RECT MASK 1 29.161 80.986 29.241 81.211 ;
      RECT MASK 1 29.493 80.986 29.573 81.211 ;
      RECT MASK 1 32.293 80.986 32.373 81.211 ;
      RECT MASK 1 32.625 80.986 32.705 81.211 ;
      RECT MASK 1 33.455 80.986 33.535 81.211 ;
      RECT MASK 1 33.787 80.986 33.867 81.211 ;
      RECT MASK 1 34.617 80.986 34.697 81.211 ;
      RECT MASK 1 34.949 80.986 35.029 81.211 ;
      RECT MASK 1 35.779 80.986 35.859 81.211 ;
      RECT MASK 1 36.111 80.986 36.191 81.211 ;
      RECT MASK 1 38.911 80.986 38.991 81.211 ;
      RECT MASK 1 39.243 80.986 39.323 81.211 ;
      RECT MASK 1 40.073 80.986 40.153 81.211 ;
      RECT MASK 1 40.405 80.986 40.485 81.211 ;
      RECT MASK 1 41.235 80.986 41.315 81.211 ;
      RECT MASK 1 41.567 80.986 41.647 81.211 ;
      RECT MASK 1 42.397 80.986 42.477 81.211 ;
      RECT MASK 1 42.729 80.986 42.809 81.211 ;
      RECT MASK 1 45.529 80.986 45.609 81.211 ;
      RECT MASK 1 45.861 80.986 45.941 81.211 ;
      RECT MASK 1 46.691 80.986 46.771 81.211 ;
      RECT MASK 1 47.023 80.986 47.103 81.211 ;
      RECT MASK 1 47.853 80.986 47.933 81.211 ;
      RECT MASK 1 48.185 80.986 48.265 81.211 ;
      RECT MASK 1 49.015 80.986 49.095 81.211 ;
      RECT MASK 1 49.347 80.986 49.427 81.211 ;
      RECT MASK 1 52.147 80.986 52.227 81.211 ;
      RECT MASK 1 52.479 80.986 52.559 81.211 ;
      RECT MASK 1 53.309 80.986 53.389 81.211 ;
      RECT MASK 1 53.641 80.986 53.721 81.211 ;
      RECT MASK 1 54.471 80.986 54.551 81.211 ;
      RECT MASK 1 54.803 80.986 54.883 81.211 ;
      RECT MASK 1 55.633 80.986 55.713 81.211 ;
      RECT MASK 1 55.965 80.986 56.045 81.211 ;
      RECT MASK 1 58.765 80.986 58.845 81.211 ;
      RECT MASK 1 59.097 80.986 59.177 81.211 ;
      RECT MASK 1 59.927 80.986 60.007 81.211 ;
      RECT MASK 1 60.259 80.986 60.339 81.211 ;
      RECT MASK 1 61.089 80.986 61.169 81.211 ;
      RECT MASK 1 61.421 80.986 61.501 81.211 ;
      RECT MASK 1 62.251 80.986 62.331 81.211 ;
      RECT MASK 1 62.583 80.986 62.663 81.211 ;
      RECT MASK 1 65.383 80.986 65.463 81.211 ;
      RECT MASK 1 65.715 80.986 65.795 81.211 ;
      RECT MASK 1 66.545 80.986 66.625 81.211 ;
      RECT MASK 1 66.877 80.986 66.957 81.211 ;
      RECT MASK 1 67.707 80.986 67.787 81.211 ;
      RECT MASK 1 68.039 80.986 68.119 81.211 ;
      RECT MASK 1 68.869 80.986 68.949 81.211 ;
      RECT MASK 1 69.201 80.986 69.281 81.211 ;
      RECT MASK 1 72.001 80.986 72.081 81.211 ;
      RECT MASK 1 72.333 80.986 72.413 81.211 ;
      RECT MASK 1 73.163 80.986 73.243 81.211 ;
      RECT MASK 1 73.495 80.986 73.575 81.211 ;
      RECT MASK 1 74.325 80.986 74.405 81.211 ;
      RECT MASK 1 74.657 80.986 74.737 81.211 ;
      RECT MASK 1 75.487 80.986 75.567 81.211 ;
      RECT MASK 1 75.819 80.986 75.899 81.211 ;
      RECT MASK 1 78.619 80.986 78.699 81.211 ;
      RECT MASK 1 78.951 80.986 79.031 81.211 ;
      RECT MASK 1 79.781 80.986 79.861 81.211 ;
      RECT MASK 1 80.113 80.986 80.193 81.211 ;
      RECT MASK 1 80.943 80.986 81.023 81.211 ;
      RECT MASK 1 81.275 80.986 81.355 81.211 ;
      RECT MASK 1 82.105 80.986 82.185 81.211 ;
      RECT MASK 1 82.437 80.986 82.517 81.211 ;
      RECT MASK 1 85.237 80.986 85.317 81.211 ;
      RECT MASK 1 85.569 80.986 85.649 81.211 ;
      RECT MASK 1 86.399 80.986 86.479 81.211 ;
      RECT MASK 1 86.731 80.986 86.811 81.211 ;
      RECT MASK 1 87.561 80.986 87.641 81.211 ;
      RECT MASK 1 87.893 80.986 87.973 81.211 ;
      RECT MASK 1 88.723 80.986 88.803 81.211 ;
      RECT MASK 1 89.055 80.986 89.135 81.211 ;
      RECT MASK 1 91.855 80.986 91.935 81.211 ;
      RECT MASK 1 92.187 80.986 92.267 81.211 ;
      RECT MASK 1 93.017 80.986 93.097 81.211 ;
      RECT MASK 1 93.349 80.986 93.429 81.211 ;
      RECT MASK 1 94.179 80.986 94.259 81.211 ;
      RECT MASK 1 94.511 80.986 94.591 81.211 ;
      RECT MASK 1 95.341 80.986 95.421 81.211 ;
      RECT MASK 1 95.673 80.986 95.753 81.211 ;
      RECT MASK 1 98.473 80.986 98.553 81.211 ;
      RECT MASK 1 98.805 80.986 98.885 81.211 ;
      RECT MASK 1 99.635 80.986 99.715 81.211 ;
      RECT MASK 1 99.967 80.986 100.047 81.211 ;
      RECT MASK 1 100.797 80.986 100.877 81.211 ;
      RECT MASK 1 101.129 80.986 101.209 81.211 ;
      RECT MASK 1 101.959 80.986 102.039 81.211 ;
      RECT MASK 1 102.291 80.986 102.371 81.211 ;
      RECT MASK 1 105.091 80.986 105.171 81.211 ;
      RECT MASK 1 105.423 80.986 105.503 81.211 ;
      RECT MASK 1 106.253 80.986 106.333 81.211 ;
      RECT MASK 1 106.585 80.986 106.665 81.211 ;
      RECT MASK 1 107.415 80.986 107.495 81.211 ;
      RECT MASK 1 107.747 80.986 107.827 81.211 ;
      RECT MASK 1 108.577 80.986 108.657 81.211 ;
      RECT MASK 1 108.909 80.986 108.989 81.211 ;
      RECT MASK 1 111.732 81.161 112.078 81.201 ;
      RECT MASK 1 112.396 81.161 112.742 81.201 ;
      RECT MASK 1 111.151 81.197 111.331 81.237 ;
      RECT MASK 1 113.143 81.197 113.323 81.237 ;
      RECT MASK 1 111.151 81.365 111.331 81.405 ;
      RECT MASK 1 113.143 81.365 113.323 81.405 ;
      RECT MASK 1 111.86 81.383 112.043 81.423 ;
      RECT MASK 1 112.524 81.383 112.707 81.423 ;
      RECT MASK 1 6.691 81.4 10.315 81.44 ;
      RECT MASK 1 12.009 81.4 16.933 81.44 ;
      RECT MASK 1 18.627 81.4 23.551 81.44 ;
      RECT MASK 1 25.245 81.4 30.169 81.44 ;
      RECT MASK 1 31.863 81.4 36.787 81.44 ;
      RECT MASK 1 38.481 81.4 43.405 81.44 ;
      RECT MASK 1 45.099 81.4 50.023 81.44 ;
      RECT MASK 1 51.717 81.4 56.641 81.44 ;
      RECT MASK 1 58.473 81.4 63.259 81.44 ;
      RECT MASK 1 64.953 81.4 69.877 81.44 ;
      RECT MASK 1 71.571 81.4 76.495 81.44 ;
      RECT MASK 1 78.189 81.4 83.113 81.44 ;
      RECT MASK 1 84.807 81.4 89.731 81.44 ;
      RECT MASK 1 91.425 81.4 96.349 81.44 ;
      RECT MASK 1 98.043 81.4 102.967 81.44 ;
      RECT MASK 1 104.661 81.4 109.585 81.44 ;
      RECT MASK 1 115.613 81.445 128.525 81.485 ;
      RECT MASK 1 11.039 81.463 11.119 81.7345 ;
      RECT MASK 1 11.371 81.463 11.451 81.7345 ;
      RECT MASK 1 17.657 81.463 17.737 81.7345 ;
      RECT MASK 1 17.989 81.463 18.069 81.7345 ;
      RECT MASK 1 24.275 81.463 24.355 81.7345 ;
      RECT MASK 1 24.607 81.463 24.687 81.7345 ;
      RECT MASK 1 30.893 81.463 30.973 81.7345 ;
      RECT MASK 1 31.225 81.463 31.305 81.7345 ;
      RECT MASK 1 37.511 81.463 37.591 81.7345 ;
      RECT MASK 1 37.843 81.463 37.923 81.7345 ;
      RECT MASK 1 44.129 81.463 44.209 81.7345 ;
      RECT MASK 1 44.461 81.463 44.541 81.7345 ;
      RECT MASK 1 50.747 81.463 50.827 81.7345 ;
      RECT MASK 1 51.079 81.463 51.159 81.7345 ;
      RECT MASK 1 57.365 81.463 57.445 81.7345 ;
      RECT MASK 1 57.697 81.463 57.777 81.7345 ;
      RECT MASK 1 63.983 81.463 64.063 81.7345 ;
      RECT MASK 1 64.315 81.463 64.395 81.7345 ;
      RECT MASK 1 70.601 81.463 70.681 81.7345 ;
      RECT MASK 1 70.933 81.463 71.013 81.7345 ;
      RECT MASK 1 77.219 81.463 77.299 81.7345 ;
      RECT MASK 1 77.551 81.463 77.631 81.7345 ;
      RECT MASK 1 83.837 81.463 83.917 81.7345 ;
      RECT MASK 1 84.169 81.463 84.249 81.7345 ;
      RECT MASK 1 90.455 81.463 90.535 81.7345 ;
      RECT MASK 1 90.787 81.463 90.867 81.7345 ;
      RECT MASK 1 97.073 81.463 97.153 81.7345 ;
      RECT MASK 1 97.405 81.463 97.485 81.7345 ;
      RECT MASK 1 103.691 81.463 103.771 81.7345 ;
      RECT MASK 1 104.023 81.463 104.103 81.7345 ;
      RECT MASK 1 111.86 81.551 112.043 81.591 ;
      RECT MASK 1 112.524 81.551 112.707 81.591 ;
      RECT MASK 1 6.983 81.6515 7.063 81.882 ;
      RECT MASK 1 7.315 81.6515 7.395 81.882 ;
      RECT MASK 1 8.145 81.6515 8.225 81.882 ;
      RECT MASK 1 8.477 81.6515 8.557 81.882 ;
      RECT MASK 1 9.307 81.6515 9.387 81.882 ;
      RECT MASK 1 9.639 81.6515 9.719 81.882 ;
      RECT MASK 1 12.439 81.6515 12.519 81.882 ;
      RECT MASK 1 12.771 81.6515 12.851 81.882 ;
      RECT MASK 1 13.601 81.6515 13.681 81.882 ;
      RECT MASK 1 13.933 81.6515 14.013 81.882 ;
      RECT MASK 1 14.763 81.6515 14.843 81.882 ;
      RECT MASK 1 15.095 81.6515 15.175 81.882 ;
      RECT MASK 1 15.925 81.6515 16.005 81.882 ;
      RECT MASK 1 16.257 81.6515 16.337 81.882 ;
      RECT MASK 1 19.057 81.6515 19.137 81.882 ;
      RECT MASK 1 19.389 81.6515 19.469 81.882 ;
      RECT MASK 1 20.219 81.6515 20.299 81.882 ;
      RECT MASK 1 20.551 81.6515 20.631 81.882 ;
      RECT MASK 1 21.381 81.6515 21.461 81.882 ;
      RECT MASK 1 21.713 81.6515 21.793 81.882 ;
      RECT MASK 1 22.543 81.6515 22.623 81.882 ;
      RECT MASK 1 22.875 81.6515 22.955 81.882 ;
      RECT MASK 1 25.675 81.6515 25.755 81.882 ;
      RECT MASK 1 26.007 81.6515 26.087 81.882 ;
      RECT MASK 1 26.837 81.6515 26.917 81.882 ;
      RECT MASK 1 27.169 81.6515 27.249 81.882 ;
      RECT MASK 1 27.999 81.6515 28.079 81.882 ;
      RECT MASK 1 28.331 81.6515 28.411 81.882 ;
      RECT MASK 1 29.161 81.6515 29.241 81.882 ;
      RECT MASK 1 29.493 81.6515 29.573 81.882 ;
      RECT MASK 1 32.293 81.6515 32.373 81.882 ;
      RECT MASK 1 32.625 81.6515 32.705 81.882 ;
      RECT MASK 1 33.455 81.6515 33.535 81.882 ;
      RECT MASK 1 33.787 81.6515 33.867 81.882 ;
      RECT MASK 1 34.617 81.6515 34.697 81.882 ;
      RECT MASK 1 34.949 81.6515 35.029 81.882 ;
      RECT MASK 1 35.779 81.6515 35.859 81.882 ;
      RECT MASK 1 36.111 81.6515 36.191 81.882 ;
      RECT MASK 1 38.911 81.6515 38.991 81.882 ;
      RECT MASK 1 39.243 81.6515 39.323 81.882 ;
      RECT MASK 1 40.073 81.6515 40.153 81.882 ;
      RECT MASK 1 40.405 81.6515 40.485 81.882 ;
      RECT MASK 1 41.235 81.6515 41.315 81.882 ;
      RECT MASK 1 41.567 81.6515 41.647 81.882 ;
      RECT MASK 1 42.397 81.6515 42.477 81.882 ;
      RECT MASK 1 42.729 81.6515 42.809 81.882 ;
      RECT MASK 1 45.529 81.6515 45.609 81.882 ;
      RECT MASK 1 45.861 81.6515 45.941 81.882 ;
      RECT MASK 1 46.691 81.6515 46.771 81.882 ;
      RECT MASK 1 47.023 81.6515 47.103 81.882 ;
      RECT MASK 1 47.853 81.6515 47.933 81.882 ;
      RECT MASK 1 48.185 81.6515 48.265 81.882 ;
      RECT MASK 1 49.015 81.6515 49.095 81.882 ;
      RECT MASK 1 49.347 81.6515 49.427 81.882 ;
      RECT MASK 1 52.147 81.6515 52.227 81.882 ;
      RECT MASK 1 52.479 81.6515 52.559 81.882 ;
      RECT MASK 1 53.309 81.6515 53.389 81.882 ;
      RECT MASK 1 53.641 81.6515 53.721 81.882 ;
      RECT MASK 1 54.471 81.6515 54.551 81.882 ;
      RECT MASK 1 54.803 81.6515 54.883 81.882 ;
      RECT MASK 1 55.633 81.6515 55.713 81.882 ;
      RECT MASK 1 55.965 81.6515 56.045 81.882 ;
      RECT MASK 1 58.765 81.6515 58.845 81.882 ;
      RECT MASK 1 59.097 81.6515 59.177 81.882 ;
      RECT MASK 1 59.927 81.6515 60.007 81.882 ;
      RECT MASK 1 60.259 81.6515 60.339 81.882 ;
      RECT MASK 1 61.089 81.6515 61.169 81.882 ;
      RECT MASK 1 61.421 81.6515 61.501 81.882 ;
      RECT MASK 1 62.251 81.6515 62.331 81.882 ;
      RECT MASK 1 62.583 81.6515 62.663 81.882 ;
      RECT MASK 1 65.383 81.6515 65.463 81.882 ;
      RECT MASK 1 65.715 81.6515 65.795 81.882 ;
      RECT MASK 1 66.545 81.6515 66.625 81.882 ;
      RECT MASK 1 66.877 81.6515 66.957 81.882 ;
      RECT MASK 1 67.707 81.6515 67.787 81.882 ;
      RECT MASK 1 68.039 81.6515 68.119 81.882 ;
      RECT MASK 1 68.869 81.6515 68.949 81.882 ;
      RECT MASK 1 69.201 81.6515 69.281 81.882 ;
      RECT MASK 1 72.001 81.6515 72.081 81.882 ;
      RECT MASK 1 72.333 81.6515 72.413 81.882 ;
      RECT MASK 1 73.163 81.6515 73.243 81.882 ;
      RECT MASK 1 73.495 81.6515 73.575 81.882 ;
      RECT MASK 1 74.325 81.6515 74.405 81.882 ;
      RECT MASK 1 74.657 81.6515 74.737 81.882 ;
      RECT MASK 1 75.487 81.6515 75.567 81.882 ;
      RECT MASK 1 75.819 81.6515 75.899 81.882 ;
      RECT MASK 1 78.619 81.6515 78.699 81.882 ;
      RECT MASK 1 78.951 81.6515 79.031 81.882 ;
      RECT MASK 1 79.781 81.6515 79.861 81.882 ;
      RECT MASK 1 80.113 81.6515 80.193 81.882 ;
      RECT MASK 1 80.943 81.6515 81.023 81.882 ;
      RECT MASK 1 81.275 81.6515 81.355 81.882 ;
      RECT MASK 1 82.105 81.6515 82.185 81.882 ;
      RECT MASK 1 82.437 81.6515 82.517 81.882 ;
      RECT MASK 1 85.237 81.6515 85.317 81.882 ;
      RECT MASK 1 85.569 81.6515 85.649 81.882 ;
      RECT MASK 1 86.399 81.6515 86.479 81.882 ;
      RECT MASK 1 86.731 81.6515 86.811 81.882 ;
      RECT MASK 1 87.561 81.6515 87.641 81.882 ;
      RECT MASK 1 87.893 81.6515 87.973 81.882 ;
      RECT MASK 1 88.723 81.6515 88.803 81.882 ;
      RECT MASK 1 89.055 81.6515 89.135 81.882 ;
      RECT MASK 1 91.855 81.6515 91.935 81.882 ;
      RECT MASK 1 92.187 81.6515 92.267 81.882 ;
      RECT MASK 1 93.017 81.6515 93.097 81.882 ;
      RECT MASK 1 93.349 81.6515 93.429 81.882 ;
      RECT MASK 1 94.179 81.6515 94.259 81.882 ;
      RECT MASK 1 94.511 81.6515 94.591 81.882 ;
      RECT MASK 1 95.341 81.6515 95.421 81.882 ;
      RECT MASK 1 95.673 81.6515 95.753 81.882 ;
      RECT MASK 1 98.473 81.6515 98.553 81.882 ;
      RECT MASK 1 98.805 81.6515 98.885 81.882 ;
      RECT MASK 1 99.635 81.6515 99.715 81.882 ;
      RECT MASK 1 99.967 81.6515 100.047 81.882 ;
      RECT MASK 1 100.797 81.6515 100.877 81.882 ;
      RECT MASK 1 101.129 81.6515 101.209 81.882 ;
      RECT MASK 1 101.959 81.6515 102.039 81.882 ;
      RECT MASK 1 102.291 81.6515 102.371 81.882 ;
      RECT MASK 1 105.091 81.6515 105.171 81.882 ;
      RECT MASK 1 105.423 81.6515 105.503 81.882 ;
      RECT MASK 1 106.253 81.6515 106.333 81.882 ;
      RECT MASK 1 106.585 81.6515 106.665 81.882 ;
      RECT MASK 1 107.415 81.6515 107.495 81.882 ;
      RECT MASK 1 107.747 81.6515 107.827 81.882 ;
      RECT MASK 1 108.577 81.6515 108.657 81.882 ;
      RECT MASK 1 108.909 81.6515 108.989 81.882 ;
      RECT MASK 1 111.151 81.735 113.323 81.775 ;
      RECT MASK 1 115.638 81.7535 115.718 86.6365 ;
      RECT MASK 1 128.42 81.7535 128.5 86.6365 ;
      RECT MASK 1 111.573 81.919 112.901 81.959 ;
      RECT MASK 1 116.462 82.05 116.522 83.1 ;
      RECT MASK 1 116.736 82.05 116.796 83.1 ;
      RECT MASK 1 117.01 82.05 117.07 83.1 ;
      RECT MASK 1 117.284 82.05 117.344 83.1 ;
      RECT MASK 1 117.558 82.05 117.618 83.1 ;
      RECT MASK 1 117.832 82.05 117.892 83.1 ;
      RECT MASK 1 118.106 82.05 118.166 83.1 ;
      RECT MASK 1 118.38 82.05 118.44 83.1 ;
      RECT MASK 1 118.654 82.05 118.714 83.1 ;
      RECT MASK 1 118.928 82.05 118.988 83.1 ;
      RECT MASK 1 119.202 82.05 119.262 83.1 ;
      RECT MASK 1 119.476 82.05 119.536 83.1 ;
      RECT MASK 1 119.75 82.05 119.81 83.1 ;
      RECT MASK 1 120.024 82.05 120.084 83.1 ;
      RECT MASK 1 120.298 82.05 120.358 83.1 ;
      RECT MASK 1 120.572 82.05 120.632 83.1 ;
      RECT MASK 1 120.846 82.05 120.906 83.1 ;
      RECT MASK 1 121.12 82.05 121.18 83.1 ;
      RECT MASK 1 121.394 82.05 121.454 83.1 ;
      RECT MASK 1 121.668 82.05 121.728 83.1 ;
      RECT MASK 1 121.942 82.05 122.002 83.1 ;
      RECT MASK 1 122.216 82.05 122.276 83.1 ;
      RECT MASK 1 122.49 82.05 122.55 83.1 ;
      RECT MASK 1 122.764 82.05 122.824 83.1 ;
      RECT MASK 1 123.038 82.05 123.098 83.1 ;
      RECT MASK 1 123.312 82.05 123.372 83.1 ;
      RECT MASK 1 123.586 82.05 123.646 83.1 ;
      RECT MASK 1 123.86 82.05 123.92 83.1 ;
      RECT MASK 1 124.134 82.05 124.194 83.1 ;
      RECT MASK 1 124.408 82.05 124.468 83.1 ;
      RECT MASK 1 124.682 82.05 124.742 83.1 ;
      RECT MASK 1 124.956 82.05 125.016 83.1 ;
      RECT MASK 1 125.23 82.05 125.29 83.1 ;
      RECT MASK 1 125.504 82.05 125.564 83.1 ;
      RECT MASK 1 125.778 82.05 125.838 83.1 ;
      RECT MASK 1 126.052 82.05 126.112 83.1 ;
      RECT MASK 1 126.326 82.05 126.386 83.1 ;
      RECT MASK 1 126.6 82.05 126.66 83.1 ;
      RECT MASK 1 126.874 82.05 126.934 83.1 ;
      RECT MASK 1 127.148 82.05 127.208 83.1 ;
      RECT MASK 1 127.422 82.05 127.482 83.1 ;
      RECT MASK 1 127.696 82.05 127.756 83.1 ;
      RECT MASK 1 7.0505 82.066 7.327 82.106 ;
      RECT MASK 1 8.2125 82.066 8.489 82.106 ;
      RECT MASK 1 9.3745 82.066 9.651 82.106 ;
      RECT MASK 1 12.5065 82.066 12.783 82.106 ;
      RECT MASK 1 13.6685 82.066 13.945 82.106 ;
      RECT MASK 1 14.8305 82.066 15.107 82.106 ;
      RECT MASK 1 15.9925 82.066 16.269 82.106 ;
      RECT MASK 1 19.1245 82.066 19.401 82.106 ;
      RECT MASK 1 20.2865 82.066 20.563 82.106 ;
      RECT MASK 1 21.4485 82.066 21.725 82.106 ;
      RECT MASK 1 22.6105 82.066 22.887 82.106 ;
      RECT MASK 1 25.7425 82.066 26.019 82.106 ;
      RECT MASK 1 26.9045 82.066 27.181 82.106 ;
      RECT MASK 1 28.0665 82.066 28.343 82.106 ;
      RECT MASK 1 29.2285 82.066 29.505 82.106 ;
      RECT MASK 1 32.3605 82.066 32.637 82.106 ;
      RECT MASK 1 33.5225 82.066 33.799 82.106 ;
      RECT MASK 1 34.6845 82.066 34.961 82.106 ;
      RECT MASK 1 35.8465 82.066 36.123 82.106 ;
      RECT MASK 1 38.9785 82.066 39.255 82.106 ;
      RECT MASK 1 40.1405 82.066 40.417 82.106 ;
      RECT MASK 1 41.3025 82.066 41.579 82.106 ;
      RECT MASK 1 42.4645 82.066 42.741 82.106 ;
      RECT MASK 1 45.5965 82.066 45.873 82.106 ;
      RECT MASK 1 46.7585 82.066 47.035 82.106 ;
      RECT MASK 1 47.9205 82.066 48.197 82.106 ;
      RECT MASK 1 49.0825 82.066 49.359 82.106 ;
      RECT MASK 1 52.2145 82.066 52.491 82.106 ;
      RECT MASK 1 53.3765 82.066 53.653 82.106 ;
      RECT MASK 1 54.5385 82.066 54.815 82.106 ;
      RECT MASK 1 55.7005 82.066 55.977 82.106 ;
      RECT MASK 1 58.8325 82.066 59.109 82.106 ;
      RECT MASK 1 59.9945 82.066 60.271 82.106 ;
      RECT MASK 1 61.1565 82.066 61.433 82.106 ;
      RECT MASK 1 62.3185 82.066 62.595 82.106 ;
      RECT MASK 1 65.4505 82.066 65.727 82.106 ;
      RECT MASK 1 66.6125 82.066 66.889 82.106 ;
      RECT MASK 1 67.7745 82.066 68.051 82.106 ;
      RECT MASK 1 68.9365 82.066 69.213 82.106 ;
      RECT MASK 1 72.0685 82.066 72.345 82.106 ;
      RECT MASK 1 73.2305 82.066 73.507 82.106 ;
      RECT MASK 1 74.3925 82.066 74.669 82.106 ;
      RECT MASK 1 75.5545 82.066 75.831 82.106 ;
      RECT MASK 1 78.6865 82.066 78.963 82.106 ;
      RECT MASK 1 79.8485 82.066 80.125 82.106 ;
      RECT MASK 1 81.0105 82.066 81.287 82.106 ;
      RECT MASK 1 82.1725 82.066 82.449 82.106 ;
      RECT MASK 1 85.3045 82.066 85.581 82.106 ;
      RECT MASK 1 86.4665 82.066 86.743 82.106 ;
      RECT MASK 1 87.6285 82.066 87.905 82.106 ;
      RECT MASK 1 88.7905 82.066 89.067 82.106 ;
      RECT MASK 1 91.9225 82.066 92.199 82.106 ;
      RECT MASK 1 93.0845 82.066 93.361 82.106 ;
      RECT MASK 1 94.2465 82.066 94.523 82.106 ;
      RECT MASK 1 95.4085 82.066 95.685 82.106 ;
      RECT MASK 1 98.5405 82.066 98.817 82.106 ;
      RECT MASK 1 99.7025 82.066 99.979 82.106 ;
      RECT MASK 1 100.8645 82.066 101.141 82.106 ;
      RECT MASK 1 102.0265 82.066 102.303 82.106 ;
      RECT MASK 1 105.1585 82.066 105.435 82.106 ;
      RECT MASK 1 106.3205 82.066 106.597 82.106 ;
      RECT MASK 1 107.4825 82.066 107.759 82.106 ;
      RECT MASK 1 108.6445 82.066 108.921 82.106 ;
      RECT MASK 1 111.186 82.255 113.288 82.295 ;
      RECT MASK 1 6.2775 82.495 109.836 82.535 ;
      RECT MASK 1 2.067 82.68 2.127 83.73 ;
      RECT MASK 1 2.341 82.68 2.401 83.73 ;
      RECT MASK 1 2.615 82.68 2.675 83.73 ;
      RECT MASK 1 2.889 82.68 2.949 83.73 ;
      RECT MASK 1 3.163 82.68 3.223 83.73 ;
      RECT MASK 1 3.437 82.68 3.497 83.73 ;
      RECT MASK 1 3.711 82.68 3.771 83.73 ;
      RECT MASK 1 3.985 82.68 4.045 83.73 ;
      RECT MASK 1 4.259 82.68 4.319 83.73 ;
      RECT MASK 1 4.533 82.68 4.593 83.73 ;
      RECT MASK 1 6.2775 82.861 109.836 82.901 ;
      RECT MASK 1 6.269 83.045 109.869 83.085 ;
      RECT MASK 1 6.978 83.229 7.161 83.269 ;
      RECT MASK 1 7.383 83.229 7.566 83.269 ;
      RECT MASK 1 8.14 83.229 8.323 83.269 ;
      RECT MASK 1 8.545 83.229 8.728 83.269 ;
      RECT MASK 1 9.302 83.229 9.485 83.269 ;
      RECT MASK 1 9.707 83.229 9.89 83.269 ;
      RECT MASK 1 12.434 83.229 12.617 83.269 ;
      RECT MASK 1 12.839 83.229 13.022 83.269 ;
      RECT MASK 1 13.596 83.229 13.779 83.269 ;
      RECT MASK 1 14.001 83.229 14.184 83.269 ;
      RECT MASK 1 14.758 83.229 14.941 83.269 ;
      RECT MASK 1 15.163 83.229 15.346 83.269 ;
      RECT MASK 1 15.92 83.229 16.103 83.269 ;
      RECT MASK 1 16.325 83.229 16.508 83.269 ;
      RECT MASK 1 19.052 83.229 19.235 83.269 ;
      RECT MASK 1 19.457 83.229 19.64 83.269 ;
      RECT MASK 1 20.214 83.229 20.397 83.269 ;
      RECT MASK 1 20.619 83.229 20.802 83.269 ;
      RECT MASK 1 21.376 83.229 21.559 83.269 ;
      RECT MASK 1 21.781 83.229 21.964 83.269 ;
      RECT MASK 1 22.538 83.229 22.721 83.269 ;
      RECT MASK 1 22.943 83.229 23.126 83.269 ;
      RECT MASK 1 25.67 83.229 25.853 83.269 ;
      RECT MASK 1 26.075 83.229 26.258 83.269 ;
      RECT MASK 1 26.832 83.229 27.015 83.269 ;
      RECT MASK 1 27.237 83.229 27.42 83.269 ;
      RECT MASK 1 27.994 83.229 28.177 83.269 ;
      RECT MASK 1 28.399 83.229 28.582 83.269 ;
      RECT MASK 1 29.156 83.229 29.339 83.269 ;
      RECT MASK 1 29.561 83.229 29.744 83.269 ;
      RECT MASK 1 32.288 83.229 32.471 83.269 ;
      RECT MASK 1 32.693 83.229 32.876 83.269 ;
      RECT MASK 1 33.45 83.229 33.633 83.269 ;
      RECT MASK 1 33.855 83.229 34.038 83.269 ;
      RECT MASK 1 34.612 83.229 34.795 83.269 ;
      RECT MASK 1 35.017 83.229 35.2 83.269 ;
      RECT MASK 1 35.774 83.229 35.957 83.269 ;
      RECT MASK 1 36.179 83.229 36.362 83.269 ;
      RECT MASK 1 38.906 83.229 39.089 83.269 ;
      RECT MASK 1 39.311 83.229 39.494 83.269 ;
      RECT MASK 1 40.068 83.229 40.251 83.269 ;
      RECT MASK 1 40.473 83.229 40.656 83.269 ;
      RECT MASK 1 41.23 83.229 41.413 83.269 ;
      RECT MASK 1 41.635 83.229 41.818 83.269 ;
      RECT MASK 1 42.392 83.229 42.575 83.269 ;
      RECT MASK 1 42.797 83.229 42.98 83.269 ;
      RECT MASK 1 45.524 83.229 45.707 83.269 ;
      RECT MASK 1 45.929 83.229 46.112 83.269 ;
      RECT MASK 1 46.686 83.229 46.869 83.269 ;
      RECT MASK 1 47.091 83.229 47.274 83.269 ;
      RECT MASK 1 47.848 83.229 48.031 83.269 ;
      RECT MASK 1 48.253 83.229 48.436 83.269 ;
      RECT MASK 1 49.01 83.229 49.193 83.269 ;
      RECT MASK 1 49.415 83.229 49.598 83.269 ;
      RECT MASK 1 52.142 83.229 52.325 83.269 ;
      RECT MASK 1 52.547 83.229 52.73 83.269 ;
      RECT MASK 1 53.304 83.229 53.487 83.269 ;
      RECT MASK 1 53.709 83.229 53.892 83.269 ;
      RECT MASK 1 54.466 83.229 54.649 83.269 ;
      RECT MASK 1 54.871 83.229 55.054 83.269 ;
      RECT MASK 1 55.628 83.229 55.811 83.269 ;
      RECT MASK 1 56.033 83.229 56.216 83.269 ;
      RECT MASK 1 58.76 83.229 58.943 83.269 ;
      RECT MASK 1 59.165 83.229 59.348 83.269 ;
      RECT MASK 1 59.922 83.229 60.105 83.269 ;
      RECT MASK 1 60.327 83.229 60.51 83.269 ;
      RECT MASK 1 61.084 83.229 61.267 83.269 ;
      RECT MASK 1 61.489 83.229 61.672 83.269 ;
      RECT MASK 1 62.246 83.229 62.429 83.269 ;
      RECT MASK 1 62.651 83.229 62.834 83.269 ;
      RECT MASK 1 65.378 83.229 65.561 83.269 ;
      RECT MASK 1 65.783 83.229 65.966 83.269 ;
      RECT MASK 1 66.54 83.229 66.723 83.269 ;
      RECT MASK 1 66.945 83.229 67.128 83.269 ;
      RECT MASK 1 67.702 83.229 67.885 83.269 ;
      RECT MASK 1 68.107 83.229 68.29 83.269 ;
      RECT MASK 1 68.864 83.229 69.047 83.269 ;
      RECT MASK 1 69.269 83.229 69.452 83.269 ;
      RECT MASK 1 71.996 83.229 72.179 83.269 ;
      RECT MASK 1 72.401 83.229 72.584 83.269 ;
      RECT MASK 1 73.158 83.229 73.341 83.269 ;
      RECT MASK 1 73.563 83.229 73.746 83.269 ;
      RECT MASK 1 74.32 83.229 74.503 83.269 ;
      RECT MASK 1 74.725 83.229 74.908 83.269 ;
      RECT MASK 1 75.482 83.229 75.665 83.269 ;
      RECT MASK 1 75.887 83.229 76.07 83.269 ;
      RECT MASK 1 78.614 83.229 78.797 83.269 ;
      RECT MASK 1 79.019 83.229 79.202 83.269 ;
      RECT MASK 1 79.776 83.229 79.959 83.269 ;
      RECT MASK 1 80.181 83.229 80.364 83.269 ;
      RECT MASK 1 80.938 83.229 81.121 83.269 ;
      RECT MASK 1 81.343 83.229 81.526 83.269 ;
      RECT MASK 1 82.1 83.229 82.283 83.269 ;
      RECT MASK 1 82.505 83.229 82.688 83.269 ;
      RECT MASK 1 85.232 83.229 85.415 83.269 ;
      RECT MASK 1 85.637 83.229 85.82 83.269 ;
      RECT MASK 1 86.394 83.229 86.577 83.269 ;
      RECT MASK 1 86.799 83.229 86.982 83.269 ;
      RECT MASK 1 87.556 83.229 87.739 83.269 ;
      RECT MASK 1 87.961 83.229 88.144 83.269 ;
      RECT MASK 1 88.718 83.229 88.901 83.269 ;
      RECT MASK 1 89.123 83.229 89.306 83.269 ;
      RECT MASK 1 91.85 83.229 92.033 83.269 ;
      RECT MASK 1 92.255 83.229 92.438 83.269 ;
      RECT MASK 1 93.012 83.229 93.195 83.269 ;
      RECT MASK 1 93.417 83.229 93.6 83.269 ;
      RECT MASK 1 94.174 83.229 94.357 83.269 ;
      RECT MASK 1 94.579 83.229 94.762 83.269 ;
      RECT MASK 1 95.336 83.229 95.519 83.269 ;
      RECT MASK 1 95.741 83.229 95.924 83.269 ;
      RECT MASK 1 98.468 83.229 98.651 83.269 ;
      RECT MASK 1 98.873 83.229 99.056 83.269 ;
      RECT MASK 1 99.63 83.229 99.813 83.269 ;
      RECT MASK 1 100.035 83.229 100.218 83.269 ;
      RECT MASK 1 100.792 83.229 100.975 83.269 ;
      RECT MASK 1 101.197 83.229 101.38 83.269 ;
      RECT MASK 1 101.954 83.229 102.137 83.269 ;
      RECT MASK 1 102.359 83.229 102.542 83.269 ;
      RECT MASK 1 105.086 83.229 105.269 83.269 ;
      RECT MASK 1 105.491 83.229 105.674 83.269 ;
      RECT MASK 1 106.248 83.229 106.431 83.269 ;
      RECT MASK 1 106.653 83.229 106.836 83.269 ;
      RECT MASK 1 107.41 83.229 107.593 83.269 ;
      RECT MASK 1 107.815 83.229 107.998 83.269 ;
      RECT MASK 1 108.572 83.229 108.755 83.269 ;
      RECT MASK 1 108.977 83.229 109.16 83.269 ;
      RECT MASK 1 6.978 83.397 7.161 83.437 ;
      RECT MASK 1 7.383 83.397 7.566 83.437 ;
      RECT MASK 1 8.14 83.397 8.323 83.437 ;
      RECT MASK 1 8.545 83.397 8.728 83.437 ;
      RECT MASK 1 9.302 83.397 9.485 83.437 ;
      RECT MASK 1 9.707 83.397 9.89 83.437 ;
      RECT MASK 1 12.434 83.397 12.617 83.437 ;
      RECT MASK 1 12.839 83.397 13.022 83.437 ;
      RECT MASK 1 13.596 83.397 13.779 83.437 ;
      RECT MASK 1 14.001 83.397 14.184 83.437 ;
      RECT MASK 1 14.758 83.397 14.941 83.437 ;
      RECT MASK 1 15.163 83.397 15.346 83.437 ;
      RECT MASK 1 15.92 83.397 16.103 83.437 ;
      RECT MASK 1 16.325 83.397 16.508 83.437 ;
      RECT MASK 1 19.052 83.397 19.235 83.437 ;
      RECT MASK 1 19.457 83.397 19.64 83.437 ;
      RECT MASK 1 20.214 83.397 20.397 83.437 ;
      RECT MASK 1 20.619 83.397 20.802 83.437 ;
      RECT MASK 1 21.376 83.397 21.559 83.437 ;
      RECT MASK 1 21.781 83.397 21.964 83.437 ;
      RECT MASK 1 22.538 83.397 22.721 83.437 ;
      RECT MASK 1 22.943 83.397 23.126 83.437 ;
      RECT MASK 1 25.67 83.397 25.853 83.437 ;
      RECT MASK 1 26.075 83.397 26.258 83.437 ;
      RECT MASK 1 26.832 83.397 27.015 83.437 ;
      RECT MASK 1 27.237 83.397 27.42 83.437 ;
      RECT MASK 1 27.994 83.397 28.177 83.437 ;
      RECT MASK 1 28.399 83.397 28.582 83.437 ;
      RECT MASK 1 29.156 83.397 29.339 83.437 ;
      RECT MASK 1 29.561 83.397 29.744 83.437 ;
      RECT MASK 1 32.288 83.397 32.471 83.437 ;
      RECT MASK 1 32.693 83.397 32.876 83.437 ;
      RECT MASK 1 33.45 83.397 33.633 83.437 ;
      RECT MASK 1 33.855 83.397 34.038 83.437 ;
      RECT MASK 1 34.612 83.397 34.795 83.437 ;
      RECT MASK 1 35.017 83.397 35.2 83.437 ;
      RECT MASK 1 35.774 83.397 35.957 83.437 ;
      RECT MASK 1 36.179 83.397 36.362 83.437 ;
      RECT MASK 1 38.906 83.397 39.089 83.437 ;
      RECT MASK 1 39.311 83.397 39.494 83.437 ;
      RECT MASK 1 40.068 83.397 40.251 83.437 ;
      RECT MASK 1 40.473 83.397 40.656 83.437 ;
      RECT MASK 1 41.23 83.397 41.413 83.437 ;
      RECT MASK 1 41.635 83.397 41.818 83.437 ;
      RECT MASK 1 42.392 83.397 42.575 83.437 ;
      RECT MASK 1 42.797 83.397 42.98 83.437 ;
      RECT MASK 1 45.524 83.397 45.707 83.437 ;
      RECT MASK 1 45.929 83.397 46.112 83.437 ;
      RECT MASK 1 46.686 83.397 46.869 83.437 ;
      RECT MASK 1 47.091 83.397 47.274 83.437 ;
      RECT MASK 1 47.848 83.397 48.031 83.437 ;
      RECT MASK 1 48.253 83.397 48.436 83.437 ;
      RECT MASK 1 49.01 83.397 49.193 83.437 ;
      RECT MASK 1 49.415 83.397 49.598 83.437 ;
      RECT MASK 1 52.142 83.397 52.325 83.437 ;
      RECT MASK 1 52.547 83.397 52.73 83.437 ;
      RECT MASK 1 53.304 83.397 53.487 83.437 ;
      RECT MASK 1 53.709 83.397 53.892 83.437 ;
      RECT MASK 1 54.466 83.397 54.649 83.437 ;
      RECT MASK 1 54.871 83.397 55.054 83.437 ;
      RECT MASK 1 55.628 83.397 55.811 83.437 ;
      RECT MASK 1 56.033 83.397 56.216 83.437 ;
      RECT MASK 1 58.76 83.397 58.943 83.437 ;
      RECT MASK 1 59.165 83.397 59.348 83.437 ;
      RECT MASK 1 59.922 83.397 60.105 83.437 ;
      RECT MASK 1 60.327 83.397 60.51 83.437 ;
      RECT MASK 1 61.084 83.397 61.267 83.437 ;
      RECT MASK 1 61.489 83.397 61.672 83.437 ;
      RECT MASK 1 62.246 83.397 62.429 83.437 ;
      RECT MASK 1 62.651 83.397 62.834 83.437 ;
      RECT MASK 1 65.378 83.397 65.561 83.437 ;
      RECT MASK 1 65.783 83.397 65.966 83.437 ;
      RECT MASK 1 66.54 83.397 66.723 83.437 ;
      RECT MASK 1 66.945 83.397 67.128 83.437 ;
      RECT MASK 1 67.702 83.397 67.885 83.437 ;
      RECT MASK 1 68.107 83.397 68.29 83.437 ;
      RECT MASK 1 68.864 83.397 69.047 83.437 ;
      RECT MASK 1 69.269 83.397 69.452 83.437 ;
      RECT MASK 1 71.996 83.397 72.179 83.437 ;
      RECT MASK 1 72.401 83.397 72.584 83.437 ;
      RECT MASK 1 73.158 83.397 73.341 83.437 ;
      RECT MASK 1 73.563 83.397 73.746 83.437 ;
      RECT MASK 1 74.32 83.397 74.503 83.437 ;
      RECT MASK 1 74.725 83.397 74.908 83.437 ;
      RECT MASK 1 75.482 83.397 75.665 83.437 ;
      RECT MASK 1 75.887 83.397 76.07 83.437 ;
      RECT MASK 1 78.614 83.397 78.797 83.437 ;
      RECT MASK 1 79.019 83.397 79.202 83.437 ;
      RECT MASK 1 79.776 83.397 79.959 83.437 ;
      RECT MASK 1 80.181 83.397 80.364 83.437 ;
      RECT MASK 1 80.938 83.397 81.121 83.437 ;
      RECT MASK 1 81.343 83.397 81.526 83.437 ;
      RECT MASK 1 82.1 83.397 82.283 83.437 ;
      RECT MASK 1 82.505 83.397 82.688 83.437 ;
      RECT MASK 1 85.232 83.397 85.415 83.437 ;
      RECT MASK 1 85.637 83.397 85.82 83.437 ;
      RECT MASK 1 86.394 83.397 86.577 83.437 ;
      RECT MASK 1 86.799 83.397 86.982 83.437 ;
      RECT MASK 1 87.556 83.397 87.739 83.437 ;
      RECT MASK 1 87.961 83.397 88.144 83.437 ;
      RECT MASK 1 88.718 83.397 88.901 83.437 ;
      RECT MASK 1 89.123 83.397 89.306 83.437 ;
      RECT MASK 1 91.85 83.397 92.033 83.437 ;
      RECT MASK 1 92.255 83.397 92.438 83.437 ;
      RECT MASK 1 93.012 83.397 93.195 83.437 ;
      RECT MASK 1 93.417 83.397 93.6 83.437 ;
      RECT MASK 1 94.174 83.397 94.357 83.437 ;
      RECT MASK 1 94.579 83.397 94.762 83.437 ;
      RECT MASK 1 95.336 83.397 95.519 83.437 ;
      RECT MASK 1 95.741 83.397 95.924 83.437 ;
      RECT MASK 1 98.468 83.397 98.651 83.437 ;
      RECT MASK 1 98.873 83.397 99.056 83.437 ;
      RECT MASK 1 99.63 83.397 99.813 83.437 ;
      RECT MASK 1 100.035 83.397 100.218 83.437 ;
      RECT MASK 1 100.792 83.397 100.975 83.437 ;
      RECT MASK 1 101.197 83.397 101.38 83.437 ;
      RECT MASK 1 101.954 83.397 102.137 83.437 ;
      RECT MASK 1 102.359 83.397 102.542 83.437 ;
      RECT MASK 1 105.086 83.397 105.269 83.437 ;
      RECT MASK 1 105.491 83.397 105.674 83.437 ;
      RECT MASK 1 106.248 83.397 106.431 83.437 ;
      RECT MASK 1 106.653 83.397 106.836 83.437 ;
      RECT MASK 1 107.41 83.397 107.593 83.437 ;
      RECT MASK 1 107.815 83.397 107.998 83.437 ;
      RECT MASK 1 108.572 83.397 108.755 83.437 ;
      RECT MASK 1 108.977 83.397 109.16 83.437 ;
      RECT MASK 1 6.269 83.415 6.449 83.455 ;
      RECT MASK 1 10.419 83.415 10.599 83.455 ;
      RECT MASK 1 11.725 83.415 11.905 83.455 ;
      RECT MASK 1 17.037 83.415 17.217 83.455 ;
      RECT MASK 1 18.343 83.415 18.523 83.455 ;
      RECT MASK 1 23.655 83.415 23.835 83.455 ;
      RECT MASK 1 24.961 83.415 25.141 83.455 ;
      RECT MASK 1 30.273 83.415 30.453 83.455 ;
      RECT MASK 1 31.579 83.415 31.759 83.455 ;
      RECT MASK 1 36.891 83.415 37.071 83.455 ;
      RECT MASK 1 38.197 83.415 38.377 83.455 ;
      RECT MASK 1 43.509 83.415 43.689 83.455 ;
      RECT MASK 1 44.815 83.415 44.995 83.455 ;
      RECT MASK 1 50.127 83.415 50.307 83.455 ;
      RECT MASK 1 51.433 83.415 51.613 83.455 ;
      RECT MASK 1 56.745 83.415 56.925 83.455 ;
      RECT MASK 1 58.051 83.415 58.231 83.455 ;
      RECT MASK 1 63.363 83.415 63.543 83.455 ;
      RECT MASK 1 64.669 83.415 64.849 83.455 ;
      RECT MASK 1 69.981 83.415 70.161 83.455 ;
      RECT MASK 1 71.287 83.415 71.467 83.455 ;
      RECT MASK 1 76.599 83.415 76.779 83.455 ;
      RECT MASK 1 77.905 83.415 78.085 83.455 ;
      RECT MASK 1 83.217 83.415 83.397 83.455 ;
      RECT MASK 1 84.523 83.415 84.703 83.455 ;
      RECT MASK 1 89.835 83.415 90.015 83.455 ;
      RECT MASK 1 91.141 83.415 91.321 83.455 ;
      RECT MASK 1 96.453 83.415 96.633 83.455 ;
      RECT MASK 1 97.759 83.415 97.939 83.455 ;
      RECT MASK 1 103.071 83.415 103.251 83.455 ;
      RECT MASK 1 104.377 83.415 104.557 83.455 ;
      RECT MASK 1 109.689 83.415 109.869 83.455 ;
      RECT MASK 1 6.269 83.583 6.449 83.623 ;
      RECT MASK 1 10.419 83.583 10.599 83.623 ;
      RECT MASK 1 11.725 83.583 11.905 83.623 ;
      RECT MASK 1 17.037 83.583 17.217 83.623 ;
      RECT MASK 1 18.343 83.583 18.523 83.623 ;
      RECT MASK 1 23.655 83.583 23.835 83.623 ;
      RECT MASK 1 24.961 83.583 25.141 83.623 ;
      RECT MASK 1 30.273 83.583 30.453 83.623 ;
      RECT MASK 1 31.579 83.583 31.759 83.623 ;
      RECT MASK 1 36.891 83.583 37.071 83.623 ;
      RECT MASK 1 38.197 83.583 38.377 83.623 ;
      RECT MASK 1 43.509 83.583 43.689 83.623 ;
      RECT MASK 1 44.815 83.583 44.995 83.623 ;
      RECT MASK 1 50.127 83.583 50.307 83.623 ;
      RECT MASK 1 51.433 83.583 51.613 83.623 ;
      RECT MASK 1 56.745 83.583 56.925 83.623 ;
      RECT MASK 1 58.051 83.583 58.231 83.623 ;
      RECT MASK 1 63.363 83.583 63.543 83.623 ;
      RECT MASK 1 64.669 83.583 64.849 83.623 ;
      RECT MASK 1 69.981 83.583 70.161 83.623 ;
      RECT MASK 1 71.287 83.583 71.467 83.623 ;
      RECT MASK 1 76.599 83.583 76.779 83.623 ;
      RECT MASK 1 77.905 83.583 78.085 83.623 ;
      RECT MASK 1 83.217 83.583 83.397 83.623 ;
      RECT MASK 1 84.523 83.583 84.703 83.623 ;
      RECT MASK 1 89.835 83.583 90.015 83.623 ;
      RECT MASK 1 91.141 83.583 91.321 83.623 ;
      RECT MASK 1 96.453 83.583 96.633 83.623 ;
      RECT MASK 1 97.759 83.583 97.939 83.623 ;
      RECT MASK 1 103.071 83.583 103.251 83.623 ;
      RECT MASK 1 104.377 83.583 104.557 83.623 ;
      RECT MASK 1 109.689 83.583 109.869 83.623 ;
      RECT MASK 1 6.85 83.619 7.03 83.659 ;
      RECT MASK 1 7.514 83.619 7.694 83.659 ;
      RECT MASK 1 8.012 83.619 8.192 83.659 ;
      RECT MASK 1 8.676 83.619 8.856 83.659 ;
      RECT MASK 1 9.174 83.619 9.354 83.659 ;
      RECT MASK 1 9.838 83.619 10.018 83.659 ;
      RECT MASK 1 12.306 83.619 12.486 83.659 ;
      RECT MASK 1 12.97 83.619 13.15 83.659 ;
      RECT MASK 1 13.468 83.619 13.648 83.659 ;
      RECT MASK 1 14.132 83.619 14.312 83.659 ;
      RECT MASK 1 14.63 83.619 14.81 83.659 ;
      RECT MASK 1 15.294 83.619 15.474 83.659 ;
      RECT MASK 1 15.792 83.619 15.972 83.659 ;
      RECT MASK 1 16.456 83.619 16.636 83.659 ;
      RECT MASK 1 18.924 83.619 19.104 83.659 ;
      RECT MASK 1 19.588 83.619 19.768 83.659 ;
      RECT MASK 1 20.086 83.619 20.266 83.659 ;
      RECT MASK 1 20.75 83.619 20.93 83.659 ;
      RECT MASK 1 21.248 83.619 21.428 83.659 ;
      RECT MASK 1 21.912 83.619 22.092 83.659 ;
      RECT MASK 1 22.41 83.619 22.59 83.659 ;
      RECT MASK 1 23.074 83.619 23.254 83.659 ;
      RECT MASK 1 25.542 83.619 25.722 83.659 ;
      RECT MASK 1 26.206 83.619 26.386 83.659 ;
      RECT MASK 1 26.704 83.619 26.884 83.659 ;
      RECT MASK 1 27.368 83.619 27.548 83.659 ;
      RECT MASK 1 27.866 83.619 28.046 83.659 ;
      RECT MASK 1 28.53 83.619 28.71 83.659 ;
      RECT MASK 1 29.028 83.619 29.208 83.659 ;
      RECT MASK 1 29.692 83.619 29.872 83.659 ;
      RECT MASK 1 32.16 83.619 32.34 83.659 ;
      RECT MASK 1 32.824 83.619 33.004 83.659 ;
      RECT MASK 1 33.322 83.619 33.502 83.659 ;
      RECT MASK 1 33.986 83.619 34.166 83.659 ;
      RECT MASK 1 34.484 83.619 34.664 83.659 ;
      RECT MASK 1 35.148 83.619 35.328 83.659 ;
      RECT MASK 1 35.646 83.619 35.826 83.659 ;
      RECT MASK 1 36.31 83.619 36.49 83.659 ;
      RECT MASK 1 38.778 83.619 38.958 83.659 ;
      RECT MASK 1 39.442 83.619 39.622 83.659 ;
      RECT MASK 1 39.94 83.619 40.12 83.659 ;
      RECT MASK 1 40.604 83.619 40.784 83.659 ;
      RECT MASK 1 41.102 83.619 41.282 83.659 ;
      RECT MASK 1 41.766 83.619 41.946 83.659 ;
      RECT MASK 1 42.264 83.619 42.444 83.659 ;
      RECT MASK 1 42.928 83.619 43.108 83.659 ;
      RECT MASK 1 45.396 83.619 45.576 83.659 ;
      RECT MASK 1 46.06 83.619 46.24 83.659 ;
      RECT MASK 1 46.558 83.619 46.738 83.659 ;
      RECT MASK 1 47.222 83.619 47.402 83.659 ;
      RECT MASK 1 47.72 83.619 47.9 83.659 ;
      RECT MASK 1 48.384 83.619 48.564 83.659 ;
      RECT MASK 1 48.882 83.619 49.062 83.659 ;
      RECT MASK 1 49.546 83.619 49.726 83.659 ;
      RECT MASK 1 52.014 83.619 52.194 83.659 ;
      RECT MASK 1 52.678 83.619 52.858 83.659 ;
      RECT MASK 1 53.176 83.619 53.356 83.659 ;
      RECT MASK 1 53.84 83.619 54.02 83.659 ;
      RECT MASK 1 54.338 83.619 54.518 83.659 ;
      RECT MASK 1 55.002 83.619 55.182 83.659 ;
      RECT MASK 1 55.5 83.619 55.68 83.659 ;
      RECT MASK 1 56.164 83.619 56.344 83.659 ;
      RECT MASK 1 58.632 83.619 58.812 83.659 ;
      RECT MASK 1 59.296 83.619 59.476 83.659 ;
      RECT MASK 1 59.794 83.619 59.974 83.659 ;
      RECT MASK 1 60.458 83.619 60.638 83.659 ;
      RECT MASK 1 60.956 83.619 61.136 83.659 ;
      RECT MASK 1 61.62 83.619 61.8 83.659 ;
      RECT MASK 1 62.118 83.619 62.298 83.659 ;
      RECT MASK 1 62.782 83.619 62.962 83.659 ;
      RECT MASK 1 65.25 83.619 65.43 83.659 ;
      RECT MASK 1 65.914 83.619 66.094 83.659 ;
      RECT MASK 1 66.412 83.619 66.592 83.659 ;
      RECT MASK 1 67.076 83.619 67.256 83.659 ;
      RECT MASK 1 67.574 83.619 67.754 83.659 ;
      RECT MASK 1 68.238 83.619 68.418 83.659 ;
      RECT MASK 1 68.736 83.619 68.916 83.659 ;
      RECT MASK 1 69.4 83.619 69.58 83.659 ;
      RECT MASK 1 71.868 83.619 72.048 83.659 ;
      RECT MASK 1 72.532 83.619 72.712 83.659 ;
      RECT MASK 1 73.03 83.619 73.21 83.659 ;
      RECT MASK 1 73.694 83.619 73.874 83.659 ;
      RECT MASK 1 74.192 83.619 74.372 83.659 ;
      RECT MASK 1 74.856 83.619 75.036 83.659 ;
      RECT MASK 1 75.354 83.619 75.534 83.659 ;
      RECT MASK 1 76.018 83.619 76.198 83.659 ;
      RECT MASK 1 78.486 83.619 78.666 83.659 ;
      RECT MASK 1 79.15 83.619 79.33 83.659 ;
      RECT MASK 1 79.648 83.619 79.828 83.659 ;
      RECT MASK 1 80.312 83.619 80.492 83.659 ;
      RECT MASK 1 80.81 83.619 80.99 83.659 ;
      RECT MASK 1 81.474 83.619 81.654 83.659 ;
      RECT MASK 1 81.972 83.619 82.152 83.659 ;
      RECT MASK 1 82.636 83.619 82.816 83.659 ;
      RECT MASK 1 85.104 83.619 85.284 83.659 ;
      RECT MASK 1 85.768 83.619 85.948 83.659 ;
      RECT MASK 1 86.266 83.619 86.446 83.659 ;
      RECT MASK 1 86.93 83.619 87.11 83.659 ;
      RECT MASK 1 87.428 83.619 87.608 83.659 ;
      RECT MASK 1 88.092 83.619 88.272 83.659 ;
      RECT MASK 1 88.59 83.619 88.77 83.659 ;
      RECT MASK 1 89.254 83.619 89.434 83.659 ;
      RECT MASK 1 91.722 83.619 91.902 83.659 ;
      RECT MASK 1 92.386 83.619 92.566 83.659 ;
      RECT MASK 1 92.884 83.619 93.064 83.659 ;
      RECT MASK 1 93.548 83.619 93.728 83.659 ;
      RECT MASK 1 94.046 83.619 94.226 83.659 ;
      RECT MASK 1 94.71 83.619 94.89 83.659 ;
      RECT MASK 1 95.208 83.619 95.388 83.659 ;
      RECT MASK 1 95.872 83.619 96.052 83.659 ;
      RECT MASK 1 98.34 83.619 98.52 83.659 ;
      RECT MASK 1 99.004 83.619 99.184 83.659 ;
      RECT MASK 1 99.502 83.619 99.682 83.659 ;
      RECT MASK 1 100.166 83.619 100.346 83.659 ;
      RECT MASK 1 100.664 83.619 100.844 83.659 ;
      RECT MASK 1 101.328 83.619 101.508 83.659 ;
      RECT MASK 1 101.826 83.619 102.006 83.659 ;
      RECT MASK 1 102.49 83.619 102.67 83.659 ;
      RECT MASK 1 104.958 83.619 105.138 83.659 ;
      RECT MASK 1 105.622 83.619 105.802 83.659 ;
      RECT MASK 1 106.12 83.619 106.3 83.659 ;
      RECT MASK 1 106.784 83.619 106.964 83.659 ;
      RECT MASK 1 107.282 83.619 107.462 83.659 ;
      RECT MASK 1 107.946 83.619 108.126 83.659 ;
      RECT MASK 1 108.444 83.619 108.624 83.659 ;
      RECT MASK 1 109.108 83.619 109.288 83.659 ;
      RECT MASK 1 116.462 83.76 116.522 84.81 ;
      RECT MASK 1 116.736 83.76 116.796 84.81 ;
      RECT MASK 1 117.01 83.76 117.07 84.81 ;
      RECT MASK 1 117.284 83.76 117.344 84.81 ;
      RECT MASK 1 117.558 83.76 117.618 84.81 ;
      RECT MASK 1 117.832 83.76 117.892 84.81 ;
      RECT MASK 1 118.106 83.76 118.166 84.81 ;
      RECT MASK 1 118.38 83.76 118.44 84.81 ;
      RECT MASK 1 118.654 83.76 118.714 84.81 ;
      RECT MASK 1 118.928 83.76 118.988 84.81 ;
      RECT MASK 1 119.202 83.76 119.262 84.81 ;
      RECT MASK 1 119.476 83.76 119.536 84.81 ;
      RECT MASK 1 119.75 83.76 119.81 84.81 ;
      RECT MASK 1 120.024 83.76 120.084 84.81 ;
      RECT MASK 1 120.298 83.76 120.358 84.81 ;
      RECT MASK 1 120.572 83.76 120.632 84.81 ;
      RECT MASK 1 120.846 83.76 120.906 84.81 ;
      RECT MASK 1 121.12 83.76 121.18 84.81 ;
      RECT MASK 1 121.394 83.76 121.454 84.81 ;
      RECT MASK 1 121.668 83.76 121.728 84.81 ;
      RECT MASK 1 121.942 83.76 122.002 84.81 ;
      RECT MASK 1 122.216 83.76 122.276 84.81 ;
      RECT MASK 1 122.49 83.76 122.55 84.81 ;
      RECT MASK 1 122.764 83.76 122.824 84.81 ;
      RECT MASK 1 123.038 83.76 123.098 84.81 ;
      RECT MASK 1 123.312 83.76 123.372 84.81 ;
      RECT MASK 1 123.586 83.76 123.646 84.81 ;
      RECT MASK 1 123.86 83.76 123.92 84.81 ;
      RECT MASK 1 124.134 83.76 124.194 84.81 ;
      RECT MASK 1 124.408 83.76 124.468 84.81 ;
      RECT MASK 1 124.682 83.76 124.742 84.81 ;
      RECT MASK 1 124.956 83.76 125.016 84.81 ;
      RECT MASK 1 125.23 83.76 125.29 84.81 ;
      RECT MASK 1 125.504 83.76 125.564 84.81 ;
      RECT MASK 1 125.778 83.76 125.838 84.81 ;
      RECT MASK 1 126.052 83.76 126.112 84.81 ;
      RECT MASK 1 126.326 83.76 126.386 84.81 ;
      RECT MASK 1 126.6 83.76 126.66 84.81 ;
      RECT MASK 1 126.874 83.76 126.934 84.81 ;
      RECT MASK 1 127.148 83.76 127.208 84.81 ;
      RECT MASK 1 127.422 83.76 127.482 84.81 ;
      RECT MASK 1 127.696 83.76 127.756 84.81 ;
      RECT MASK 1 6.193 83.841 109.945 83.881 ;
      RECT MASK 1 6.193 84.109 6.857 84.149 ;
      RECT MASK 1 10.177 84.109 10.675 84.149 ;
      RECT MASK 1 11.649 84.109 12.313 84.149 ;
      RECT MASK 1 16.795 84.109 17.293 84.149 ;
      RECT MASK 1 18.267 84.109 18.931 84.149 ;
      RECT MASK 1 23.413 84.109 23.911 84.149 ;
      RECT MASK 1 24.885 84.109 25.549 84.149 ;
      RECT MASK 1 30.031 84.109 30.529 84.149 ;
      RECT MASK 1 31.503 84.109 32.167 84.149 ;
      RECT MASK 1 36.649 84.109 37.147 84.149 ;
      RECT MASK 1 38.121 84.109 38.785 84.149 ;
      RECT MASK 1 43.267 84.109 43.765 84.149 ;
      RECT MASK 1 44.739 84.109 45.403 84.149 ;
      RECT MASK 1 49.885 84.109 50.383 84.149 ;
      RECT MASK 1 51.357 84.109 52.021 84.149 ;
      RECT MASK 1 56.503 84.109 57.001 84.149 ;
      RECT MASK 1 57.975 84.109 58.6695 84.149 ;
      RECT MASK 1 63.121 84.109 63.619 84.149 ;
      RECT MASK 1 64.593 84.109 65.257 84.149 ;
      RECT MASK 1 69.739 84.109 70.237 84.149 ;
      RECT MASK 1 71.211 84.109 71.875 84.149 ;
      RECT MASK 1 76.357 84.109 76.855 84.149 ;
      RECT MASK 1 77.829 84.109 78.493 84.149 ;
      RECT MASK 1 82.975 84.109 83.473 84.149 ;
      RECT MASK 1 84.447 84.109 85.111 84.149 ;
      RECT MASK 1 89.593 84.109 90.091 84.149 ;
      RECT MASK 1 91.065 84.109 91.729 84.149 ;
      RECT MASK 1 96.211 84.109 96.709 84.149 ;
      RECT MASK 1 97.683 84.109 98.347 84.149 ;
      RECT MASK 1 102.829 84.109 103.327 84.149 ;
      RECT MASK 1 104.301 84.109 104.965 84.149 ;
      RECT MASK 1 109.447 84.109 109.945 84.149 ;
      RECT MASK 1 7.051 84.19 7.66 84.23 ;
      RECT MASK 1 8.213 84.19 8.822 84.23 ;
      RECT MASK 1 9.375 84.19 9.984 84.23 ;
      RECT MASK 1 12.507 84.19 13.116 84.23 ;
      RECT MASK 1 13.669 84.19 14.278 84.23 ;
      RECT MASK 1 14.831 84.19 15.44 84.23 ;
      RECT MASK 1 15.993 84.19 16.602 84.23 ;
      RECT MASK 1 19.125 84.19 19.734 84.23 ;
      RECT MASK 1 20.287 84.19 20.896 84.23 ;
      RECT MASK 1 21.449 84.19 22.058 84.23 ;
      RECT MASK 1 22.611 84.19 23.22 84.23 ;
      RECT MASK 1 25.743 84.19 26.352 84.23 ;
      RECT MASK 1 26.905 84.19 27.514 84.23 ;
      RECT MASK 1 28.067 84.19 28.676 84.23 ;
      RECT MASK 1 29.229 84.19 29.838 84.23 ;
      RECT MASK 1 32.361 84.19 32.97 84.23 ;
      RECT MASK 1 33.523 84.19 34.132 84.23 ;
      RECT MASK 1 34.685 84.19 35.294 84.23 ;
      RECT MASK 1 35.847 84.19 36.456 84.23 ;
      RECT MASK 1 38.979 84.19 39.588 84.23 ;
      RECT MASK 1 40.141 84.19 40.75 84.23 ;
      RECT MASK 1 41.303 84.19 41.912 84.23 ;
      RECT MASK 1 42.465 84.19 43.074 84.23 ;
      RECT MASK 1 45.597 84.19 46.206 84.23 ;
      RECT MASK 1 46.759 84.19 47.368 84.23 ;
      RECT MASK 1 47.921 84.19 48.53 84.23 ;
      RECT MASK 1 49.083 84.19 49.692 84.23 ;
      RECT MASK 1 52.215 84.19 52.824 84.23 ;
      RECT MASK 1 53.377 84.19 53.986 84.23 ;
      RECT MASK 1 54.539 84.19 55.148 84.23 ;
      RECT MASK 1 55.701 84.19 56.31 84.23 ;
      RECT MASK 1 58.833 84.19 59.442 84.23 ;
      RECT MASK 1 59.995 84.19 60.604 84.23 ;
      RECT MASK 1 61.157 84.19 61.766 84.23 ;
      RECT MASK 1 62.319 84.19 62.928 84.23 ;
      RECT MASK 1 65.451 84.19 66.06 84.23 ;
      RECT MASK 1 66.613 84.19 67.222 84.23 ;
      RECT MASK 1 67.775 84.19 68.384 84.23 ;
      RECT MASK 1 68.937 84.19 69.546 84.23 ;
      RECT MASK 1 72.069 84.19 72.678 84.23 ;
      RECT MASK 1 73.231 84.19 73.84 84.23 ;
      RECT MASK 1 74.393 84.19 75.002 84.23 ;
      RECT MASK 1 75.555 84.19 76.164 84.23 ;
      RECT MASK 1 78.687 84.19 79.296 84.23 ;
      RECT MASK 1 79.849 84.19 80.458 84.23 ;
      RECT MASK 1 81.011 84.19 81.62 84.23 ;
      RECT MASK 1 82.173 84.19 82.782 84.23 ;
      RECT MASK 1 85.305 84.19 85.914 84.23 ;
      RECT MASK 1 86.467 84.19 87.076 84.23 ;
      RECT MASK 1 87.629 84.19 88.238 84.23 ;
      RECT MASK 1 88.791 84.19 89.4 84.23 ;
      RECT MASK 1 91.923 84.19 92.532 84.23 ;
      RECT MASK 1 93.085 84.19 93.694 84.23 ;
      RECT MASK 1 94.247 84.19 94.856 84.23 ;
      RECT MASK 1 95.409 84.19 96.018 84.23 ;
      RECT MASK 1 98.541 84.19 99.15 84.23 ;
      RECT MASK 1 99.703 84.19 100.312 84.23 ;
      RECT MASK 1 100.865 84.19 101.474 84.23 ;
      RECT MASK 1 102.027 84.19 102.636 84.23 ;
      RECT MASK 1 105.159 84.19 105.768 84.23 ;
      RECT MASK 1 106.321 84.19 106.93 84.23 ;
      RECT MASK 1 107.483 84.19 108.092 84.23 ;
      RECT MASK 1 108.645 84.19 109.254 84.23 ;
      RECT MASK 1 2.067 84.39 2.127 85.44 ;
      RECT MASK 1 2.341 84.39 2.401 85.44 ;
      RECT MASK 1 2.615 84.39 2.675 85.44 ;
      RECT MASK 1 2.889 84.39 2.949 85.44 ;
      RECT MASK 1 3.163 84.39 3.223 85.44 ;
      RECT MASK 1 3.437 84.39 3.497 85.44 ;
      RECT MASK 1 3.711 84.39 3.771 85.44 ;
      RECT MASK 1 3.985 84.39 4.045 85.44 ;
      RECT MASK 1 4.259 84.39 4.319 85.44 ;
      RECT MASK 1 4.533 84.39 4.593 85.44 ;
      RECT MASK 1 6.224 84.569 109.907 84.609 ;
      RECT MASK 1 6.269 84.791 6.449 84.831 ;
      RECT MASK 1 6.85 84.791 7.03 84.831 ;
      RECT MASK 1 7.514 84.791 7.694 84.831 ;
      RECT MASK 1 8.012 84.791 8.192 84.831 ;
      RECT MASK 1 8.676 84.791 8.856 84.831 ;
      RECT MASK 1 9.174 84.791 9.354 84.831 ;
      RECT MASK 1 9.838 84.791 10.018 84.831 ;
      RECT MASK 1 10.419 84.791 10.599 84.831 ;
      RECT MASK 1 11.725 84.791 11.905 84.831 ;
      RECT MASK 1 12.306 84.791 12.486 84.831 ;
      RECT MASK 1 12.97 84.791 13.15 84.831 ;
      RECT MASK 1 13.468 84.791 13.648 84.831 ;
      RECT MASK 1 14.132 84.791 14.312 84.831 ;
      RECT MASK 1 14.63 84.791 14.81 84.831 ;
      RECT MASK 1 15.294 84.791 15.474 84.831 ;
      RECT MASK 1 15.792 84.791 15.972 84.831 ;
      RECT MASK 1 16.456 84.791 16.636 84.831 ;
      RECT MASK 1 17.037 84.791 17.217 84.831 ;
      RECT MASK 1 18.343 84.791 18.523 84.831 ;
      RECT MASK 1 18.924 84.791 19.104 84.831 ;
      RECT MASK 1 19.588 84.791 19.768 84.831 ;
      RECT MASK 1 20.086 84.791 20.266 84.831 ;
      RECT MASK 1 20.75 84.791 20.93 84.831 ;
      RECT MASK 1 21.248 84.791 21.428 84.831 ;
      RECT MASK 1 21.912 84.791 22.092 84.831 ;
      RECT MASK 1 22.41 84.791 22.59 84.831 ;
      RECT MASK 1 23.074 84.791 23.254 84.831 ;
      RECT MASK 1 23.655 84.791 23.835 84.831 ;
      RECT MASK 1 24.961 84.791 25.141 84.831 ;
      RECT MASK 1 25.542 84.791 25.722 84.831 ;
      RECT MASK 1 26.206 84.791 26.386 84.831 ;
      RECT MASK 1 26.704 84.791 26.884 84.831 ;
      RECT MASK 1 27.368 84.791 27.548 84.831 ;
      RECT MASK 1 27.866 84.791 28.046 84.831 ;
      RECT MASK 1 28.53 84.791 28.71 84.831 ;
      RECT MASK 1 29.028 84.791 29.208 84.831 ;
      RECT MASK 1 29.692 84.791 29.872 84.831 ;
      RECT MASK 1 30.273 84.791 30.453 84.831 ;
      RECT MASK 1 31.579 84.791 31.759 84.831 ;
      RECT MASK 1 32.16 84.791 32.34 84.831 ;
      RECT MASK 1 32.824 84.791 33.004 84.831 ;
      RECT MASK 1 33.322 84.791 33.502 84.831 ;
      RECT MASK 1 33.986 84.791 34.166 84.831 ;
      RECT MASK 1 34.484 84.791 34.664 84.831 ;
      RECT MASK 1 35.148 84.791 35.328 84.831 ;
      RECT MASK 1 35.646 84.791 35.826 84.831 ;
      RECT MASK 1 36.31 84.791 36.49 84.831 ;
      RECT MASK 1 36.891 84.791 37.071 84.831 ;
      RECT MASK 1 38.197 84.791 38.377 84.831 ;
      RECT MASK 1 38.778 84.791 38.958 84.831 ;
      RECT MASK 1 39.442 84.791 39.622 84.831 ;
      RECT MASK 1 39.94 84.791 40.12 84.831 ;
      RECT MASK 1 40.604 84.791 40.784 84.831 ;
      RECT MASK 1 41.102 84.791 41.282 84.831 ;
      RECT MASK 1 41.766 84.791 41.946 84.831 ;
      RECT MASK 1 42.264 84.791 42.444 84.831 ;
      RECT MASK 1 42.928 84.791 43.108 84.831 ;
      RECT MASK 1 43.509 84.791 43.689 84.831 ;
      RECT MASK 1 44.815 84.791 44.995 84.831 ;
      RECT MASK 1 45.396 84.791 45.576 84.831 ;
      RECT MASK 1 46.06 84.791 46.24 84.831 ;
      RECT MASK 1 46.558 84.791 46.738 84.831 ;
      RECT MASK 1 47.222 84.791 47.402 84.831 ;
      RECT MASK 1 47.72 84.791 47.9 84.831 ;
      RECT MASK 1 48.384 84.791 48.564 84.831 ;
      RECT MASK 1 48.882 84.791 49.062 84.831 ;
      RECT MASK 1 49.546 84.791 49.726 84.831 ;
      RECT MASK 1 50.127 84.791 50.307 84.831 ;
      RECT MASK 1 51.433 84.791 51.613 84.831 ;
      RECT MASK 1 52.014 84.791 52.194 84.831 ;
      RECT MASK 1 52.678 84.791 52.858 84.831 ;
      RECT MASK 1 53.176 84.791 53.356 84.831 ;
      RECT MASK 1 53.84 84.791 54.02 84.831 ;
      RECT MASK 1 54.338 84.791 54.518 84.831 ;
      RECT MASK 1 55.002 84.791 55.182 84.831 ;
      RECT MASK 1 55.5 84.791 55.68 84.831 ;
      RECT MASK 1 56.164 84.791 56.344 84.831 ;
      RECT MASK 1 56.745 84.791 56.925 84.831 ;
      RECT MASK 1 58.051 84.791 58.231 84.831 ;
      RECT MASK 1 58.632 84.791 58.812 84.831 ;
      RECT MASK 1 59.296 84.791 59.476 84.831 ;
      RECT MASK 1 59.794 84.791 59.974 84.831 ;
      RECT MASK 1 60.458 84.791 60.638 84.831 ;
      RECT MASK 1 60.956 84.791 61.136 84.831 ;
      RECT MASK 1 61.62 84.791 61.8 84.831 ;
      RECT MASK 1 62.118 84.791 62.298 84.831 ;
      RECT MASK 1 62.782 84.791 62.962 84.831 ;
      RECT MASK 1 63.363 84.791 63.543 84.831 ;
      RECT MASK 1 64.669 84.791 64.849 84.831 ;
      RECT MASK 1 65.25 84.791 65.43 84.831 ;
      RECT MASK 1 65.914 84.791 66.094 84.831 ;
      RECT MASK 1 66.412 84.791 66.592 84.831 ;
      RECT MASK 1 67.076 84.791 67.256 84.831 ;
      RECT MASK 1 67.574 84.791 67.754 84.831 ;
      RECT MASK 1 68.238 84.791 68.418 84.831 ;
      RECT MASK 1 68.736 84.791 68.916 84.831 ;
      RECT MASK 1 69.4 84.791 69.58 84.831 ;
      RECT MASK 1 69.981 84.791 70.161 84.831 ;
      RECT MASK 1 71.287 84.791 71.467 84.831 ;
      RECT MASK 1 71.868 84.791 72.048 84.831 ;
      RECT MASK 1 72.532 84.791 72.712 84.831 ;
      RECT MASK 1 73.03 84.791 73.21 84.831 ;
      RECT MASK 1 73.694 84.791 73.874 84.831 ;
      RECT MASK 1 74.192 84.791 74.372 84.831 ;
      RECT MASK 1 74.856 84.791 75.036 84.831 ;
      RECT MASK 1 75.354 84.791 75.534 84.831 ;
      RECT MASK 1 76.018 84.791 76.198 84.831 ;
      RECT MASK 1 76.599 84.791 76.779 84.831 ;
      RECT MASK 1 77.905 84.791 78.085 84.831 ;
      RECT MASK 1 78.486 84.791 78.666 84.831 ;
      RECT MASK 1 79.15 84.791 79.33 84.831 ;
      RECT MASK 1 79.648 84.791 79.828 84.831 ;
      RECT MASK 1 80.312 84.791 80.492 84.831 ;
      RECT MASK 1 80.81 84.791 80.99 84.831 ;
      RECT MASK 1 81.474 84.791 81.654 84.831 ;
      RECT MASK 1 81.972 84.791 82.152 84.831 ;
      RECT MASK 1 82.636 84.791 82.816 84.831 ;
      RECT MASK 1 83.217 84.791 83.397 84.831 ;
      RECT MASK 1 84.523 84.791 84.703 84.831 ;
      RECT MASK 1 85.104 84.791 85.284 84.831 ;
      RECT MASK 1 85.768 84.791 85.948 84.831 ;
      RECT MASK 1 86.266 84.791 86.446 84.831 ;
      RECT MASK 1 86.93 84.791 87.11 84.831 ;
      RECT MASK 1 87.428 84.791 87.608 84.831 ;
      RECT MASK 1 88.092 84.791 88.272 84.831 ;
      RECT MASK 1 88.59 84.791 88.77 84.831 ;
      RECT MASK 1 89.254 84.791 89.434 84.831 ;
      RECT MASK 1 89.835 84.791 90.015 84.831 ;
      RECT MASK 1 91.141 84.791 91.321 84.831 ;
      RECT MASK 1 91.722 84.791 91.902 84.831 ;
      RECT MASK 1 92.386 84.791 92.566 84.831 ;
      RECT MASK 1 92.884 84.791 93.064 84.831 ;
      RECT MASK 1 93.548 84.791 93.728 84.831 ;
      RECT MASK 1 94.046 84.791 94.226 84.831 ;
      RECT MASK 1 94.71 84.791 94.89 84.831 ;
      RECT MASK 1 95.208 84.791 95.388 84.831 ;
      RECT MASK 1 95.872 84.791 96.052 84.831 ;
      RECT MASK 1 96.453 84.791 96.633 84.831 ;
      RECT MASK 1 97.759 84.791 97.939 84.831 ;
      RECT MASK 1 98.34 84.791 98.52 84.831 ;
      RECT MASK 1 99.004 84.791 99.184 84.831 ;
      RECT MASK 1 99.502 84.791 99.682 84.831 ;
      RECT MASK 1 100.166 84.791 100.346 84.831 ;
      RECT MASK 1 100.664 84.791 100.844 84.831 ;
      RECT MASK 1 101.328 84.791 101.508 84.831 ;
      RECT MASK 1 101.826 84.791 102.006 84.831 ;
      RECT MASK 1 102.49 84.791 102.67 84.831 ;
      RECT MASK 1 103.071 84.791 103.251 84.831 ;
      RECT MASK 1 104.377 84.791 104.557 84.831 ;
      RECT MASK 1 104.958 84.791 105.138 84.831 ;
      RECT MASK 1 105.622 84.791 105.802 84.831 ;
      RECT MASK 1 106.12 84.791 106.3 84.831 ;
      RECT MASK 1 106.784 84.791 106.964 84.831 ;
      RECT MASK 1 107.282 84.791 107.462 84.831 ;
      RECT MASK 1 107.946 84.791 108.126 84.831 ;
      RECT MASK 1 108.444 84.791 108.624 84.831 ;
      RECT MASK 1 109.108 84.791 109.288 84.831 ;
      RECT MASK 1 109.689 84.791 109.869 84.831 ;
      RECT MASK 1 11.039 84.9185 11.119 85.141 ;
      RECT MASK 1 11.371 84.9185 11.451 85.141 ;
      RECT MASK 1 17.657 84.9185 17.737 85.141 ;
      RECT MASK 1 17.989 84.9185 18.069 85.141 ;
      RECT MASK 1 24.275 84.9185 24.355 85.141 ;
      RECT MASK 1 24.607 84.9185 24.687 85.141 ;
      RECT MASK 1 30.893 84.9185 30.973 85.141 ;
      RECT MASK 1 31.225 84.9185 31.305 85.141 ;
      RECT MASK 1 37.511 84.9185 37.591 85.141 ;
      RECT MASK 1 37.843 84.9185 37.923 85.141 ;
      RECT MASK 1 44.129 84.9185 44.209 85.141 ;
      RECT MASK 1 44.461 84.9185 44.541 85.141 ;
      RECT MASK 1 50.747 84.9185 50.827 85.141 ;
      RECT MASK 1 51.079 84.9185 51.159 85.141 ;
      RECT MASK 1 57.365 84.9185 57.445 85.141 ;
      RECT MASK 1 57.697 84.9185 57.777 85.141 ;
      RECT MASK 1 63.983 84.9185 64.063 85.141 ;
      RECT MASK 1 64.315 84.9185 64.395 85.141 ;
      RECT MASK 1 70.601 84.9185 70.681 85.141 ;
      RECT MASK 1 70.933 84.9185 71.013 85.141 ;
      RECT MASK 1 77.219 84.9185 77.299 85.141 ;
      RECT MASK 1 77.551 84.9185 77.631 85.141 ;
      RECT MASK 1 83.837 84.9185 83.917 85.141 ;
      RECT MASK 1 84.169 84.9185 84.249 85.141 ;
      RECT MASK 1 90.455 84.9185 90.535 85.141 ;
      RECT MASK 1 90.787 84.9185 90.867 85.141 ;
      RECT MASK 1 97.073 84.9185 97.153 85.141 ;
      RECT MASK 1 97.405 84.9185 97.485 85.141 ;
      RECT MASK 1 103.691 84.9185 103.771 85.141 ;
      RECT MASK 1 104.023 84.9185 104.103 85.141 ;
      RECT MASK 1 6.269 84.959 6.449 84.999 ;
      RECT MASK 1 10.419 84.959 10.599 84.999 ;
      RECT MASK 1 11.725 84.959 11.905 84.999 ;
      RECT MASK 1 17.037 84.959 17.217 84.999 ;
      RECT MASK 1 18.343 84.959 18.523 84.999 ;
      RECT MASK 1 23.655 84.959 23.835 84.999 ;
      RECT MASK 1 24.961 84.959 25.141 84.999 ;
      RECT MASK 1 30.273 84.959 30.453 84.999 ;
      RECT MASK 1 31.579 84.959 31.759 84.999 ;
      RECT MASK 1 36.891 84.959 37.071 84.999 ;
      RECT MASK 1 38.197 84.959 38.377 84.999 ;
      RECT MASK 1 43.509 84.959 43.689 84.999 ;
      RECT MASK 1 44.815 84.959 44.995 84.999 ;
      RECT MASK 1 50.127 84.959 50.307 84.999 ;
      RECT MASK 1 51.433 84.959 51.613 84.999 ;
      RECT MASK 1 56.745 84.959 56.925 84.999 ;
      RECT MASK 1 58.051 84.959 58.231 84.999 ;
      RECT MASK 1 63.363 84.959 63.543 84.999 ;
      RECT MASK 1 64.669 84.959 64.849 84.999 ;
      RECT MASK 1 69.981 84.959 70.161 84.999 ;
      RECT MASK 1 71.287 84.959 71.467 84.999 ;
      RECT MASK 1 76.599 84.959 76.779 84.999 ;
      RECT MASK 1 77.905 84.959 78.085 84.999 ;
      RECT MASK 1 83.217 84.959 83.397 84.999 ;
      RECT MASK 1 84.523 84.959 84.703 84.999 ;
      RECT MASK 1 89.835 84.959 90.015 84.999 ;
      RECT MASK 1 91.141 84.959 91.321 84.999 ;
      RECT MASK 1 96.453 84.959 96.633 84.999 ;
      RECT MASK 1 97.759 84.959 97.939 84.999 ;
      RECT MASK 1 103.071 84.959 103.251 84.999 ;
      RECT MASK 1 104.377 84.959 104.557 84.999 ;
      RECT MASK 1 109.689 84.959 109.869 84.999 ;
      RECT MASK 1 6.978 85.013 7.161 85.053 ;
      RECT MASK 1 7.383 85.013 7.566 85.053 ;
      RECT MASK 1 8.14 85.013 8.323 85.053 ;
      RECT MASK 1 8.545 85.013 8.728 85.053 ;
      RECT MASK 1 9.302 85.013 9.485 85.053 ;
      RECT MASK 1 9.707 85.013 9.89 85.053 ;
      RECT MASK 1 12.434 85.013 12.617 85.053 ;
      RECT MASK 1 12.839 85.013 13.022 85.053 ;
      RECT MASK 1 13.596 85.013 13.779 85.053 ;
      RECT MASK 1 14.001 85.013 14.184 85.053 ;
      RECT MASK 1 14.758 85.013 14.941 85.053 ;
      RECT MASK 1 15.163 85.013 15.346 85.053 ;
      RECT MASK 1 15.92 85.013 16.103 85.053 ;
      RECT MASK 1 16.325 85.013 16.508 85.053 ;
      RECT MASK 1 19.052 85.013 19.235 85.053 ;
      RECT MASK 1 19.457 85.013 19.64 85.053 ;
      RECT MASK 1 20.214 85.013 20.397 85.053 ;
      RECT MASK 1 20.619 85.013 20.802 85.053 ;
      RECT MASK 1 21.376 85.013 21.559 85.053 ;
      RECT MASK 1 21.781 85.013 21.964 85.053 ;
      RECT MASK 1 22.538 85.013 22.721 85.053 ;
      RECT MASK 1 22.943 85.013 23.126 85.053 ;
      RECT MASK 1 25.67 85.013 25.853 85.053 ;
      RECT MASK 1 26.075 85.013 26.258 85.053 ;
      RECT MASK 1 26.832 85.013 27.015 85.053 ;
      RECT MASK 1 27.237 85.013 27.42 85.053 ;
      RECT MASK 1 27.994 85.013 28.177 85.053 ;
      RECT MASK 1 28.399 85.013 28.582 85.053 ;
      RECT MASK 1 29.156 85.013 29.339 85.053 ;
      RECT MASK 1 29.561 85.013 29.744 85.053 ;
      RECT MASK 1 32.288 85.013 32.471 85.053 ;
      RECT MASK 1 32.693 85.013 32.876 85.053 ;
      RECT MASK 1 33.45 85.013 33.633 85.053 ;
      RECT MASK 1 33.855 85.013 34.038 85.053 ;
      RECT MASK 1 34.612 85.013 34.795 85.053 ;
      RECT MASK 1 35.017 85.013 35.2 85.053 ;
      RECT MASK 1 35.774 85.013 35.957 85.053 ;
      RECT MASK 1 36.179 85.013 36.362 85.053 ;
      RECT MASK 1 38.906 85.013 39.089 85.053 ;
      RECT MASK 1 39.311 85.013 39.494 85.053 ;
      RECT MASK 1 40.068 85.013 40.251 85.053 ;
      RECT MASK 1 40.473 85.013 40.656 85.053 ;
      RECT MASK 1 41.23 85.013 41.413 85.053 ;
      RECT MASK 1 41.635 85.013 41.818 85.053 ;
      RECT MASK 1 42.392 85.013 42.575 85.053 ;
      RECT MASK 1 42.797 85.013 42.98 85.053 ;
      RECT MASK 1 45.524 85.013 45.707 85.053 ;
      RECT MASK 1 45.929 85.013 46.112 85.053 ;
      RECT MASK 1 46.686 85.013 46.869 85.053 ;
      RECT MASK 1 47.091 85.013 47.274 85.053 ;
      RECT MASK 1 47.848 85.013 48.031 85.053 ;
      RECT MASK 1 48.253 85.013 48.436 85.053 ;
      RECT MASK 1 49.01 85.013 49.193 85.053 ;
      RECT MASK 1 49.415 85.013 49.598 85.053 ;
      RECT MASK 1 52.142 85.013 52.325 85.053 ;
      RECT MASK 1 52.547 85.013 52.73 85.053 ;
      RECT MASK 1 53.304 85.013 53.487 85.053 ;
      RECT MASK 1 53.709 85.013 53.892 85.053 ;
      RECT MASK 1 54.466 85.013 54.649 85.053 ;
      RECT MASK 1 54.871 85.013 55.054 85.053 ;
      RECT MASK 1 55.628 85.013 55.811 85.053 ;
      RECT MASK 1 56.033 85.013 56.216 85.053 ;
      RECT MASK 1 58.76 85.013 58.943 85.053 ;
      RECT MASK 1 59.165 85.013 59.348 85.053 ;
      RECT MASK 1 59.922 85.013 60.105 85.053 ;
      RECT MASK 1 60.327 85.013 60.51 85.053 ;
      RECT MASK 1 61.084 85.013 61.267 85.053 ;
      RECT MASK 1 61.489 85.013 61.672 85.053 ;
      RECT MASK 1 62.246 85.013 62.429 85.053 ;
      RECT MASK 1 62.651 85.013 62.834 85.053 ;
      RECT MASK 1 65.378 85.013 65.561 85.053 ;
      RECT MASK 1 65.783 85.013 65.966 85.053 ;
      RECT MASK 1 66.54 85.013 66.723 85.053 ;
      RECT MASK 1 66.945 85.013 67.128 85.053 ;
      RECT MASK 1 67.702 85.013 67.885 85.053 ;
      RECT MASK 1 68.107 85.013 68.29 85.053 ;
      RECT MASK 1 68.864 85.013 69.047 85.053 ;
      RECT MASK 1 69.269 85.013 69.452 85.053 ;
      RECT MASK 1 71.996 85.013 72.179 85.053 ;
      RECT MASK 1 72.401 85.013 72.584 85.053 ;
      RECT MASK 1 73.158 85.013 73.341 85.053 ;
      RECT MASK 1 73.563 85.013 73.746 85.053 ;
      RECT MASK 1 74.32 85.013 74.503 85.053 ;
      RECT MASK 1 74.725 85.013 74.908 85.053 ;
      RECT MASK 1 75.482 85.013 75.665 85.053 ;
      RECT MASK 1 75.887 85.013 76.07 85.053 ;
      RECT MASK 1 78.614 85.013 78.797 85.053 ;
      RECT MASK 1 79.019 85.013 79.202 85.053 ;
      RECT MASK 1 79.776 85.013 79.959 85.053 ;
      RECT MASK 1 80.181 85.013 80.364 85.053 ;
      RECT MASK 1 80.938 85.013 81.121 85.053 ;
      RECT MASK 1 81.343 85.013 81.526 85.053 ;
      RECT MASK 1 82.1 85.013 82.283 85.053 ;
      RECT MASK 1 82.505 85.013 82.688 85.053 ;
      RECT MASK 1 85.232 85.013 85.415 85.053 ;
      RECT MASK 1 85.637 85.013 85.82 85.053 ;
      RECT MASK 1 86.394 85.013 86.577 85.053 ;
      RECT MASK 1 86.799 85.013 86.982 85.053 ;
      RECT MASK 1 87.556 85.013 87.739 85.053 ;
      RECT MASK 1 87.961 85.013 88.144 85.053 ;
      RECT MASK 1 88.718 85.013 88.901 85.053 ;
      RECT MASK 1 89.123 85.013 89.306 85.053 ;
      RECT MASK 1 91.85 85.013 92.033 85.053 ;
      RECT MASK 1 92.255 85.013 92.438 85.053 ;
      RECT MASK 1 93.012 85.013 93.195 85.053 ;
      RECT MASK 1 93.417 85.013 93.6 85.053 ;
      RECT MASK 1 94.174 85.013 94.357 85.053 ;
      RECT MASK 1 94.579 85.013 94.762 85.053 ;
      RECT MASK 1 95.336 85.013 95.519 85.053 ;
      RECT MASK 1 95.741 85.013 95.924 85.053 ;
      RECT MASK 1 98.468 85.013 98.651 85.053 ;
      RECT MASK 1 98.873 85.013 99.056 85.053 ;
      RECT MASK 1 99.63 85.013 99.813 85.053 ;
      RECT MASK 1 100.035 85.013 100.218 85.053 ;
      RECT MASK 1 100.792 85.013 100.975 85.053 ;
      RECT MASK 1 101.197 85.013 101.38 85.053 ;
      RECT MASK 1 101.954 85.013 102.137 85.053 ;
      RECT MASK 1 102.359 85.013 102.542 85.053 ;
      RECT MASK 1 105.086 85.013 105.269 85.053 ;
      RECT MASK 1 105.491 85.013 105.674 85.053 ;
      RECT MASK 1 106.248 85.013 106.431 85.053 ;
      RECT MASK 1 106.653 85.013 106.836 85.053 ;
      RECT MASK 1 107.41 85.013 107.593 85.053 ;
      RECT MASK 1 107.815 85.013 107.998 85.053 ;
      RECT MASK 1 108.572 85.013 108.755 85.053 ;
      RECT MASK 1 108.977 85.013 109.16 85.053 ;
      RECT MASK 1 6.978 85.181 7.161 85.221 ;
      RECT MASK 1 7.383 85.181 7.566 85.221 ;
      RECT MASK 1 8.14 85.181 8.323 85.221 ;
      RECT MASK 1 8.545 85.181 8.728 85.221 ;
      RECT MASK 1 9.302 85.181 9.485 85.221 ;
      RECT MASK 1 9.707 85.181 9.89 85.221 ;
      RECT MASK 1 12.434 85.181 12.617 85.221 ;
      RECT MASK 1 12.839 85.181 13.022 85.221 ;
      RECT MASK 1 13.596 85.181 13.779 85.221 ;
      RECT MASK 1 14.001 85.181 14.184 85.221 ;
      RECT MASK 1 14.758 85.181 14.941 85.221 ;
      RECT MASK 1 15.163 85.181 15.346 85.221 ;
      RECT MASK 1 15.92 85.181 16.103 85.221 ;
      RECT MASK 1 16.325 85.181 16.508 85.221 ;
      RECT MASK 1 19.052 85.181 19.235 85.221 ;
      RECT MASK 1 19.457 85.181 19.64 85.221 ;
      RECT MASK 1 20.214 85.181 20.397 85.221 ;
      RECT MASK 1 20.619 85.181 20.802 85.221 ;
      RECT MASK 1 21.376 85.181 21.559 85.221 ;
      RECT MASK 1 21.781 85.181 21.964 85.221 ;
      RECT MASK 1 22.538 85.181 22.721 85.221 ;
      RECT MASK 1 22.943 85.181 23.126 85.221 ;
      RECT MASK 1 25.67 85.181 25.853 85.221 ;
      RECT MASK 1 26.075 85.181 26.258 85.221 ;
      RECT MASK 1 26.832 85.181 27.015 85.221 ;
      RECT MASK 1 27.237 85.181 27.42 85.221 ;
      RECT MASK 1 27.994 85.181 28.177 85.221 ;
      RECT MASK 1 28.399 85.181 28.582 85.221 ;
      RECT MASK 1 29.156 85.181 29.339 85.221 ;
      RECT MASK 1 29.561 85.181 29.744 85.221 ;
      RECT MASK 1 32.288 85.181 32.471 85.221 ;
      RECT MASK 1 32.693 85.181 32.876 85.221 ;
      RECT MASK 1 33.45 85.181 33.633 85.221 ;
      RECT MASK 1 33.855 85.181 34.038 85.221 ;
      RECT MASK 1 34.612 85.181 34.795 85.221 ;
      RECT MASK 1 35.017 85.181 35.2 85.221 ;
      RECT MASK 1 35.774 85.181 35.957 85.221 ;
      RECT MASK 1 36.179 85.181 36.362 85.221 ;
      RECT MASK 1 38.906 85.181 39.089 85.221 ;
      RECT MASK 1 39.311 85.181 39.494 85.221 ;
      RECT MASK 1 40.068 85.181 40.251 85.221 ;
      RECT MASK 1 40.473 85.181 40.656 85.221 ;
      RECT MASK 1 41.23 85.181 41.413 85.221 ;
      RECT MASK 1 41.635 85.181 41.818 85.221 ;
      RECT MASK 1 42.392 85.181 42.575 85.221 ;
      RECT MASK 1 42.797 85.181 42.98 85.221 ;
      RECT MASK 1 45.524 85.181 45.707 85.221 ;
      RECT MASK 1 45.929 85.181 46.112 85.221 ;
      RECT MASK 1 46.686 85.181 46.869 85.221 ;
      RECT MASK 1 47.091 85.181 47.274 85.221 ;
      RECT MASK 1 47.848 85.181 48.031 85.221 ;
      RECT MASK 1 48.253 85.181 48.436 85.221 ;
      RECT MASK 1 49.01 85.181 49.193 85.221 ;
      RECT MASK 1 49.415 85.181 49.598 85.221 ;
      RECT MASK 1 52.142 85.181 52.325 85.221 ;
      RECT MASK 1 52.547 85.181 52.73 85.221 ;
      RECT MASK 1 53.304 85.181 53.487 85.221 ;
      RECT MASK 1 53.709 85.181 53.892 85.221 ;
      RECT MASK 1 54.466 85.181 54.649 85.221 ;
      RECT MASK 1 54.871 85.181 55.054 85.221 ;
      RECT MASK 1 55.628 85.181 55.811 85.221 ;
      RECT MASK 1 56.033 85.181 56.216 85.221 ;
      RECT MASK 1 58.76 85.181 58.943 85.221 ;
      RECT MASK 1 59.165 85.181 59.348 85.221 ;
      RECT MASK 1 59.922 85.181 60.105 85.221 ;
      RECT MASK 1 60.327 85.181 60.51 85.221 ;
      RECT MASK 1 61.084 85.181 61.267 85.221 ;
      RECT MASK 1 61.489 85.181 61.672 85.221 ;
      RECT MASK 1 62.246 85.181 62.429 85.221 ;
      RECT MASK 1 62.651 85.181 62.834 85.221 ;
      RECT MASK 1 65.378 85.181 65.561 85.221 ;
      RECT MASK 1 65.783 85.181 65.966 85.221 ;
      RECT MASK 1 66.54 85.181 66.723 85.221 ;
      RECT MASK 1 66.945 85.181 67.128 85.221 ;
      RECT MASK 1 67.702 85.181 67.885 85.221 ;
      RECT MASK 1 68.107 85.181 68.29 85.221 ;
      RECT MASK 1 68.864 85.181 69.047 85.221 ;
      RECT MASK 1 69.269 85.181 69.452 85.221 ;
      RECT MASK 1 71.996 85.181 72.179 85.221 ;
      RECT MASK 1 72.401 85.181 72.584 85.221 ;
      RECT MASK 1 73.158 85.181 73.341 85.221 ;
      RECT MASK 1 73.563 85.181 73.746 85.221 ;
      RECT MASK 1 74.32 85.181 74.503 85.221 ;
      RECT MASK 1 74.725 85.181 74.908 85.221 ;
      RECT MASK 1 75.482 85.181 75.665 85.221 ;
      RECT MASK 1 75.887 85.181 76.07 85.221 ;
      RECT MASK 1 78.614 85.181 78.797 85.221 ;
      RECT MASK 1 79.019 85.181 79.202 85.221 ;
      RECT MASK 1 79.776 85.181 79.959 85.221 ;
      RECT MASK 1 80.181 85.181 80.364 85.221 ;
      RECT MASK 1 80.938 85.181 81.121 85.221 ;
      RECT MASK 1 81.343 85.181 81.526 85.221 ;
      RECT MASK 1 82.1 85.181 82.283 85.221 ;
      RECT MASK 1 82.505 85.181 82.688 85.221 ;
      RECT MASK 1 85.232 85.181 85.415 85.221 ;
      RECT MASK 1 85.637 85.181 85.82 85.221 ;
      RECT MASK 1 86.394 85.181 86.577 85.221 ;
      RECT MASK 1 86.799 85.181 86.982 85.221 ;
      RECT MASK 1 87.556 85.181 87.739 85.221 ;
      RECT MASK 1 87.961 85.181 88.144 85.221 ;
      RECT MASK 1 88.718 85.181 88.901 85.221 ;
      RECT MASK 1 89.123 85.181 89.306 85.221 ;
      RECT MASK 1 91.85 85.181 92.033 85.221 ;
      RECT MASK 1 92.255 85.181 92.438 85.221 ;
      RECT MASK 1 93.012 85.181 93.195 85.221 ;
      RECT MASK 1 93.417 85.181 93.6 85.221 ;
      RECT MASK 1 94.174 85.181 94.357 85.221 ;
      RECT MASK 1 94.579 85.181 94.762 85.221 ;
      RECT MASK 1 95.336 85.181 95.519 85.221 ;
      RECT MASK 1 95.741 85.181 95.924 85.221 ;
      RECT MASK 1 98.468 85.181 98.651 85.221 ;
      RECT MASK 1 98.873 85.181 99.056 85.221 ;
      RECT MASK 1 99.63 85.181 99.813 85.221 ;
      RECT MASK 1 100.035 85.181 100.218 85.221 ;
      RECT MASK 1 100.792 85.181 100.975 85.221 ;
      RECT MASK 1 101.197 85.181 101.38 85.221 ;
      RECT MASK 1 101.954 85.181 102.137 85.221 ;
      RECT MASK 1 102.359 85.181 102.542 85.221 ;
      RECT MASK 1 105.086 85.181 105.269 85.221 ;
      RECT MASK 1 105.491 85.181 105.674 85.221 ;
      RECT MASK 1 106.248 85.181 106.431 85.221 ;
      RECT MASK 1 106.653 85.181 106.836 85.221 ;
      RECT MASK 1 107.41 85.181 107.593 85.221 ;
      RECT MASK 1 107.815 85.181 107.998 85.221 ;
      RECT MASK 1 108.572 85.181 108.755 85.221 ;
      RECT MASK 1 108.977 85.181 109.16 85.221 ;
      RECT MASK 1 6.224 85.365 109.898 85.405 ;
      RECT MASK 1 116.462 85.47 116.522 86.52 ;
      RECT MASK 1 116.736 85.47 116.796 86.52 ;
      RECT MASK 1 117.01 85.47 117.07 86.52 ;
      RECT MASK 1 117.284 85.47 117.344 86.52 ;
      RECT MASK 1 117.558 85.47 117.618 86.52 ;
      RECT MASK 1 117.832 85.47 117.892 86.52 ;
      RECT MASK 1 118.106 85.47 118.166 86.52 ;
      RECT MASK 1 118.38 85.47 118.44 86.52 ;
      RECT MASK 1 118.654 85.47 118.714 86.52 ;
      RECT MASK 1 118.928 85.47 118.988 86.52 ;
      RECT MASK 1 119.202 85.47 119.262 86.52 ;
      RECT MASK 1 119.476 85.47 119.536 86.52 ;
      RECT MASK 1 119.75 85.47 119.81 86.52 ;
      RECT MASK 1 120.024 85.47 120.084 86.52 ;
      RECT MASK 1 120.298 85.47 120.358 86.52 ;
      RECT MASK 1 120.572 85.47 120.632 86.52 ;
      RECT MASK 1 120.846 85.47 120.906 86.52 ;
      RECT MASK 1 121.12 85.47 121.18 86.52 ;
      RECT MASK 1 121.394 85.47 121.454 86.52 ;
      RECT MASK 1 121.668 85.47 121.728 86.52 ;
      RECT MASK 1 121.942 85.47 122.002 86.52 ;
      RECT MASK 1 122.216 85.47 122.276 86.52 ;
      RECT MASK 1 122.49 85.47 122.55 86.52 ;
      RECT MASK 1 122.764 85.47 122.824 86.52 ;
      RECT MASK 1 123.038 85.47 123.098 86.52 ;
      RECT MASK 1 123.312 85.47 123.372 86.52 ;
      RECT MASK 1 123.586 85.47 123.646 86.52 ;
      RECT MASK 1 123.86 85.47 123.92 86.52 ;
      RECT MASK 1 124.134 85.47 124.194 86.52 ;
      RECT MASK 1 124.408 85.47 124.468 86.52 ;
      RECT MASK 1 124.682 85.47 124.742 86.52 ;
      RECT MASK 1 124.956 85.47 125.016 86.52 ;
      RECT MASK 1 125.23 85.47 125.29 86.52 ;
      RECT MASK 1 125.504 85.47 125.564 86.52 ;
      RECT MASK 1 125.778 85.47 125.838 86.52 ;
      RECT MASK 1 126.052 85.47 126.112 86.52 ;
      RECT MASK 1 126.326 85.47 126.386 86.52 ;
      RECT MASK 1 126.6 85.47 126.66 86.52 ;
      RECT MASK 1 126.874 85.47 126.934 86.52 ;
      RECT MASK 1 127.148 85.47 127.208 86.52 ;
      RECT MASK 1 127.422 85.47 127.482 86.52 ;
      RECT MASK 1 127.696 85.47 127.756 86.52 ;
      RECT MASK 1 6.224 85.549 109.819 85.589 ;
      RECT MASK 1 6.224 85.885 109.826 85.925 ;
      RECT MASK 1 2.067 86.1 2.127 87.15 ;
      RECT MASK 1 2.341 86.1 2.401 87.15 ;
      RECT MASK 1 2.615 86.1 2.675 87.15 ;
      RECT MASK 1 2.889 86.1 2.949 87.15 ;
      RECT MASK 1 3.163 86.1 3.223 87.15 ;
      RECT MASK 1 3.437 86.1 3.497 87.15 ;
      RECT MASK 1 3.711 86.1 3.771 87.15 ;
      RECT MASK 1 3.985 86.1 4.045 87.15 ;
      RECT MASK 1 4.259 86.1 4.319 87.15 ;
      RECT MASK 1 4.533 86.1 4.593 87.15 ;
      RECT MASK 1 69.797 86.365 71.728 86.405 ;
      RECT MASK 1 103.854 86.365 105.785 86.405 ;
      RECT MASK 1 35.702 86.411 35.782 86.629 ;
      RECT MASK 1 67.02 86.411 67.1 86.629 ;
      RECT MASK 1 72.092 86.411 72.172 86.629 ;
      RECT MASK 1 103.41 86.411 103.49 86.629 ;
      RECT MASK 1 33.407 86.455 35.338 86.495 ;
      RECT MASK 1 67.472 86.455 69.229 86.495 ;
      RECT MASK 1 36.1535 86.469 66.6485 86.569 ;
      RECT MASK 1 72.5435 86.469 103.0385 86.569 ;
      RECT MASK 1 69.807 86.6735 69.887 95.0065 ;
      RECT MASK 1 105.695 86.6735 105.775 95.0065 ;
      RECT MASK 1 33.417 86.7635 33.497 94.9165 ;
      RECT MASK 1 69.139 86.7635 69.219 94.9165 ;
      RECT MASK 1 70.129 86.815 71.728 86.855 ;
      RECT MASK 1 103.854 86.815 105.453 86.855 ;
      RECT MASK 1 33.739 86.905 35.338 86.945 ;
      RECT MASK 1 67.472 86.905 68.897 86.945 ;
      RECT MASK 1 115.613 86.905 128.525 86.945 ;
      RECT MASK 1 35.702 87.011 35.782 94.668 ;
      RECT MASK 1 67.02 87.011 67.1 94.668 ;
      RECT MASK 1 72.102 87.011 72.162 87.452 ;
      RECT MASK 1 103.42 87.011 103.48 87.452 ;
      RECT MASK 1 70.139 87.1235 70.219 94.5565 ;
      RECT MASK 1 105.363 87.1235 105.443 94.5565 ;
      RECT MASK 1 36.326 87.147 66.476 87.207 ;
      RECT MASK 1 72.716 87.147 102.866 87.207 ;
      RECT MASK 1 33.749 87.2135 33.829 94.4665 ;
      RECT MASK 1 68.807 87.2135 68.887 94.4665 ;
      RECT MASK 1 25.67 87.237 30.62 87.297 ;
      RECT MASK 1 5.984 87.325 12.811 87.365 ;
      RECT MASK 1 13.208 87.325 17.19 87.365 ;
      RECT MASK 1 17.592 87.325 22.239 87.365 ;
      RECT MASK 1 107.479 87.355 128.525 87.395 ;
      RECT MASK 1 36.326 87.399 66.476 87.459 ;
      RECT MASK 1 72.716 87.399 102.866 87.459 ;
      RECT MASK 1 34.36 87.46 35.134 87.5 ;
      RECT MASK 1 67.676 87.46 68.276 87.5 ;
      RECT MASK 1 70.75 87.46 71.524 87.5 ;
      RECT MASK 1 104.058 87.46 104.832 87.5 ;
      RECT MASK 1 22.444 87.49 24.198 87.53 ;
      RECT MASK 1 8.205 87.6335 8.285 90.2665 ;
      RECT MASK 1 12.687 87.6335 12.767 90.2665 ;
      RECT MASK 1 13.253 87.6335 13.333 90.2665 ;
      RECT MASK 1 17.071 87.6335 17.151 90.2665 ;
      RECT MASK 1 17.637 87.6335 17.717 90.2665 ;
      RECT MASK 1 22.119 87.6335 22.199 90.2665 ;
      RECT MASK 1 6.205 87.661 6.869 87.701 ;
      RECT MASK 1 107.504 87.6635 107.584 96.6565 ;
      RECT MASK 1 128.42 87.6635 128.5 96.6565 ;
      RECT MASK 1 8.7735 87.775 12.2035 87.815 ;
      RECT MASK 1 13.8215 87.775 16.5875 87.815 ;
      RECT MASK 1 18.2055 87.775 21.6355 87.815 ;
      RECT MASK 1 2.067 87.81 2.127 88.86 ;
      RECT MASK 1 2.341 87.81 2.401 88.86 ;
      RECT MASK 1 2.615 87.81 2.675 88.86 ;
      RECT MASK 1 2.889 87.81 2.949 88.86 ;
      RECT MASK 1 3.163 87.81 3.223 88.86 ;
      RECT MASK 1 3.437 87.81 3.497 88.86 ;
      RECT MASK 1 3.711 87.81 3.771 88.86 ;
      RECT MASK 1 3.985 87.81 4.045 88.86 ;
      RECT MASK 1 4.259 87.81 4.319 88.86 ;
      RECT MASK 1 4.533 87.81 4.593 88.86 ;
      RECT MASK 1 25.67 87.821 25.941 87.881 ;
      RECT MASK 1 26.211 87.821 30.079 87.881 ;
      RECT MASK 1 30.349 87.821 30.62 87.881 ;
      RECT MASK 1 5.92 87.845 7.154 87.885 ;
      RECT MASK 1 22.444 87.91 24.198 87.95 ;
      RECT MASK 1 72.102 87.922 72.162 88.352 ;
      RECT MASK 1 103.42 87.922 103.48 88.352 ;
      RECT MASK 1 108.242 87.93 108.302 88.98 ;
      RECT MASK 1 108.516 87.93 108.576 88.98 ;
      RECT MASK 1 108.79 87.93 108.85 88.98 ;
      RECT MASK 1 109.064 87.93 109.124 88.98 ;
      RECT MASK 1 109.338 87.93 109.398 88.98 ;
      RECT MASK 1 109.612 87.93 109.672 88.98 ;
      RECT MASK 1 109.886 87.93 109.946 88.98 ;
      RECT MASK 1 110.16 87.93 110.22 88.98 ;
      RECT MASK 1 110.434 87.93 110.494 88.98 ;
      RECT MASK 1 110.708 87.93 110.768 88.98 ;
      RECT MASK 1 110.982 87.93 111.042 88.98 ;
      RECT MASK 1 111.256 87.93 111.316 88.98 ;
      RECT MASK 1 111.53 87.93 111.59 88.98 ;
      RECT MASK 1 111.804 87.93 111.864 88.98 ;
      RECT MASK 1 112.078 87.93 112.138 88.98 ;
      RECT MASK 1 112.352 87.93 112.412 88.98 ;
      RECT MASK 1 112.626 87.93 112.686 88.98 ;
      RECT MASK 1 112.9 87.93 112.96 88.98 ;
      RECT MASK 1 113.174 87.93 113.234 88.98 ;
      RECT MASK 1 113.448 87.93 113.508 88.98 ;
      RECT MASK 1 113.722 87.93 113.782 88.98 ;
      RECT MASK 1 113.996 87.93 114.056 88.98 ;
      RECT MASK 1 114.27 87.93 114.33 88.98 ;
      RECT MASK 1 114.544 87.93 114.604 88.98 ;
      RECT MASK 1 114.818 87.93 114.878 88.98 ;
      RECT MASK 1 115.092 87.93 115.152 88.98 ;
      RECT MASK 1 115.366 87.93 115.426 88.98 ;
      RECT MASK 1 115.64 87.93 115.7 88.98 ;
      RECT MASK 1 115.914 87.93 115.974 88.98 ;
      RECT MASK 1 116.188 87.93 116.248 88.98 ;
      RECT MASK 1 116.462 87.93 116.522 88.98 ;
      RECT MASK 1 116.736 87.93 116.796 88.98 ;
      RECT MASK 1 117.01 87.93 117.07 88.98 ;
      RECT MASK 1 117.284 87.93 117.344 88.98 ;
      RECT MASK 1 117.558 87.93 117.618 88.98 ;
      RECT MASK 1 117.832 87.93 117.892 88.98 ;
      RECT MASK 1 118.106 87.93 118.166 88.98 ;
      RECT MASK 1 118.38 87.93 118.44 88.98 ;
      RECT MASK 1 118.654 87.93 118.714 88.98 ;
      RECT MASK 1 118.928 87.93 118.988 88.98 ;
      RECT MASK 1 119.202 87.93 119.262 88.98 ;
      RECT MASK 1 119.476 87.93 119.536 88.98 ;
      RECT MASK 1 119.75 87.93 119.81 88.98 ;
      RECT MASK 1 120.024 87.93 120.084 88.98 ;
      RECT MASK 1 120.298 87.93 120.358 88.98 ;
      RECT MASK 1 120.572 87.93 120.632 88.98 ;
      RECT MASK 1 120.846 87.93 120.906 88.98 ;
      RECT MASK 1 121.12 87.93 121.18 88.98 ;
      RECT MASK 1 121.394 87.93 121.454 88.98 ;
      RECT MASK 1 121.668 87.93 121.728 88.98 ;
      RECT MASK 1 121.942 87.93 122.002 88.98 ;
      RECT MASK 1 122.216 87.93 122.276 88.98 ;
      RECT MASK 1 122.49 87.93 122.55 88.98 ;
      RECT MASK 1 122.764 87.93 122.824 88.98 ;
      RECT MASK 1 123.038 87.93 123.098 88.98 ;
      RECT MASK 1 123.312 87.93 123.372 88.98 ;
      RECT MASK 1 123.586 87.93 123.646 88.98 ;
      RECT MASK 1 123.86 87.93 123.92 88.98 ;
      RECT MASK 1 124.134 87.93 124.194 88.98 ;
      RECT MASK 1 124.408 87.93 124.468 88.98 ;
      RECT MASK 1 124.682 87.93 124.742 88.98 ;
      RECT MASK 1 124.956 87.93 125.016 88.98 ;
      RECT MASK 1 125.23 87.93 125.29 88.98 ;
      RECT MASK 1 125.504 87.93 125.564 88.98 ;
      RECT MASK 1 125.778 87.93 125.838 88.98 ;
      RECT MASK 1 126.052 87.93 126.112 88.98 ;
      RECT MASK 1 126.326 87.93 126.386 88.98 ;
      RECT MASK 1 126.6 87.93 126.66 88.98 ;
      RECT MASK 1 126.874 87.93 126.934 88.98 ;
      RECT MASK 1 127.148 87.93 127.208 88.98 ;
      RECT MASK 1 127.422 87.93 127.482 88.98 ;
      RECT MASK 1 127.696 87.93 127.756 88.98 ;
      RECT MASK 1 6.492 88.029 6.675 88.069 ;
      RECT MASK 1 36.326 88.047 36.778 88.107 ;
      RECT MASK 1 37.048 88.047 65.754 88.107 ;
      RECT MASK 1 66.024 88.047 66.476 88.107 ;
      RECT MASK 1 72.716 88.047 73.168 88.107 ;
      RECT MASK 1 73.438 88.047 102.144 88.107 ;
      RECT MASK 1 102.414 88.047 102.866 88.107 ;
      RECT MASK 1 34.36 88.07 35.134 88.15 ;
      RECT MASK 1 67.676 88.07 68.276 88.15 ;
      RECT MASK 1 70.75 88.07 71.524 88.15 ;
      RECT MASK 1 104.058 88.07 104.832 88.15 ;
      RECT MASK 1 25.67 88.083 25.938 88.143 ;
      RECT MASK 1 26.212 88.083 30.078 88.143 ;
      RECT MASK 1 30.352 88.083 30.62 88.143 ;
      RECT MASK 1 8.7885 88.0835 8.8685 89.8165 ;
      RECT MASK 1 12.1085 88.0835 12.1885 89.8165 ;
      RECT MASK 1 13.8365 88.0835 13.9165 89.8165 ;
      RECT MASK 1 16.4925 88.0835 16.5725 89.8165 ;
      RECT MASK 1 18.2205 88.0835 18.3005 89.8165 ;
      RECT MASK 1 21.5405 88.0835 21.6205 89.8165 ;
      RECT MASK 1 6.492 88.197 6.675 88.237 ;
      RECT MASK 1 9.1055 88.225 11.8715 88.265 ;
      RECT MASK 1 14.1405 88.225 16.2815 88.265 ;
      RECT MASK 1 18.5375 88.225 21.3035 88.265 ;
      RECT MASK 1 5.949 88.251 6.129 88.291 ;
      RECT MASK 1 6.945 88.251 7.125 88.291 ;
      RECT MASK 1 36.326 88.299 36.778 88.359 ;
      RECT MASK 1 37.048 88.299 65.754 88.359 ;
      RECT MASK 1 66.024 88.299 66.476 88.359 ;
      RECT MASK 1 72.716 88.299 73.168 88.359 ;
      RECT MASK 1 73.438 88.299 102.144 88.359 ;
      RECT MASK 1 102.414 88.299 102.866 88.359 ;
      RECT MASK 1 22.444 88.33 24.198 88.37 ;
      RECT MASK 1 5.949 88.419 6.129 88.459 ;
      RECT MASK 1 6.364 88.419 6.71 88.459 ;
      RECT MASK 1 6.945 88.419 7.125 88.459 ;
      RECT MASK 1 71.997 88.46 72.269 88.52 ;
      RECT MASK 1 103.313 88.46 103.585 88.52 ;
      RECT MASK 1 5.911 88.641 7.163 88.681 ;
      RECT MASK 1 25.67 88.677 30.62 88.737 ;
      RECT MASK 1 9.1305 88.688 9.1905 88.912 ;
      RECT MASK 1 9.4625 88.688 9.5225 88.912 ;
      RECT MASK 1 9.7945 88.688 9.8545 88.912 ;
      RECT MASK 1 10.1265 88.688 10.1865 88.912 ;
      RECT MASK 1 10.4585 88.688 10.5185 88.912 ;
      RECT MASK 1 10.7905 88.688 10.8505 88.912 ;
      RECT MASK 1 11.1225 88.688 11.1825 88.912 ;
      RECT MASK 1 11.4545 88.688 11.5145 88.912 ;
      RECT MASK 1 11.7865 88.688 11.8465 88.912 ;
      RECT MASK 1 14.1785 88.688 14.2385 88.912 ;
      RECT MASK 1 14.5105 88.688 14.5705 88.912 ;
      RECT MASK 1 14.8425 88.688 14.9025 88.912 ;
      RECT MASK 1 15.1745 88.688 15.2345 88.912 ;
      RECT MASK 1 15.5065 88.688 15.5665 88.912 ;
      RECT MASK 1 15.8385 88.688 15.8985 88.912 ;
      RECT MASK 1 16.1705 88.688 16.2305 88.912 ;
      RECT MASK 1 18.7285 88.688 18.7885 88.912 ;
      RECT MASK 1 19.0605 88.688 19.1205 88.912 ;
      RECT MASK 1 19.3925 88.688 19.4525 88.912 ;
      RECT MASK 1 19.7245 88.688 19.7845 88.912 ;
      RECT MASK 1 20.0565 88.688 20.1165 88.912 ;
      RECT MASK 1 20.3885 88.688 20.4485 88.912 ;
      RECT MASK 1 20.7205 88.688 20.7805 88.912 ;
      RECT MASK 1 21.0525 88.688 21.1125 88.912 ;
      RECT MASK 1 22.444 88.75 24.198 88.79 ;
      RECT MASK 1 72.102 88.811 72.162 89.252 ;
      RECT MASK 1 103.42 88.811 103.48 89.252 ;
      RECT MASK 1 34.36 88.91 35.134 88.99 ;
      RECT MASK 1 67.676 88.91 68.276 88.99 ;
      RECT MASK 1 70.75 88.91 71.524 88.99 ;
      RECT MASK 1 104.058 88.91 104.832 88.99 ;
      RECT MASK 1 36.326 88.947 66.476 89.007 ;
      RECT MASK 1 72.716 88.947 102.866 89.007 ;
      RECT MASK 1 6.57 89.01 7.717 89.07 ;
      RECT MASK 1 9.4855 89.17 11.491 89.21 ;
      RECT MASK 1 14.5335 89.17 15.875 89.21 ;
      RECT MASK 1 18.9175 89.17 20.923 89.21 ;
      RECT MASK 1 22.444 89.17 24.198 89.21 ;
      RECT MASK 1 36.326 89.199 66.476 89.259 ;
      RECT MASK 1 72.716 89.199 102.866 89.259 ;
      RECT MASK 1 5.873 89.369 7.201 89.409 ;
      RECT MASK 1 108.242 89.43 108.302 90.48 ;
      RECT MASK 1 108.516 89.43 108.576 90.48 ;
      RECT MASK 1 108.79 89.43 108.85 90.48 ;
      RECT MASK 1 109.064 89.43 109.124 90.48 ;
      RECT MASK 1 109.338 89.43 109.398 90.48 ;
      RECT MASK 1 109.612 89.43 109.672 90.48 ;
      RECT MASK 1 109.886 89.43 109.946 90.48 ;
      RECT MASK 1 110.16 89.43 110.22 90.48 ;
      RECT MASK 1 110.434 89.43 110.494 90.48 ;
      RECT MASK 1 110.708 89.43 110.768 90.48 ;
      RECT MASK 1 110.982 89.43 111.042 90.48 ;
      RECT MASK 1 111.256 89.43 111.316 90.48 ;
      RECT MASK 1 111.53 89.43 111.59 90.48 ;
      RECT MASK 1 111.804 89.43 111.864 90.48 ;
      RECT MASK 1 112.078 89.43 112.138 90.48 ;
      RECT MASK 1 112.352 89.43 112.412 90.48 ;
      RECT MASK 1 112.626 89.43 112.686 90.48 ;
      RECT MASK 1 112.9 89.43 112.96 90.48 ;
      RECT MASK 1 113.174 89.43 113.234 90.48 ;
      RECT MASK 1 113.448 89.43 113.508 90.48 ;
      RECT MASK 1 113.722 89.43 113.782 90.48 ;
      RECT MASK 1 113.996 89.43 114.056 90.48 ;
      RECT MASK 1 114.27 89.43 114.33 90.48 ;
      RECT MASK 1 114.544 89.43 114.604 90.48 ;
      RECT MASK 1 114.818 89.43 114.878 90.48 ;
      RECT MASK 1 115.092 89.43 115.152 90.48 ;
      RECT MASK 1 115.366 89.43 115.426 90.48 ;
      RECT MASK 1 115.64 89.43 115.7 90.48 ;
      RECT MASK 1 115.914 89.43 115.974 90.48 ;
      RECT MASK 1 116.188 89.43 116.248 90.48 ;
      RECT MASK 1 116.462 89.43 116.522 90.48 ;
      RECT MASK 1 116.736 89.43 116.796 90.48 ;
      RECT MASK 1 117.01 89.43 117.07 90.48 ;
      RECT MASK 1 117.284 89.43 117.344 90.48 ;
      RECT MASK 1 117.558 89.43 117.618 90.48 ;
      RECT MASK 1 117.832 89.43 117.892 90.48 ;
      RECT MASK 1 118.106 89.43 118.166 90.48 ;
      RECT MASK 1 118.38 89.43 118.44 90.48 ;
      RECT MASK 1 118.654 89.43 118.714 90.48 ;
      RECT MASK 1 118.928 89.43 118.988 90.48 ;
      RECT MASK 1 119.202 89.43 119.262 90.48 ;
      RECT MASK 1 119.476 89.43 119.536 90.48 ;
      RECT MASK 1 119.75 89.43 119.81 90.48 ;
      RECT MASK 1 120.024 89.43 120.084 90.48 ;
      RECT MASK 1 120.298 89.43 120.358 90.48 ;
      RECT MASK 1 120.572 89.43 120.632 90.48 ;
      RECT MASK 1 120.846 89.43 120.906 90.48 ;
      RECT MASK 1 121.12 89.43 121.18 90.48 ;
      RECT MASK 1 121.394 89.43 121.454 90.48 ;
      RECT MASK 1 121.668 89.43 121.728 90.48 ;
      RECT MASK 1 121.942 89.43 122.002 90.48 ;
      RECT MASK 1 122.216 89.43 122.276 90.48 ;
      RECT MASK 1 122.49 89.43 122.55 90.48 ;
      RECT MASK 1 122.764 89.43 122.824 90.48 ;
      RECT MASK 1 123.038 89.43 123.098 90.48 ;
      RECT MASK 1 123.312 89.43 123.372 90.48 ;
      RECT MASK 1 123.586 89.43 123.646 90.48 ;
      RECT MASK 1 123.86 89.43 123.92 90.48 ;
      RECT MASK 1 124.134 89.43 124.194 90.48 ;
      RECT MASK 1 124.408 89.43 124.468 90.48 ;
      RECT MASK 1 124.682 89.43 124.742 90.48 ;
      RECT MASK 1 124.956 89.43 125.016 90.48 ;
      RECT MASK 1 125.23 89.43 125.29 90.48 ;
      RECT MASK 1 125.504 89.43 125.564 90.48 ;
      RECT MASK 1 125.778 89.43 125.838 90.48 ;
      RECT MASK 1 126.052 89.43 126.112 90.48 ;
      RECT MASK 1 126.326 89.43 126.386 90.48 ;
      RECT MASK 1 126.6 89.43 126.66 90.48 ;
      RECT MASK 1 126.874 89.43 126.934 90.48 ;
      RECT MASK 1 127.148 89.43 127.208 90.48 ;
      RECT MASK 1 127.422 89.43 127.482 90.48 ;
      RECT MASK 1 127.696 89.43 127.756 90.48 ;
      RECT MASK 1 9.1305 89.468 9.1905 89.692 ;
      RECT MASK 1 9.4625 89.468 9.5225 89.692 ;
      RECT MASK 1 9.7945 89.468 9.8545 89.692 ;
      RECT MASK 1 10.1265 89.468 10.1865 89.692 ;
      RECT MASK 1 10.4585 89.468 10.5185 89.692 ;
      RECT MASK 1 10.7905 89.468 10.8505 89.692 ;
      RECT MASK 1 11.1225 89.468 11.1825 89.692 ;
      RECT MASK 1 11.4545 89.468 11.5145 89.692 ;
      RECT MASK 1 11.7865 89.468 11.8465 89.692 ;
      RECT MASK 1 14.1785 89.468 14.2385 89.692 ;
      RECT MASK 1 14.5105 89.468 14.5705 89.692 ;
      RECT MASK 1 14.8425 89.468 14.9025 89.692 ;
      RECT MASK 1 15.1745 89.468 15.2345 89.692 ;
      RECT MASK 1 15.5065 89.468 15.5665 89.692 ;
      RECT MASK 1 15.8385 89.468 15.8985 89.692 ;
      RECT MASK 1 16.1705 89.468 16.2305 89.692 ;
      RECT MASK 1 18.7285 89.468 18.7885 89.692 ;
      RECT MASK 1 19.0605 89.468 19.1205 89.692 ;
      RECT MASK 1 19.3925 89.468 19.4525 89.692 ;
      RECT MASK 1 19.7245 89.468 19.7845 89.692 ;
      RECT MASK 1 20.0565 89.468 20.1165 89.692 ;
      RECT MASK 1 20.3885 89.468 20.4485 89.692 ;
      RECT MASK 1 20.7205 89.468 20.7805 89.692 ;
      RECT MASK 1 21.0525 89.468 21.1125 89.692 ;
      RECT MASK 1 2.067 89.52 2.127 90.57 ;
      RECT MASK 1 2.341 89.52 2.401 90.57 ;
      RECT MASK 1 2.615 89.52 2.675 90.57 ;
      RECT MASK 1 2.889 89.52 2.949 90.57 ;
      RECT MASK 1 3.163 89.52 3.223 90.57 ;
      RECT MASK 1 3.437 89.52 3.497 90.57 ;
      RECT MASK 1 3.711 89.52 3.771 90.57 ;
      RECT MASK 1 3.985 89.52 4.045 90.57 ;
      RECT MASK 1 4.259 89.52 4.319 90.57 ;
      RECT MASK 1 4.533 89.52 4.593 90.57 ;
      RECT MASK 1 25.67 89.577 30.62 89.637 ;
      RECT MASK 1 22.444 89.59 24.198 89.63 ;
      RECT MASK 1 6.364 89.591 6.71 89.631 ;
      RECT MASK 1 5.949 89.627 6.129 89.667 ;
      RECT MASK 1 6.945 89.627 7.125 89.667 ;
      RECT MASK 1 72.102 89.722 72.162 90.152 ;
      RECT MASK 1 103.42 89.722 103.48 90.152 ;
      RECT MASK 1 34.36 89.75 35.134 89.83 ;
      RECT MASK 1 67.676 89.75 68.276 89.83 ;
      RECT MASK 1 70.75 89.75 71.524 89.83 ;
      RECT MASK 1 104.058 89.75 104.832 89.83 ;
      RECT MASK 1 5.949 89.795 6.129 89.835 ;
      RECT MASK 1 6.945 89.795 7.125 89.835 ;
      RECT MASK 1 6.399 89.813 6.582 89.853 ;
      RECT MASK 1 36.326 89.847 36.778 89.907 ;
      RECT MASK 1 37.048 89.847 65.754 89.907 ;
      RECT MASK 1 66.024 89.847 66.476 89.907 ;
      RECT MASK 1 72.716 89.847 73.168 89.907 ;
      RECT MASK 1 73.438 89.847 102.144 89.907 ;
      RECT MASK 1 102.414 89.847 102.866 89.907 ;
      RECT MASK 1 6.399 89.981 6.582 90.021 ;
      RECT MASK 1 22.444 90.01 24.198 90.05 ;
      RECT MASK 1 8.7735 90.085 12.2035 90.125 ;
      RECT MASK 1 13.8215 90.085 16.5875 90.125 ;
      RECT MASK 1 18.2055 90.085 21.6355 90.125 ;
      RECT MASK 1 36.326 90.099 36.778 90.159 ;
      RECT MASK 1 37.048 90.099 65.754 90.159 ;
      RECT MASK 1 66.024 90.099 66.476 90.159 ;
      RECT MASK 1 72.716 90.099 73.168 90.159 ;
      RECT MASK 1 73.438 90.099 102.144 90.159 ;
      RECT MASK 1 102.414 90.099 102.866 90.159 ;
      RECT MASK 1 25.67 90.161 25.941 90.221 ;
      RECT MASK 1 26.211 90.161 30.079 90.221 ;
      RECT MASK 1 30.349 90.161 30.62 90.221 ;
      RECT MASK 1 5.949 90.165 7.125 90.205 ;
      RECT MASK 1 71.997 90.26 72.269 90.32 ;
      RECT MASK 1 103.313 90.26 103.585 90.32 ;
      RECT MASK 1 6.205 90.349 6.869 90.389 ;
      RECT MASK 1 25.67 90.423 25.938 90.483 ;
      RECT MASK 1 26.212 90.423 30.078 90.483 ;
      RECT MASK 1 30.352 90.423 30.62 90.483 ;
      RECT MASK 1 22.444 90.43 24.198 90.47 ;
      RECT MASK 1 8.16 90.535 12.807 90.575 ;
      RECT MASK 1 13.208 90.535 17.19 90.575 ;
      RECT MASK 1 17.592 90.535 22.239 90.575 ;
      RECT MASK 1 34.36 90.59 35.134 90.67 ;
      RECT MASK 1 67.676 90.59 68.276 90.67 ;
      RECT MASK 1 70.75 90.59 71.524 90.67 ;
      RECT MASK 1 104.058 90.59 104.832 90.67 ;
      RECT MASK 1 72.102 90.611 72.162 91.052 ;
      RECT MASK 1 103.42 90.611 103.48 91.052 ;
      RECT MASK 1 5.984 90.745 7.09 90.785 ;
      RECT MASK 1 36.326 90.747 66.476 90.807 ;
      RECT MASK 1 72.716 90.747 102.866 90.807 ;
      RECT MASK 1 22.444 90.85 24.198 90.89 ;
      RECT MASK 1 108.242 90.93 108.302 91.98 ;
      RECT MASK 1 108.516 90.93 108.576 91.98 ;
      RECT MASK 1 108.79 90.93 108.85 91.98 ;
      RECT MASK 1 109.064 90.93 109.124 91.98 ;
      RECT MASK 1 109.338 90.93 109.398 91.98 ;
      RECT MASK 1 109.612 90.93 109.672 91.98 ;
      RECT MASK 1 109.886 90.93 109.946 91.98 ;
      RECT MASK 1 110.16 90.93 110.22 91.98 ;
      RECT MASK 1 110.434 90.93 110.494 91.98 ;
      RECT MASK 1 110.708 90.93 110.768 91.98 ;
      RECT MASK 1 110.982 90.93 111.042 91.98 ;
      RECT MASK 1 111.256 90.93 111.316 91.98 ;
      RECT MASK 1 111.53 90.93 111.59 91.98 ;
      RECT MASK 1 111.804 90.93 111.864 91.98 ;
      RECT MASK 1 112.078 90.93 112.138 91.98 ;
      RECT MASK 1 112.352 90.93 112.412 91.98 ;
      RECT MASK 1 112.626 90.93 112.686 91.98 ;
      RECT MASK 1 112.9 90.93 112.96 91.98 ;
      RECT MASK 1 113.174 90.93 113.234 91.98 ;
      RECT MASK 1 113.448 90.93 113.508 91.98 ;
      RECT MASK 1 113.722 90.93 113.782 91.98 ;
      RECT MASK 1 113.996 90.93 114.056 91.98 ;
      RECT MASK 1 114.27 90.93 114.33 91.98 ;
      RECT MASK 1 114.544 90.93 114.604 91.98 ;
      RECT MASK 1 114.818 90.93 114.878 91.98 ;
      RECT MASK 1 115.092 90.93 115.152 91.98 ;
      RECT MASK 1 115.366 90.93 115.426 91.98 ;
      RECT MASK 1 115.64 90.93 115.7 91.98 ;
      RECT MASK 1 115.914 90.93 115.974 91.98 ;
      RECT MASK 1 116.188 90.93 116.248 91.98 ;
      RECT MASK 1 116.462 90.93 116.522 91.98 ;
      RECT MASK 1 116.736 90.93 116.796 91.98 ;
      RECT MASK 1 117.01 90.93 117.07 91.98 ;
      RECT MASK 1 117.284 90.93 117.344 91.98 ;
      RECT MASK 1 117.558 90.93 117.618 91.98 ;
      RECT MASK 1 117.832 90.93 117.892 91.98 ;
      RECT MASK 1 118.106 90.93 118.166 91.98 ;
      RECT MASK 1 118.38 90.93 118.44 91.98 ;
      RECT MASK 1 118.654 90.93 118.714 91.98 ;
      RECT MASK 1 118.928 90.93 118.988 91.98 ;
      RECT MASK 1 119.202 90.93 119.262 91.98 ;
      RECT MASK 1 119.476 90.93 119.536 91.98 ;
      RECT MASK 1 119.75 90.93 119.81 91.98 ;
      RECT MASK 1 120.024 90.93 120.084 91.98 ;
      RECT MASK 1 120.298 90.93 120.358 91.98 ;
      RECT MASK 1 120.572 90.93 120.632 91.98 ;
      RECT MASK 1 120.846 90.93 120.906 91.98 ;
      RECT MASK 1 121.12 90.93 121.18 91.98 ;
      RECT MASK 1 121.394 90.93 121.454 91.98 ;
      RECT MASK 1 121.668 90.93 121.728 91.98 ;
      RECT MASK 1 121.942 90.93 122.002 91.98 ;
      RECT MASK 1 122.216 90.93 122.276 91.98 ;
      RECT MASK 1 122.49 90.93 122.55 91.98 ;
      RECT MASK 1 122.764 90.93 122.824 91.98 ;
      RECT MASK 1 123.038 90.93 123.098 91.98 ;
      RECT MASK 1 123.312 90.93 123.372 91.98 ;
      RECT MASK 1 123.586 90.93 123.646 91.98 ;
      RECT MASK 1 123.86 90.93 123.92 91.98 ;
      RECT MASK 1 124.134 90.93 124.194 91.98 ;
      RECT MASK 1 124.408 90.93 124.468 91.98 ;
      RECT MASK 1 124.682 90.93 124.742 91.98 ;
      RECT MASK 1 124.956 90.93 125.016 91.98 ;
      RECT MASK 1 125.23 90.93 125.29 91.98 ;
      RECT MASK 1 125.504 90.93 125.564 91.98 ;
      RECT MASK 1 125.778 90.93 125.838 91.98 ;
      RECT MASK 1 126.052 90.93 126.112 91.98 ;
      RECT MASK 1 126.326 90.93 126.386 91.98 ;
      RECT MASK 1 126.6 90.93 126.66 91.98 ;
      RECT MASK 1 126.874 90.93 126.934 91.98 ;
      RECT MASK 1 127.148 90.93 127.208 91.98 ;
      RECT MASK 1 127.422 90.93 127.482 91.98 ;
      RECT MASK 1 127.696 90.93 127.756 91.98 ;
      RECT MASK 1 7.8125 90.985 12.807 91.025 ;
      RECT MASK 1 13.208 90.985 17.19 91.025 ;
      RECT MASK 1 17.592 90.985 22.239 91.025 ;
      RECT MASK 1 36.326 90.999 66.476 91.059 ;
      RECT MASK 1 72.716 90.999 102.866 91.059 ;
      RECT MASK 1 25.67 91.017 30.62 91.077 ;
      RECT MASK 1 6.205 91.171 6.869 91.211 ;
      RECT MASK 1 2.067 91.23 2.127 92.28 ;
      RECT MASK 1 2.341 91.23 2.401 92.28 ;
      RECT MASK 1 2.615 91.23 2.675 92.28 ;
      RECT MASK 1 2.889 91.23 2.949 92.28 ;
      RECT MASK 1 3.163 91.23 3.223 92.28 ;
      RECT MASK 1 3.437 91.23 3.497 92.28 ;
      RECT MASK 1 3.711 91.23 3.771 92.28 ;
      RECT MASK 1 3.985 91.23 4.045 92.28 ;
      RECT MASK 1 4.259 91.23 4.319 92.28 ;
      RECT MASK 1 4.533 91.23 4.593 92.28 ;
      RECT MASK 1 22.444 91.27 24.198 91.31 ;
      RECT MASK 1 7.873 91.2935 7.953 93.9265 ;
      RECT MASK 1 12.687 91.2935 12.767 93.9265 ;
      RECT MASK 1 13.253 91.2935 13.333 93.9265 ;
      RECT MASK 1 17.071 91.2935 17.151 93.9265 ;
      RECT MASK 1 17.637 91.2935 17.717 93.9265 ;
      RECT MASK 1 22.119 91.2935 22.199 93.9265 ;
      RECT MASK 1 5.949 91.355 7.125 91.395 ;
      RECT MASK 1 34.36 91.43 35.134 91.51 ;
      RECT MASK 1 67.676 91.43 68.276 91.51 ;
      RECT MASK 1 70.75 91.43 71.524 91.51 ;
      RECT MASK 1 104.058 91.43 104.832 91.51 ;
      RECT MASK 1 8.446 91.435 11.876 91.475 ;
      RECT MASK 1 13.8215 91.435 16.5875 91.475 ;
      RECT MASK 1 18.2055 91.435 21.6355 91.475 ;
      RECT MASK 1 72.102 91.522 72.162 91.952 ;
      RECT MASK 1 103.42 91.522 103.48 91.952 ;
      RECT MASK 1 6.492 91.539 6.675 91.579 ;
      RECT MASK 1 25.188 91.63 31.092 91.67 ;
      RECT MASK 1 36.326 91.647 36.778 91.707 ;
      RECT MASK 1 37.048 91.647 65.754 91.707 ;
      RECT MASK 1 66.024 91.647 66.476 91.707 ;
      RECT MASK 1 72.716 91.647 73.168 91.707 ;
      RECT MASK 1 73.438 91.647 102.144 91.707 ;
      RECT MASK 1 102.414 91.647 102.866 91.707 ;
      RECT MASK 1 22.444 91.69 24.198 91.73 ;
      RECT MASK 1 6.492 91.707 6.675 91.747 ;
      RECT MASK 1 5.949 91.725 6.129 91.765 ;
      RECT MASK 1 6.945 91.725 7.125 91.765 ;
      RECT MASK 1 8.461 91.7435 8.541 93.4765 ;
      RECT MASK 1 11.781 91.7435 11.861 93.4765 ;
      RECT MASK 1 13.8365 91.7435 13.9165 93.4765 ;
      RECT MASK 1 16.4925 91.7435 16.5725 93.4765 ;
      RECT MASK 1 18.2205 91.7435 18.3005 93.4765 ;
      RECT MASK 1 21.5405 91.7435 21.6205 93.4765 ;
      RECT MASK 1 8.803 91.868 8.863 92.092 ;
      RECT MASK 1 9.135 91.868 9.195 92.092 ;
      RECT MASK 1 9.467 91.868 9.527 92.092 ;
      RECT MASK 1 9.799 91.868 9.859 92.092 ;
      RECT MASK 1 10.131 91.868 10.191 92.092 ;
      RECT MASK 1 10.463 91.868 10.523 92.092 ;
      RECT MASK 1 10.795 91.868 10.855 92.092 ;
      RECT MASK 1 11.127 91.868 11.187 92.092 ;
      RECT MASK 1 11.459 91.868 11.519 92.092 ;
      RECT MASK 1 14.1785 91.868 14.2385 92.092 ;
      RECT MASK 1 14.5105 91.868 14.5705 92.092 ;
      RECT MASK 1 14.8425 91.868 14.9025 92.092 ;
      RECT MASK 1 15.1745 91.868 15.2345 92.092 ;
      RECT MASK 1 15.5065 91.868 15.5665 92.092 ;
      RECT MASK 1 15.8385 91.868 15.8985 92.092 ;
      RECT MASK 1 16.1705 91.868 16.2305 92.092 ;
      RECT MASK 1 18.7285 91.868 18.7885 92.092 ;
      RECT MASK 1 19.0605 91.868 19.1205 92.092 ;
      RECT MASK 1 19.3925 91.868 19.4525 92.092 ;
      RECT MASK 1 19.7245 91.868 19.7845 92.092 ;
      RECT MASK 1 20.0565 91.868 20.1165 92.092 ;
      RECT MASK 1 20.3885 91.868 20.4485 92.092 ;
      RECT MASK 1 20.7205 91.868 20.7805 92.092 ;
      RECT MASK 1 21.0525 91.868 21.1125 92.092 ;
      RECT MASK 1 5.949 91.893 6.129 91.933 ;
      RECT MASK 1 6.945 91.893 7.125 91.933 ;
      RECT MASK 1 36.326 91.899 36.778 91.959 ;
      RECT MASK 1 37.048 91.899 65.754 91.959 ;
      RECT MASK 1 66.024 91.899 66.476 91.959 ;
      RECT MASK 1 72.716 91.899 73.168 91.959 ;
      RECT MASK 1 73.438 91.899 102.144 91.959 ;
      RECT MASK 1 102.414 91.899 102.866 91.959 ;
      RECT MASK 1 6.364 91.929 6.71 91.969 ;
      RECT MASK 1 71.997 92.06 72.269 92.12 ;
      RECT MASK 1 103.313 92.06 103.585 92.12 ;
      RECT MASK 1 22.444 92.11 24.198 92.15 ;
      RECT MASK 1 5.873 92.151 7.201 92.191 ;
      RECT MASK 1 34.36 92.27 35.134 92.35 ;
      RECT MASK 1 67.676 92.27 68.276 92.35 ;
      RECT MASK 1 70.75 92.27 71.524 92.35 ;
      RECT MASK 1 104.058 92.27 104.832 92.35 ;
      RECT MASK 1 9.158 92.35 11.1635 92.39 ;
      RECT MASK 1 14.5335 92.35 15.875 92.39 ;
      RECT MASK 1 18.9175 92.35 20.923 92.39 ;
      RECT MASK 1 72.102 92.411 72.162 92.852 ;
      RECT MASK 1 103.42 92.411 103.48 92.852 ;
      RECT MASK 1 108.242 92.43 108.302 93.48 ;
      RECT MASK 1 108.516 92.43 108.576 93.48 ;
      RECT MASK 1 108.79 92.43 108.85 93.48 ;
      RECT MASK 1 109.064 92.43 109.124 93.48 ;
      RECT MASK 1 109.338 92.43 109.398 93.48 ;
      RECT MASK 1 109.612 92.43 109.672 93.48 ;
      RECT MASK 1 109.886 92.43 109.946 93.48 ;
      RECT MASK 1 110.16 92.43 110.22 93.48 ;
      RECT MASK 1 110.434 92.43 110.494 93.48 ;
      RECT MASK 1 110.708 92.43 110.768 93.48 ;
      RECT MASK 1 110.982 92.43 111.042 93.48 ;
      RECT MASK 1 111.256 92.43 111.316 93.48 ;
      RECT MASK 1 111.53 92.43 111.59 93.48 ;
      RECT MASK 1 111.804 92.43 111.864 93.48 ;
      RECT MASK 1 112.078 92.43 112.138 93.48 ;
      RECT MASK 1 112.352 92.43 112.412 93.48 ;
      RECT MASK 1 112.626 92.43 112.686 93.48 ;
      RECT MASK 1 112.9 92.43 112.96 93.48 ;
      RECT MASK 1 113.174 92.43 113.234 93.48 ;
      RECT MASK 1 113.448 92.43 113.508 93.48 ;
      RECT MASK 1 113.722 92.43 113.782 93.48 ;
      RECT MASK 1 113.996 92.43 114.056 93.48 ;
      RECT MASK 1 114.27 92.43 114.33 93.48 ;
      RECT MASK 1 114.544 92.43 114.604 93.48 ;
      RECT MASK 1 114.818 92.43 114.878 93.48 ;
      RECT MASK 1 115.092 92.43 115.152 93.48 ;
      RECT MASK 1 115.366 92.43 115.426 93.48 ;
      RECT MASK 1 115.64 92.43 115.7 93.48 ;
      RECT MASK 1 115.914 92.43 115.974 93.48 ;
      RECT MASK 1 116.188 92.43 116.248 93.48 ;
      RECT MASK 1 116.462 92.43 116.522 93.48 ;
      RECT MASK 1 116.736 92.43 116.796 93.48 ;
      RECT MASK 1 117.01 92.43 117.07 93.48 ;
      RECT MASK 1 117.284 92.43 117.344 93.48 ;
      RECT MASK 1 117.558 92.43 117.618 93.48 ;
      RECT MASK 1 117.832 92.43 117.892 93.48 ;
      RECT MASK 1 118.106 92.43 118.166 93.48 ;
      RECT MASK 1 118.38 92.43 118.44 93.48 ;
      RECT MASK 1 118.654 92.43 118.714 93.48 ;
      RECT MASK 1 118.928 92.43 118.988 93.48 ;
      RECT MASK 1 119.202 92.43 119.262 93.48 ;
      RECT MASK 1 119.476 92.43 119.536 93.48 ;
      RECT MASK 1 119.75 92.43 119.81 93.48 ;
      RECT MASK 1 120.024 92.43 120.084 93.48 ;
      RECT MASK 1 120.298 92.43 120.358 93.48 ;
      RECT MASK 1 120.572 92.43 120.632 93.48 ;
      RECT MASK 1 120.846 92.43 120.906 93.48 ;
      RECT MASK 1 121.12 92.43 121.18 93.48 ;
      RECT MASK 1 121.394 92.43 121.454 93.48 ;
      RECT MASK 1 121.668 92.43 121.728 93.48 ;
      RECT MASK 1 121.942 92.43 122.002 93.48 ;
      RECT MASK 1 122.216 92.43 122.276 93.48 ;
      RECT MASK 1 122.49 92.43 122.55 93.48 ;
      RECT MASK 1 122.764 92.43 122.824 93.48 ;
      RECT MASK 1 123.038 92.43 123.098 93.48 ;
      RECT MASK 1 123.312 92.43 123.372 93.48 ;
      RECT MASK 1 123.586 92.43 123.646 93.48 ;
      RECT MASK 1 123.86 92.43 123.92 93.48 ;
      RECT MASK 1 124.134 92.43 124.194 93.48 ;
      RECT MASK 1 124.408 92.43 124.468 93.48 ;
      RECT MASK 1 124.682 92.43 124.742 93.48 ;
      RECT MASK 1 124.956 92.43 125.016 93.48 ;
      RECT MASK 1 125.23 92.43 125.29 93.48 ;
      RECT MASK 1 125.504 92.43 125.564 93.48 ;
      RECT MASK 1 125.778 92.43 125.838 93.48 ;
      RECT MASK 1 126.052 92.43 126.112 93.48 ;
      RECT MASK 1 126.326 92.43 126.386 93.48 ;
      RECT MASK 1 126.6 92.43 126.66 93.48 ;
      RECT MASK 1 126.874 92.43 126.934 93.48 ;
      RECT MASK 1 127.148 92.43 127.208 93.48 ;
      RECT MASK 1 127.422 92.43 127.482 93.48 ;
      RECT MASK 1 127.696 92.43 127.756 93.48 ;
      RECT MASK 1 22.444 92.53 24.198 92.57 ;
      RECT MASK 1 36.326 92.547 66.476 92.607 ;
      RECT MASK 1 72.716 92.547 102.866 92.607 ;
      RECT MASK 1 8.803 92.648 8.863 92.872 ;
      RECT MASK 1 9.135 92.648 9.195 92.872 ;
      RECT MASK 1 9.467 92.648 9.527 92.872 ;
      RECT MASK 1 9.799 92.648 9.859 92.872 ;
      RECT MASK 1 10.131 92.648 10.191 92.872 ;
      RECT MASK 1 10.463 92.648 10.523 92.872 ;
      RECT MASK 1 10.795 92.648 10.855 92.872 ;
      RECT MASK 1 11.127 92.648 11.187 92.872 ;
      RECT MASK 1 11.459 92.648 11.519 92.872 ;
      RECT MASK 1 14.1785 92.648 14.2385 92.872 ;
      RECT MASK 1 14.5105 92.648 14.5705 92.872 ;
      RECT MASK 1 14.8425 92.648 14.9025 92.872 ;
      RECT MASK 1 15.1745 92.648 15.2345 92.872 ;
      RECT MASK 1 15.5065 92.648 15.5665 92.872 ;
      RECT MASK 1 15.8385 92.648 15.8985 92.872 ;
      RECT MASK 1 16.1705 92.648 16.2305 92.872 ;
      RECT MASK 1 18.7285 92.648 18.7885 92.872 ;
      RECT MASK 1 19.0605 92.648 19.1205 92.872 ;
      RECT MASK 1 19.3925 92.648 19.4525 92.872 ;
      RECT MASK 1 19.7245 92.648 19.7845 92.872 ;
      RECT MASK 1 20.0565 92.648 20.1165 92.872 ;
      RECT MASK 1 20.3885 92.648 20.4485 92.872 ;
      RECT MASK 1 20.7205 92.648 20.7805 92.872 ;
      RECT MASK 1 21.0525 92.648 21.1125 92.872 ;
      RECT MASK 1 36.326 92.799 66.476 92.859 ;
      RECT MASK 1 72.716 92.799 102.866 92.859 ;
      RECT MASK 1 5.911 92.879 7.163 92.919 ;
      RECT MASK 1 2.067 92.94 2.127 93.99 ;
      RECT MASK 1 2.341 92.94 2.401 93.99 ;
      RECT MASK 1 2.615 92.94 2.675 93.99 ;
      RECT MASK 1 2.889 92.94 2.949 93.99 ;
      RECT MASK 1 3.163 92.94 3.223 93.99 ;
      RECT MASK 1 3.437 92.94 3.497 93.99 ;
      RECT MASK 1 3.711 92.94 3.771 93.99 ;
      RECT MASK 1 3.985 92.94 4.045 93.99 ;
      RECT MASK 1 4.259 92.94 4.319 93.99 ;
      RECT MASK 1 4.533 92.94 4.593 93.99 ;
      RECT MASK 1 22.444 92.95 24.198 92.99 ;
      RECT MASK 1 5.949 93.101 6.129 93.141 ;
      RECT MASK 1 6.364 93.101 6.71 93.141 ;
      RECT MASK 1 6.945 93.101 7.125 93.141 ;
      RECT MASK 1 34.36 93.11 35.134 93.19 ;
      RECT MASK 1 67.676 93.11 68.276 93.19 ;
      RECT MASK 1 70.75 93.11 71.524 93.19 ;
      RECT MASK 1 104.058 93.11 104.832 93.19 ;
      RECT MASK 1 5.949 93.269 6.129 93.309 ;
      RECT MASK 1 6.945 93.269 7.125 93.309 ;
      RECT MASK 1 8.778 93.295 11.544 93.335 ;
      RECT MASK 1 14.1405 93.295 16.2815 93.335 ;
      RECT MASK 1 18.5375 93.295 21.3035 93.335 ;
      RECT MASK 1 72.102 93.322 72.162 93.752 ;
      RECT MASK 1 103.42 93.322 103.48 93.752 ;
      RECT MASK 1 6.399 93.323 6.582 93.363 ;
      RECT MASK 1 22.444 93.37 24.198 93.41 ;
      RECT MASK 1 36.326 93.447 36.778 93.507 ;
      RECT MASK 1 37.048 93.447 65.754 93.507 ;
      RECT MASK 1 66.024 93.447 66.476 93.507 ;
      RECT MASK 1 72.716 93.447 73.168 93.507 ;
      RECT MASK 1 73.438 93.447 102.144 93.507 ;
      RECT MASK 1 102.414 93.447 102.866 93.507 ;
      RECT MASK 1 6.399 93.491 6.582 93.531 ;
      RECT MASK 1 5.92 93.675 7.154 93.715 ;
      RECT MASK 1 36.326 93.699 36.778 93.759 ;
      RECT MASK 1 37.048 93.699 65.754 93.759 ;
      RECT MASK 1 66.024 93.699 66.476 93.759 ;
      RECT MASK 1 72.716 93.699 73.168 93.759 ;
      RECT MASK 1 73.438 93.699 102.144 93.759 ;
      RECT MASK 1 102.414 93.699 102.866 93.759 ;
      RECT MASK 1 8.446 93.745 11.876 93.785 ;
      RECT MASK 1 13.8215 93.745 16.5875 93.785 ;
      RECT MASK 1 18.2055 93.745 21.6355 93.785 ;
      RECT MASK 1 22.444 93.79 24.198 93.83 ;
      RECT MASK 1 6.205 93.859 7.732 93.899 ;
      RECT MASK 1 71.997 93.86 72.269 93.92 ;
      RECT MASK 1 103.313 93.86 103.585 93.92 ;
      RECT MASK 1 108.242 93.93 108.302 94.98 ;
      RECT MASK 1 108.516 93.93 108.576 94.98 ;
      RECT MASK 1 108.79 93.93 108.85 94.98 ;
      RECT MASK 1 109.064 93.93 109.124 94.98 ;
      RECT MASK 1 109.338 93.93 109.398 94.98 ;
      RECT MASK 1 109.612 93.93 109.672 94.98 ;
      RECT MASK 1 109.886 93.93 109.946 94.98 ;
      RECT MASK 1 110.16 93.93 110.22 94.98 ;
      RECT MASK 1 110.434 93.93 110.494 94.98 ;
      RECT MASK 1 110.708 93.93 110.768 94.98 ;
      RECT MASK 1 110.982 93.93 111.042 94.98 ;
      RECT MASK 1 111.256 93.93 111.316 94.98 ;
      RECT MASK 1 111.53 93.93 111.59 94.98 ;
      RECT MASK 1 111.804 93.93 111.864 94.98 ;
      RECT MASK 1 112.078 93.93 112.138 94.98 ;
      RECT MASK 1 112.352 93.93 112.412 94.98 ;
      RECT MASK 1 112.626 93.93 112.686 94.98 ;
      RECT MASK 1 112.9 93.93 112.96 94.98 ;
      RECT MASK 1 113.174 93.93 113.234 94.98 ;
      RECT MASK 1 113.448 93.93 113.508 94.98 ;
      RECT MASK 1 113.722 93.93 113.782 94.98 ;
      RECT MASK 1 113.996 93.93 114.056 94.98 ;
      RECT MASK 1 114.27 93.93 114.33 94.98 ;
      RECT MASK 1 114.544 93.93 114.604 94.98 ;
      RECT MASK 1 114.818 93.93 114.878 94.98 ;
      RECT MASK 1 115.092 93.93 115.152 94.98 ;
      RECT MASK 1 115.366 93.93 115.426 94.98 ;
      RECT MASK 1 115.64 93.93 115.7 94.98 ;
      RECT MASK 1 115.914 93.93 115.974 94.98 ;
      RECT MASK 1 116.188 93.93 116.248 94.98 ;
      RECT MASK 1 116.462 93.93 116.522 94.98 ;
      RECT MASK 1 116.736 93.93 116.796 94.98 ;
      RECT MASK 1 117.01 93.93 117.07 94.98 ;
      RECT MASK 1 117.284 93.93 117.344 94.98 ;
      RECT MASK 1 117.558 93.93 117.618 94.98 ;
      RECT MASK 1 117.832 93.93 117.892 94.98 ;
      RECT MASK 1 118.106 93.93 118.166 94.98 ;
      RECT MASK 1 118.38 93.93 118.44 94.98 ;
      RECT MASK 1 118.654 93.93 118.714 94.98 ;
      RECT MASK 1 118.928 93.93 118.988 94.98 ;
      RECT MASK 1 119.202 93.93 119.262 94.98 ;
      RECT MASK 1 119.476 93.93 119.536 94.98 ;
      RECT MASK 1 119.75 93.93 119.81 94.98 ;
      RECT MASK 1 120.024 93.93 120.084 94.98 ;
      RECT MASK 1 120.298 93.93 120.358 94.98 ;
      RECT MASK 1 120.572 93.93 120.632 94.98 ;
      RECT MASK 1 120.846 93.93 120.906 94.98 ;
      RECT MASK 1 121.12 93.93 121.18 94.98 ;
      RECT MASK 1 121.394 93.93 121.454 94.98 ;
      RECT MASK 1 121.668 93.93 121.728 94.98 ;
      RECT MASK 1 121.942 93.93 122.002 94.98 ;
      RECT MASK 1 122.216 93.93 122.276 94.98 ;
      RECT MASK 1 122.49 93.93 122.55 94.98 ;
      RECT MASK 1 122.764 93.93 122.824 94.98 ;
      RECT MASK 1 123.038 93.93 123.098 94.98 ;
      RECT MASK 1 123.312 93.93 123.372 94.98 ;
      RECT MASK 1 123.586 93.93 123.646 94.98 ;
      RECT MASK 1 123.86 93.93 123.92 94.98 ;
      RECT MASK 1 124.134 93.93 124.194 94.98 ;
      RECT MASK 1 124.408 93.93 124.468 94.98 ;
      RECT MASK 1 124.682 93.93 124.742 94.98 ;
      RECT MASK 1 124.956 93.93 125.016 94.98 ;
      RECT MASK 1 125.23 93.93 125.29 94.98 ;
      RECT MASK 1 125.504 93.93 125.564 94.98 ;
      RECT MASK 1 125.778 93.93 125.838 94.98 ;
      RECT MASK 1 126.052 93.93 126.112 94.98 ;
      RECT MASK 1 126.326 93.93 126.386 94.98 ;
      RECT MASK 1 126.6 93.93 126.66 94.98 ;
      RECT MASK 1 126.874 93.93 126.934 94.98 ;
      RECT MASK 1 127.148 93.93 127.208 94.98 ;
      RECT MASK 1 127.422 93.93 127.482 94.98 ;
      RECT MASK 1 127.696 93.93 127.756 94.98 ;
      RECT MASK 1 34.36 93.95 35.134 94.03 ;
      RECT MASK 1 67.676 93.95 68.276 94.03 ;
      RECT MASK 1 70.75 93.95 71.524 94.03 ;
      RECT MASK 1 104.058 93.95 104.832 94.03 ;
      RECT MASK 1 5.984 94.195 12.811 94.235 ;
      RECT MASK 1 13.208 94.195 17.19 94.235 ;
      RECT MASK 1 17.592 94.195 22.239 94.235 ;
      RECT MASK 1 22.444 94.21 24.198 94.25 ;
      RECT MASK 1 72.102 94.227 72.162 94.652 ;
      RECT MASK 1 103.42 94.227 103.48 94.652 ;
      RECT MASK 1 36.326 94.347 66.476 94.407 ;
      RECT MASK 1 72.716 94.347 102.866 94.407 ;
      RECT MASK 1 36.326 94.599 66.476 94.659 ;
      RECT MASK 1 72.716 94.599 102.866 94.659 ;
      RECT MASK 1 22.444 94.63 31.502 94.67 ;
      RECT MASK 1 2.067 94.65 2.127 95.7 ;
      RECT MASK 1 2.341 94.65 2.401 95.7 ;
      RECT MASK 1 2.615 94.65 2.675 95.7 ;
      RECT MASK 1 2.889 94.65 2.949 95.7 ;
      RECT MASK 1 3.163 94.65 3.223 95.7 ;
      RECT MASK 1 3.437 94.65 3.497 95.7 ;
      RECT MASK 1 3.711 94.65 3.771 95.7 ;
      RECT MASK 1 3.985 94.65 4.045 95.7 ;
      RECT MASK 1 4.259 94.65 4.319 95.7 ;
      RECT MASK 1 4.533 94.65 4.593 95.7 ;
      RECT MASK 1 33.739 94.735 35.338 94.775 ;
      RECT MASK 1 67.467 94.735 68.897 94.775 ;
      RECT MASK 1 70.129 94.825 71.728 94.865 ;
      RECT MASK 1 103.854 94.825 105.453 94.865 ;
      RECT MASK 1 22.444 95.05 31.502 95.09 ;
      RECT MASK 1 35.702 95.051 35.782 95.269 ;
      RECT MASK 1 67.02 95.051 67.1 95.269 ;
      RECT MASK 1 72.092 95.051 72.172 95.269 ;
      RECT MASK 1 103.41 95.051 103.49 95.269 ;
      RECT MASK 1 36.1535 95.111 66.6485 95.211 ;
      RECT MASK 1 72.5435 95.111 103.0385 95.211 ;
      RECT MASK 1 33.407 95.185 35.338 95.225 ;
      RECT MASK 1 67.467 95.185 69.229 95.225 ;
      RECT MASK 1 69.797 95.275 71.728 95.315 ;
      RECT MASK 1 103.854 95.275 105.785 95.315 ;
      RECT MASK 1 108.242 95.43 108.302 96.48 ;
      RECT MASK 1 108.516 95.43 108.576 96.48 ;
      RECT MASK 1 108.79 95.43 108.85 96.48 ;
      RECT MASK 1 109.064 95.43 109.124 96.48 ;
      RECT MASK 1 109.338 95.43 109.398 96.48 ;
      RECT MASK 1 109.612 95.43 109.672 96.48 ;
      RECT MASK 1 109.886 95.43 109.946 96.48 ;
      RECT MASK 1 110.16 95.43 110.22 96.48 ;
      RECT MASK 1 110.434 95.43 110.494 96.48 ;
      RECT MASK 1 110.708 95.43 110.768 96.48 ;
      RECT MASK 1 110.982 95.43 111.042 96.48 ;
      RECT MASK 1 111.256 95.43 111.316 96.48 ;
      RECT MASK 1 111.53 95.43 111.59 96.48 ;
      RECT MASK 1 111.804 95.43 111.864 96.48 ;
      RECT MASK 1 112.078 95.43 112.138 96.48 ;
      RECT MASK 1 112.352 95.43 112.412 96.48 ;
      RECT MASK 1 112.626 95.43 112.686 96.48 ;
      RECT MASK 1 112.9 95.43 112.96 96.48 ;
      RECT MASK 1 113.174 95.43 113.234 96.48 ;
      RECT MASK 1 113.448 95.43 113.508 96.48 ;
      RECT MASK 1 113.722 95.43 113.782 96.48 ;
      RECT MASK 1 113.996 95.43 114.056 96.48 ;
      RECT MASK 1 114.27 95.43 114.33 96.48 ;
      RECT MASK 1 114.544 95.43 114.604 96.48 ;
      RECT MASK 1 114.818 95.43 114.878 96.48 ;
      RECT MASK 1 115.092 95.43 115.152 96.48 ;
      RECT MASK 1 115.366 95.43 115.426 96.48 ;
      RECT MASK 1 115.64 95.43 115.7 96.48 ;
      RECT MASK 1 115.914 95.43 115.974 96.48 ;
      RECT MASK 1 116.188 95.43 116.248 96.48 ;
      RECT MASK 1 116.462 95.43 116.522 96.48 ;
      RECT MASK 1 116.736 95.43 116.796 96.48 ;
      RECT MASK 1 117.01 95.43 117.07 96.48 ;
      RECT MASK 1 117.284 95.43 117.344 96.48 ;
      RECT MASK 1 117.558 95.43 117.618 96.48 ;
      RECT MASK 1 117.832 95.43 117.892 96.48 ;
      RECT MASK 1 118.106 95.43 118.166 96.48 ;
      RECT MASK 1 118.38 95.43 118.44 96.48 ;
      RECT MASK 1 118.654 95.43 118.714 96.48 ;
      RECT MASK 1 118.928 95.43 118.988 96.48 ;
      RECT MASK 1 119.202 95.43 119.262 96.48 ;
      RECT MASK 1 119.476 95.43 119.536 96.48 ;
      RECT MASK 1 119.75 95.43 119.81 96.48 ;
      RECT MASK 1 120.024 95.43 120.084 96.48 ;
      RECT MASK 1 120.298 95.43 120.358 96.48 ;
      RECT MASK 1 120.572 95.43 120.632 96.48 ;
      RECT MASK 1 120.846 95.43 120.906 96.48 ;
      RECT MASK 1 121.12 95.43 121.18 96.48 ;
      RECT MASK 1 121.394 95.43 121.454 96.48 ;
      RECT MASK 1 121.668 95.43 121.728 96.48 ;
      RECT MASK 1 121.942 95.43 122.002 96.48 ;
      RECT MASK 1 122.216 95.43 122.276 96.48 ;
      RECT MASK 1 122.49 95.43 122.55 96.48 ;
      RECT MASK 1 122.764 95.43 122.824 96.48 ;
      RECT MASK 1 123.038 95.43 123.098 96.48 ;
      RECT MASK 1 123.312 95.43 123.372 96.48 ;
      RECT MASK 1 123.586 95.43 123.646 96.48 ;
      RECT MASK 1 123.86 95.43 123.92 96.48 ;
      RECT MASK 1 124.134 95.43 124.194 96.48 ;
      RECT MASK 1 124.408 95.43 124.468 96.48 ;
      RECT MASK 1 124.682 95.43 124.742 96.48 ;
      RECT MASK 1 124.956 95.43 125.016 96.48 ;
      RECT MASK 1 125.23 95.43 125.29 96.48 ;
      RECT MASK 1 125.504 95.43 125.564 96.48 ;
      RECT MASK 1 125.778 95.43 125.838 96.48 ;
      RECT MASK 1 126.052 95.43 126.112 96.48 ;
      RECT MASK 1 126.326 95.43 126.386 96.48 ;
      RECT MASK 1 126.6 95.43 126.66 96.48 ;
      RECT MASK 1 126.874 95.43 126.934 96.48 ;
      RECT MASK 1 127.148 95.43 127.208 96.48 ;
      RECT MASK 1 127.422 95.43 127.482 96.48 ;
      RECT MASK 1 127.696 95.43 127.756 96.48 ;
      RECT MASK 1 22.444 95.47 31.502 95.51 ;
      RECT MASK 1 22.444 95.89 36.656 95.93 ;
      RECT MASK 1 1.248 96.235 5.362 96.275 ;
      RECT MASK 1 22.444 96.31 36.656 96.35 ;
      RECT MASK 1 107.479 96.925 128.525 96.965 ;
      RECT MASK 1 1.439 97.375 44.397 97.415 ;
      RECT MASK 1 44.831 97.375 87.789 97.415 ;
      RECT MASK 1 88.223 97.375 128.525 97.415 ;
      RECT MASK 1 1.464 97.6835 1.544 107.5765 ;
      RECT MASK 1 44.292 97.6835 44.372 107.5765 ;
      RECT MASK 1 44.856 97.6835 44.936 107.5765 ;
      RECT MASK 1 87.684 97.6835 87.764 107.5765 ;
      RECT MASK 1 88.248 97.6835 88.328 107.5765 ;
      RECT MASK 1 128.42 97.6835 128.5 107.5765 ;
      RECT MASK 1 2.201 97.83 2.261 98.88 ;
      RECT MASK 1 2.475 97.83 2.535 98.88 ;
      RECT MASK 1 2.749 97.83 2.809 98.88 ;
      RECT MASK 1 3.023 97.83 3.083 98.88 ;
      RECT MASK 1 3.297 97.83 3.357 98.88 ;
      RECT MASK 1 3.571 97.83 3.631 98.88 ;
      RECT MASK 1 3.845 97.83 3.905 98.88 ;
      RECT MASK 1 4.119 97.83 4.179 98.88 ;
      RECT MASK 1 4.393 97.83 4.453 98.88 ;
      RECT MASK 1 4.667 97.83 4.727 98.88 ;
      RECT MASK 1 4.941 97.83 5.001 98.88 ;
      RECT MASK 1 5.215 97.83 5.275 98.88 ;
      RECT MASK 1 5.489 97.83 5.549 98.88 ;
      RECT MASK 1 5.763 97.83 5.823 98.88 ;
      RECT MASK 1 6.037 97.83 6.097 98.88 ;
      RECT MASK 1 6.311 97.83 6.371 98.88 ;
      RECT MASK 1 6.585 97.83 6.645 98.88 ;
      RECT MASK 1 6.859 97.83 6.919 98.88 ;
      RECT MASK 1 7.133 97.83 7.193 98.88 ;
      RECT MASK 1 7.407 97.83 7.467 98.88 ;
      RECT MASK 1 7.681 97.83 7.741 98.88 ;
      RECT MASK 1 7.955 97.83 8.015 98.88 ;
      RECT MASK 1 8.229 97.83 8.289 98.88 ;
      RECT MASK 1 8.503 97.83 8.563 98.88 ;
      RECT MASK 1 8.777 97.83 8.837 98.88 ;
      RECT MASK 1 9.051 97.83 9.111 98.88 ;
      RECT MASK 1 9.325 97.83 9.385 98.88 ;
      RECT MASK 1 9.599 97.83 9.659 98.88 ;
      RECT MASK 1 9.873 97.83 9.933 98.88 ;
      RECT MASK 1 10.147 97.83 10.207 98.88 ;
      RECT MASK 1 10.421 97.83 10.481 98.88 ;
      RECT MASK 1 10.695 97.83 10.755 98.88 ;
      RECT MASK 1 10.969 97.83 11.029 98.88 ;
      RECT MASK 1 11.243 97.83 11.303 98.88 ;
      RECT MASK 1 11.517 97.83 11.577 98.88 ;
      RECT MASK 1 11.791 97.83 11.851 98.88 ;
      RECT MASK 1 12.065 97.83 12.125 98.88 ;
      RECT MASK 1 12.339 97.83 12.399 98.88 ;
      RECT MASK 1 12.613 97.83 12.673 98.88 ;
      RECT MASK 1 12.887 97.83 12.947 98.88 ;
      RECT MASK 1 13.161 97.83 13.221 98.88 ;
      RECT MASK 1 13.435 97.83 13.495 98.88 ;
      RECT MASK 1 13.709 97.83 13.769 98.88 ;
      RECT MASK 1 13.983 97.83 14.043 98.88 ;
      RECT MASK 1 14.257 97.83 14.317 98.88 ;
      RECT MASK 1 14.531 97.83 14.591 98.88 ;
      RECT MASK 1 14.805 97.83 14.865 98.88 ;
      RECT MASK 1 15.079 97.83 15.139 98.88 ;
      RECT MASK 1 15.353 97.83 15.413 98.88 ;
      RECT MASK 1 15.627 97.83 15.687 98.88 ;
      RECT MASK 1 15.901 97.83 15.961 98.88 ;
      RECT MASK 1 16.175 97.83 16.235 98.88 ;
      RECT MASK 1 16.449 97.83 16.509 98.88 ;
      RECT MASK 1 16.723 97.83 16.783 98.88 ;
      RECT MASK 1 16.997 97.83 17.057 98.88 ;
      RECT MASK 1 17.271 97.83 17.331 98.88 ;
      RECT MASK 1 17.545 97.83 17.605 98.88 ;
      RECT MASK 1 17.819 97.83 17.879 98.88 ;
      RECT MASK 1 18.093 97.83 18.153 98.88 ;
      RECT MASK 1 18.367 97.83 18.427 98.88 ;
      RECT MASK 1 18.641 97.83 18.701 98.88 ;
      RECT MASK 1 18.915 97.83 18.975 98.88 ;
      RECT MASK 1 19.189 97.83 19.249 98.88 ;
      RECT MASK 1 19.463 97.83 19.523 98.88 ;
      RECT MASK 1 19.737 97.83 19.797 98.88 ;
      RECT MASK 1 20.011 97.83 20.071 98.88 ;
      RECT MASK 1 20.285 97.83 20.345 98.88 ;
      RECT MASK 1 20.559 97.83 20.619 98.88 ;
      RECT MASK 1 20.833 97.83 20.893 98.88 ;
      RECT MASK 1 21.107 97.83 21.167 98.88 ;
      RECT MASK 1 21.381 97.83 21.441 98.88 ;
      RECT MASK 1 21.655 97.83 21.715 98.88 ;
      RECT MASK 1 21.929 97.83 21.989 98.88 ;
      RECT MASK 1 22.203 97.83 22.263 98.88 ;
      RECT MASK 1 22.477 97.83 22.537 98.88 ;
      RECT MASK 1 22.751 97.83 22.811 98.88 ;
      RECT MASK 1 23.025 97.83 23.085 98.88 ;
      RECT MASK 1 23.299 97.83 23.359 98.88 ;
      RECT MASK 1 23.573 97.83 23.633 98.88 ;
      RECT MASK 1 23.847 97.83 23.907 98.88 ;
      RECT MASK 1 24.121 97.83 24.181 98.88 ;
      RECT MASK 1 24.395 97.83 24.455 98.88 ;
      RECT MASK 1 24.669 97.83 24.729 98.88 ;
      RECT MASK 1 24.943 97.83 25.003 98.88 ;
      RECT MASK 1 25.217 97.83 25.277 98.88 ;
      RECT MASK 1 25.491 97.83 25.551 98.88 ;
      RECT MASK 1 25.765 97.83 25.825 98.88 ;
      RECT MASK 1 26.039 97.83 26.099 98.88 ;
      RECT MASK 1 26.313 97.83 26.373 98.88 ;
      RECT MASK 1 26.587 97.83 26.647 98.88 ;
      RECT MASK 1 26.861 97.83 26.921 98.88 ;
      RECT MASK 1 27.135 97.83 27.195 98.88 ;
      RECT MASK 1 27.409 97.83 27.469 98.88 ;
      RECT MASK 1 27.683 97.83 27.743 98.88 ;
      RECT MASK 1 27.957 97.83 28.017 98.88 ;
      RECT MASK 1 28.231 97.83 28.291 98.88 ;
      RECT MASK 1 28.505 97.83 28.565 98.88 ;
      RECT MASK 1 28.779 97.83 28.839 98.88 ;
      RECT MASK 1 29.053 97.83 29.113 98.88 ;
      RECT MASK 1 29.327 97.83 29.387 98.88 ;
      RECT MASK 1 29.601 97.83 29.661 98.88 ;
      RECT MASK 1 29.875 97.83 29.935 98.88 ;
      RECT MASK 1 30.149 97.83 30.209 98.88 ;
      RECT MASK 1 30.423 97.83 30.483 98.88 ;
      RECT MASK 1 30.697 97.83 30.757 98.88 ;
      RECT MASK 1 30.971 97.83 31.031 98.88 ;
      RECT MASK 1 31.245 97.83 31.305 98.88 ;
      RECT MASK 1 31.519 97.83 31.579 98.88 ;
      RECT MASK 1 31.793 97.83 31.853 98.88 ;
      RECT MASK 1 32.067 97.83 32.127 98.88 ;
      RECT MASK 1 32.341 97.83 32.401 98.88 ;
      RECT MASK 1 32.615 97.83 32.675 98.88 ;
      RECT MASK 1 32.889 97.83 32.949 98.88 ;
      RECT MASK 1 33.163 97.83 33.223 98.88 ;
      RECT MASK 1 33.437 97.83 33.497 98.88 ;
      RECT MASK 1 33.711 97.83 33.771 98.88 ;
      RECT MASK 1 33.985 97.83 34.045 98.88 ;
      RECT MASK 1 34.259 97.83 34.319 98.88 ;
      RECT MASK 1 34.533 97.83 34.593 98.88 ;
      RECT MASK 1 34.807 97.83 34.867 98.88 ;
      RECT MASK 1 35.081 97.83 35.141 98.88 ;
      RECT MASK 1 35.355 97.83 35.415 98.88 ;
      RECT MASK 1 35.629 97.83 35.689 98.88 ;
      RECT MASK 1 35.903 97.83 35.963 98.88 ;
      RECT MASK 1 36.177 97.83 36.237 98.88 ;
      RECT MASK 1 36.451 97.83 36.511 98.88 ;
      RECT MASK 1 36.725 97.83 36.785 98.88 ;
      RECT MASK 1 36.999 97.83 37.059 98.88 ;
      RECT MASK 1 37.273 97.83 37.333 98.88 ;
      RECT MASK 1 37.547 97.83 37.607 98.88 ;
      RECT MASK 1 37.821 97.83 37.881 98.88 ;
      RECT MASK 1 38.095 97.83 38.155 98.88 ;
      RECT MASK 1 38.369 97.83 38.429 98.88 ;
      RECT MASK 1 38.643 97.83 38.703 98.88 ;
      RECT MASK 1 38.917 97.83 38.977 98.88 ;
      RECT MASK 1 39.191 97.83 39.251 98.88 ;
      RECT MASK 1 39.465 97.83 39.525 98.88 ;
      RECT MASK 1 39.739 97.83 39.799 98.88 ;
      RECT MASK 1 40.013 97.83 40.073 98.88 ;
      RECT MASK 1 40.287 97.83 40.347 98.88 ;
      RECT MASK 1 40.561 97.83 40.621 98.88 ;
      RECT MASK 1 40.835 97.83 40.895 98.88 ;
      RECT MASK 1 41.109 97.83 41.169 98.88 ;
      RECT MASK 1 41.383 97.83 41.443 98.88 ;
      RECT MASK 1 41.657 97.83 41.717 98.88 ;
      RECT MASK 1 41.931 97.83 41.991 98.88 ;
      RECT MASK 1 42.205 97.83 42.265 98.88 ;
      RECT MASK 1 42.479 97.83 42.539 98.88 ;
      RECT MASK 1 42.753 97.83 42.813 98.88 ;
      RECT MASK 1 43.027 97.83 43.087 98.88 ;
      RECT MASK 1 43.301 97.83 43.361 98.88 ;
      RECT MASK 1 43.575 97.83 43.635 98.88 ;
      RECT MASK 1 45.593 97.83 45.653 98.88 ;
      RECT MASK 1 45.867 97.83 45.927 98.88 ;
      RECT MASK 1 46.141 97.83 46.201 98.88 ;
      RECT MASK 1 46.415 97.83 46.475 98.88 ;
      RECT MASK 1 46.689 97.83 46.749 98.88 ;
      RECT MASK 1 46.963 97.83 47.023 98.88 ;
      RECT MASK 1 47.237 97.83 47.297 98.88 ;
      RECT MASK 1 47.511 97.83 47.571 98.88 ;
      RECT MASK 1 47.785 97.83 47.845 98.88 ;
      RECT MASK 1 48.059 97.83 48.119 98.88 ;
      RECT MASK 1 48.333 97.83 48.393 98.88 ;
      RECT MASK 1 48.607 97.83 48.667 98.88 ;
      RECT MASK 1 48.881 97.83 48.941 98.88 ;
      RECT MASK 1 49.155 97.83 49.215 98.88 ;
      RECT MASK 1 49.429 97.83 49.489 98.88 ;
      RECT MASK 1 49.703 97.83 49.763 98.88 ;
      RECT MASK 1 49.977 97.83 50.037 98.88 ;
      RECT MASK 1 50.251 97.83 50.311 98.88 ;
      RECT MASK 1 50.525 97.83 50.585 98.88 ;
      RECT MASK 1 50.799 97.83 50.859 98.88 ;
      RECT MASK 1 51.073 97.83 51.133 98.88 ;
      RECT MASK 1 51.347 97.83 51.407 98.88 ;
      RECT MASK 1 51.621 97.83 51.681 98.88 ;
      RECT MASK 1 51.895 97.83 51.955 98.88 ;
      RECT MASK 1 52.169 97.83 52.229 98.88 ;
      RECT MASK 1 52.443 97.83 52.503 98.88 ;
      RECT MASK 1 52.717 97.83 52.777 98.88 ;
      RECT MASK 1 52.991 97.83 53.051 98.88 ;
      RECT MASK 1 53.265 97.83 53.325 98.88 ;
      RECT MASK 1 53.539 97.83 53.599 98.88 ;
      RECT MASK 1 53.813 97.83 53.873 98.88 ;
      RECT MASK 1 54.087 97.83 54.147 98.88 ;
      RECT MASK 1 54.361 97.83 54.421 98.88 ;
      RECT MASK 1 54.635 97.83 54.695 98.88 ;
      RECT MASK 1 54.909 97.83 54.969 98.88 ;
      RECT MASK 1 55.183 97.83 55.243 98.88 ;
      RECT MASK 1 55.457 97.83 55.517 98.88 ;
      RECT MASK 1 55.731 97.83 55.791 98.88 ;
      RECT MASK 1 56.005 97.83 56.065 98.88 ;
      RECT MASK 1 56.279 97.83 56.339 98.88 ;
      RECT MASK 1 56.553 97.83 56.613 98.88 ;
      RECT MASK 1 56.827 97.83 56.887 98.88 ;
      RECT MASK 1 57.101 97.83 57.161 98.88 ;
      RECT MASK 1 57.375 97.83 57.435 98.88 ;
      RECT MASK 1 57.649 97.83 57.709 98.88 ;
      RECT MASK 1 57.923 97.83 57.983 98.88 ;
      RECT MASK 1 58.197 97.83 58.257 98.88 ;
      RECT MASK 1 58.471 97.83 58.531 98.88 ;
      RECT MASK 1 58.745 97.83 58.805 98.88 ;
      RECT MASK 1 59.019 97.83 59.079 98.88 ;
      RECT MASK 1 59.293 97.83 59.353 98.88 ;
      RECT MASK 1 59.567 97.83 59.627 98.88 ;
      RECT MASK 1 59.841 97.83 59.901 98.88 ;
      RECT MASK 1 60.115 97.83 60.175 98.88 ;
      RECT MASK 1 60.389 97.83 60.449 98.88 ;
      RECT MASK 1 60.663 97.83 60.723 98.88 ;
      RECT MASK 1 60.937 97.83 60.997 98.88 ;
      RECT MASK 1 61.211 97.83 61.271 98.88 ;
      RECT MASK 1 61.485 97.83 61.545 98.88 ;
      RECT MASK 1 61.759 97.83 61.819 98.88 ;
      RECT MASK 1 62.033 97.83 62.093 98.88 ;
      RECT MASK 1 62.307 97.83 62.367 98.88 ;
      RECT MASK 1 62.581 97.83 62.641 98.88 ;
      RECT MASK 1 62.855 97.83 62.915 98.88 ;
      RECT MASK 1 63.129 97.83 63.189 98.88 ;
      RECT MASK 1 63.403 97.83 63.463 98.88 ;
      RECT MASK 1 63.677 97.83 63.737 98.88 ;
      RECT MASK 1 63.951 97.83 64.011 98.88 ;
      RECT MASK 1 64.225 97.83 64.285 98.88 ;
      RECT MASK 1 64.499 97.83 64.559 98.88 ;
      RECT MASK 1 64.773 97.83 64.833 98.88 ;
      RECT MASK 1 65.047 97.83 65.107 98.88 ;
      RECT MASK 1 65.321 97.83 65.381 98.88 ;
      RECT MASK 1 65.595 97.83 65.655 98.88 ;
      RECT MASK 1 65.869 97.83 65.929 98.88 ;
      RECT MASK 1 66.143 97.83 66.203 98.88 ;
      RECT MASK 1 66.417 97.83 66.477 98.88 ;
      RECT MASK 1 66.691 97.83 66.751 98.88 ;
      RECT MASK 1 66.965 97.83 67.025 98.88 ;
      RECT MASK 1 67.239 97.83 67.299 98.88 ;
      RECT MASK 1 67.513 97.83 67.573 98.88 ;
      RECT MASK 1 67.787 97.83 67.847 98.88 ;
      RECT MASK 1 68.061 97.83 68.121 98.88 ;
      RECT MASK 1 68.335 97.83 68.395 98.88 ;
      RECT MASK 1 68.609 97.83 68.669 98.88 ;
      RECT MASK 1 68.883 97.83 68.943 98.88 ;
      RECT MASK 1 69.157 97.83 69.217 98.88 ;
      RECT MASK 1 69.431 97.83 69.491 98.88 ;
      RECT MASK 1 69.705 97.83 69.765 98.88 ;
      RECT MASK 1 69.979 97.83 70.039 98.88 ;
      RECT MASK 1 70.253 97.83 70.313 98.88 ;
      RECT MASK 1 70.527 97.83 70.587 98.88 ;
      RECT MASK 1 70.801 97.83 70.861 98.88 ;
      RECT MASK 1 71.075 97.83 71.135 98.88 ;
      RECT MASK 1 71.349 97.83 71.409 98.88 ;
      RECT MASK 1 71.623 97.83 71.683 98.88 ;
      RECT MASK 1 71.897 97.83 71.957 98.88 ;
      RECT MASK 1 72.171 97.83 72.231 98.88 ;
      RECT MASK 1 72.445 97.83 72.505 98.88 ;
      RECT MASK 1 72.719 97.83 72.779 98.88 ;
      RECT MASK 1 72.993 97.83 73.053 98.88 ;
      RECT MASK 1 73.267 97.83 73.327 98.88 ;
      RECT MASK 1 73.541 97.83 73.601 98.88 ;
      RECT MASK 1 73.815 97.83 73.875 98.88 ;
      RECT MASK 1 74.089 97.83 74.149 98.88 ;
      RECT MASK 1 74.363 97.83 74.423 98.88 ;
      RECT MASK 1 74.637 97.83 74.697 98.88 ;
      RECT MASK 1 74.911 97.83 74.971 98.88 ;
      RECT MASK 1 75.185 97.83 75.245 98.88 ;
      RECT MASK 1 75.459 97.83 75.519 98.88 ;
      RECT MASK 1 75.733 97.83 75.793 98.88 ;
      RECT MASK 1 76.007 97.83 76.067 98.88 ;
      RECT MASK 1 76.281 97.83 76.341 98.88 ;
      RECT MASK 1 76.555 97.83 76.615 98.88 ;
      RECT MASK 1 76.829 97.83 76.889 98.88 ;
      RECT MASK 1 77.103 97.83 77.163 98.88 ;
      RECT MASK 1 77.377 97.83 77.437 98.88 ;
      RECT MASK 1 77.651 97.83 77.711 98.88 ;
      RECT MASK 1 77.925 97.83 77.985 98.88 ;
      RECT MASK 1 78.199 97.83 78.259 98.88 ;
      RECT MASK 1 78.473 97.83 78.533 98.88 ;
      RECT MASK 1 78.747 97.83 78.807 98.88 ;
      RECT MASK 1 79.021 97.83 79.081 98.88 ;
      RECT MASK 1 79.295 97.83 79.355 98.88 ;
      RECT MASK 1 79.569 97.83 79.629 98.88 ;
      RECT MASK 1 79.843 97.83 79.903 98.88 ;
      RECT MASK 1 80.117 97.83 80.177 98.88 ;
      RECT MASK 1 80.391 97.83 80.451 98.88 ;
      RECT MASK 1 80.665 97.83 80.725 98.88 ;
      RECT MASK 1 80.939 97.83 80.999 98.88 ;
      RECT MASK 1 81.213 97.83 81.273 98.88 ;
      RECT MASK 1 81.487 97.83 81.547 98.88 ;
      RECT MASK 1 81.761 97.83 81.821 98.88 ;
      RECT MASK 1 82.035 97.83 82.095 98.88 ;
      RECT MASK 1 82.309 97.83 82.369 98.88 ;
      RECT MASK 1 82.583 97.83 82.643 98.88 ;
      RECT MASK 1 82.857 97.83 82.917 98.88 ;
      RECT MASK 1 83.131 97.83 83.191 98.88 ;
      RECT MASK 1 83.405 97.83 83.465 98.88 ;
      RECT MASK 1 83.679 97.83 83.739 98.88 ;
      RECT MASK 1 83.953 97.83 84.013 98.88 ;
      RECT MASK 1 84.227 97.83 84.287 98.88 ;
      RECT MASK 1 84.501 97.83 84.561 98.88 ;
      RECT MASK 1 84.775 97.83 84.835 98.88 ;
      RECT MASK 1 85.049 97.83 85.109 98.88 ;
      RECT MASK 1 85.323 97.83 85.383 98.88 ;
      RECT MASK 1 85.597 97.83 85.657 98.88 ;
      RECT MASK 1 85.871 97.83 85.931 98.88 ;
      RECT MASK 1 86.145 97.83 86.205 98.88 ;
      RECT MASK 1 86.419 97.83 86.479 98.88 ;
      RECT MASK 1 86.693 97.83 86.753 98.88 ;
      RECT MASK 1 86.967 97.83 87.027 98.88 ;
      RECT MASK 1 88.952 97.83 89.012 98.88 ;
      RECT MASK 1 89.226 97.83 89.286 98.88 ;
      RECT MASK 1 89.5 97.83 89.56 98.88 ;
      RECT MASK 1 89.774 97.83 89.834 98.88 ;
      RECT MASK 1 90.048 97.83 90.108 98.88 ;
      RECT MASK 1 90.322 97.83 90.382 98.88 ;
      RECT MASK 1 90.596 97.83 90.656 98.88 ;
      RECT MASK 1 90.87 97.83 90.93 98.88 ;
      RECT MASK 1 91.144 97.83 91.204 98.88 ;
      RECT MASK 1 91.418 97.83 91.478 98.88 ;
      RECT MASK 1 91.692 97.83 91.752 98.88 ;
      RECT MASK 1 91.966 97.83 92.026 98.88 ;
      RECT MASK 1 92.24 97.83 92.3 98.88 ;
      RECT MASK 1 92.514 97.83 92.574 98.88 ;
      RECT MASK 1 92.788 97.83 92.848 98.88 ;
      RECT MASK 1 93.062 97.83 93.122 98.88 ;
      RECT MASK 1 93.336 97.83 93.396 98.88 ;
      RECT MASK 1 93.61 97.83 93.67 98.88 ;
      RECT MASK 1 93.884 97.83 93.944 98.88 ;
      RECT MASK 1 94.158 97.83 94.218 98.88 ;
      RECT MASK 1 94.432 97.83 94.492 98.88 ;
      RECT MASK 1 94.706 97.83 94.766 98.88 ;
      RECT MASK 1 94.98 97.83 95.04 98.88 ;
      RECT MASK 1 95.254 97.83 95.314 98.88 ;
      RECT MASK 1 95.528 97.83 95.588 98.88 ;
      RECT MASK 1 95.802 97.83 95.862 98.88 ;
      RECT MASK 1 96.076 97.83 96.136 98.88 ;
      RECT MASK 1 96.35 97.83 96.41 98.88 ;
      RECT MASK 1 96.624 97.83 96.684 98.88 ;
      RECT MASK 1 96.898 97.83 96.958 98.88 ;
      RECT MASK 1 97.172 97.83 97.232 98.88 ;
      RECT MASK 1 97.446 97.83 97.506 98.88 ;
      RECT MASK 1 97.72 97.83 97.78 98.88 ;
      RECT MASK 1 97.994 97.83 98.054 98.88 ;
      RECT MASK 1 98.268 97.83 98.328 98.88 ;
      RECT MASK 1 98.542 97.83 98.602 98.88 ;
      RECT MASK 1 98.816 97.83 98.876 98.88 ;
      RECT MASK 1 99.09 97.83 99.15 98.88 ;
      RECT MASK 1 99.364 97.83 99.424 98.88 ;
      RECT MASK 1 99.638 97.83 99.698 98.88 ;
      RECT MASK 1 99.912 97.83 99.972 98.88 ;
      RECT MASK 1 100.186 97.83 100.246 98.88 ;
      RECT MASK 1 100.46 97.83 100.52 98.88 ;
      RECT MASK 1 100.734 97.83 100.794 98.88 ;
      RECT MASK 1 101.008 97.83 101.068 98.88 ;
      RECT MASK 1 101.282 97.83 101.342 98.88 ;
      RECT MASK 1 101.556 97.83 101.616 98.88 ;
      RECT MASK 1 101.83 97.83 101.89 98.88 ;
      RECT MASK 1 102.104 97.83 102.164 98.88 ;
      RECT MASK 1 102.378 97.83 102.438 98.88 ;
      RECT MASK 1 102.652 97.83 102.712 98.88 ;
      RECT MASK 1 102.926 97.83 102.986 98.88 ;
      RECT MASK 1 103.2 97.83 103.26 98.88 ;
      RECT MASK 1 103.474 97.83 103.534 98.88 ;
      RECT MASK 1 103.748 97.83 103.808 98.88 ;
      RECT MASK 1 104.022 97.83 104.082 98.88 ;
      RECT MASK 1 104.296 97.83 104.356 98.88 ;
      RECT MASK 1 104.57 97.83 104.63 98.88 ;
      RECT MASK 1 104.844 97.83 104.904 98.88 ;
      RECT MASK 1 105.118 97.83 105.178 98.88 ;
      RECT MASK 1 105.392 97.83 105.452 98.88 ;
      RECT MASK 1 105.666 97.83 105.726 98.88 ;
      RECT MASK 1 105.94 97.83 106 98.88 ;
      RECT MASK 1 106.214 97.83 106.274 98.88 ;
      RECT MASK 1 106.488 97.83 106.548 98.88 ;
      RECT MASK 1 106.762 97.83 106.822 98.88 ;
      RECT MASK 1 107.036 97.83 107.096 98.88 ;
      RECT MASK 1 107.31 97.83 107.37 98.88 ;
      RECT MASK 1 107.584 97.83 107.644 98.88 ;
      RECT MASK 1 107.858 97.83 107.918 98.88 ;
      RECT MASK 1 108.132 97.83 108.192 98.88 ;
      RECT MASK 1 108.406 97.83 108.466 98.88 ;
      RECT MASK 1 108.68 97.83 108.74 98.88 ;
      RECT MASK 1 108.954 97.83 109.014 98.88 ;
      RECT MASK 1 109.228 97.83 109.288 98.88 ;
      RECT MASK 1 109.502 97.83 109.562 98.88 ;
      RECT MASK 1 109.776 97.83 109.836 98.88 ;
      RECT MASK 1 110.05 97.83 110.11 98.88 ;
      RECT MASK 1 110.324 97.83 110.384 98.88 ;
      RECT MASK 1 110.598 97.83 110.658 98.88 ;
      RECT MASK 1 110.872 97.83 110.932 98.88 ;
      RECT MASK 1 111.146 97.83 111.206 98.88 ;
      RECT MASK 1 111.42 97.83 111.48 98.88 ;
      RECT MASK 1 111.694 97.83 111.754 98.88 ;
      RECT MASK 1 111.968 97.83 112.028 98.88 ;
      RECT MASK 1 112.242 97.83 112.302 98.88 ;
      RECT MASK 1 112.516 97.83 112.576 98.88 ;
      RECT MASK 1 112.79 97.83 112.85 98.88 ;
      RECT MASK 1 113.064 97.83 113.124 98.88 ;
      RECT MASK 1 113.338 97.83 113.398 98.88 ;
      RECT MASK 1 113.612 97.83 113.672 98.88 ;
      RECT MASK 1 113.886 97.83 113.946 98.88 ;
      RECT MASK 1 114.16 97.83 114.22 98.88 ;
      RECT MASK 1 114.434 97.83 114.494 98.88 ;
      RECT MASK 1 114.708 97.83 114.768 98.88 ;
      RECT MASK 1 114.982 97.83 115.042 98.88 ;
      RECT MASK 1 115.256 97.83 115.316 98.88 ;
      RECT MASK 1 115.53 97.83 115.59 98.88 ;
      RECT MASK 1 115.804 97.83 115.864 98.88 ;
      RECT MASK 1 116.078 97.83 116.138 98.88 ;
      RECT MASK 1 116.352 97.83 116.412 98.88 ;
      RECT MASK 1 116.626 97.83 116.686 98.88 ;
      RECT MASK 1 116.9 97.83 116.96 98.88 ;
      RECT MASK 1 117.174 97.83 117.234 98.88 ;
      RECT MASK 1 117.448 97.83 117.508 98.88 ;
      RECT MASK 1 117.722 97.83 117.782 98.88 ;
      RECT MASK 1 117.996 97.83 118.056 98.88 ;
      RECT MASK 1 118.27 97.83 118.33 98.88 ;
      RECT MASK 1 118.544 97.83 118.604 98.88 ;
      RECT MASK 1 118.818 97.83 118.878 98.88 ;
      RECT MASK 1 119.092 97.83 119.152 98.88 ;
      RECT MASK 1 119.366 97.83 119.426 98.88 ;
      RECT MASK 1 119.64 97.83 119.7 98.88 ;
      RECT MASK 1 119.914 97.83 119.974 98.88 ;
      RECT MASK 1 120.188 97.83 120.248 98.88 ;
      RECT MASK 1 120.462 97.83 120.522 98.88 ;
      RECT MASK 1 120.736 97.83 120.796 98.88 ;
      RECT MASK 1 121.01 97.83 121.07 98.88 ;
      RECT MASK 1 121.284 97.83 121.344 98.88 ;
      RECT MASK 1 121.558 97.83 121.618 98.88 ;
      RECT MASK 1 121.832 97.83 121.892 98.88 ;
      RECT MASK 1 122.106 97.83 122.166 98.88 ;
      RECT MASK 1 122.38 97.83 122.44 98.88 ;
      RECT MASK 1 122.654 97.83 122.714 98.88 ;
      RECT MASK 1 122.928 97.83 122.988 98.88 ;
      RECT MASK 1 123.202 97.83 123.262 98.88 ;
      RECT MASK 1 123.476 97.83 123.536 98.88 ;
      RECT MASK 1 123.75 97.83 123.81 98.88 ;
      RECT MASK 1 124.024 97.83 124.084 98.88 ;
      RECT MASK 1 124.298 97.83 124.358 98.88 ;
      RECT MASK 1 124.572 97.83 124.632 98.88 ;
      RECT MASK 1 124.846 97.83 124.906 98.88 ;
      RECT MASK 1 125.12 97.83 125.18 98.88 ;
      RECT MASK 1 125.394 97.83 125.454 98.88 ;
      RECT MASK 1 125.668 97.83 125.728 98.88 ;
      RECT MASK 1 125.942 97.83 126.002 98.88 ;
      RECT MASK 1 126.216 97.83 126.276 98.88 ;
      RECT MASK 1 126.49 97.83 126.55 98.88 ;
      RECT MASK 1 126.764 97.83 126.824 98.88 ;
      RECT MASK 1 127.038 97.83 127.098 98.88 ;
      RECT MASK 1 127.312 97.83 127.372 98.88 ;
      RECT MASK 1 127.586 97.83 127.646 98.88 ;
      RECT MASK 1 2.201 99.54 2.261 100.59 ;
      RECT MASK 1 2.475 99.54 2.535 100.59 ;
      RECT MASK 1 2.749 99.54 2.809 100.59 ;
      RECT MASK 1 3.023 99.54 3.083 100.59 ;
      RECT MASK 1 3.297 99.54 3.357 100.59 ;
      RECT MASK 1 3.571 99.54 3.631 100.59 ;
      RECT MASK 1 3.845 99.54 3.905 100.59 ;
      RECT MASK 1 4.119 99.54 4.179 100.59 ;
      RECT MASK 1 4.393 99.54 4.453 100.59 ;
      RECT MASK 1 4.667 99.54 4.727 100.59 ;
      RECT MASK 1 4.941 99.54 5.001 100.59 ;
      RECT MASK 1 5.215 99.54 5.275 100.59 ;
      RECT MASK 1 5.489 99.54 5.549 100.59 ;
      RECT MASK 1 5.763 99.54 5.823 100.59 ;
      RECT MASK 1 6.037 99.54 6.097 100.59 ;
      RECT MASK 1 6.311 99.54 6.371 100.59 ;
      RECT MASK 1 6.585 99.54 6.645 100.59 ;
      RECT MASK 1 6.859 99.54 6.919 100.59 ;
      RECT MASK 1 7.133 99.54 7.193 100.59 ;
      RECT MASK 1 7.407 99.54 7.467 100.59 ;
      RECT MASK 1 7.681 99.54 7.741 100.59 ;
      RECT MASK 1 7.955 99.54 8.015 100.59 ;
      RECT MASK 1 8.229 99.54 8.289 100.59 ;
      RECT MASK 1 8.503 99.54 8.563 100.59 ;
      RECT MASK 1 8.777 99.54 8.837 100.59 ;
      RECT MASK 1 9.051 99.54 9.111 100.59 ;
      RECT MASK 1 9.325 99.54 9.385 100.59 ;
      RECT MASK 1 9.599 99.54 9.659 100.59 ;
      RECT MASK 1 9.873 99.54 9.933 100.59 ;
      RECT MASK 1 10.147 99.54 10.207 100.59 ;
      RECT MASK 1 10.421 99.54 10.481 100.59 ;
      RECT MASK 1 10.695 99.54 10.755 100.59 ;
      RECT MASK 1 10.969 99.54 11.029 100.59 ;
      RECT MASK 1 11.243 99.54 11.303 100.59 ;
      RECT MASK 1 11.517 99.54 11.577 100.59 ;
      RECT MASK 1 11.791 99.54 11.851 100.59 ;
      RECT MASK 1 12.065 99.54 12.125 100.59 ;
      RECT MASK 1 12.339 99.54 12.399 100.59 ;
      RECT MASK 1 12.613 99.54 12.673 100.59 ;
      RECT MASK 1 12.887 99.54 12.947 100.59 ;
      RECT MASK 1 13.161 99.54 13.221 100.59 ;
      RECT MASK 1 13.435 99.54 13.495 100.59 ;
      RECT MASK 1 13.709 99.54 13.769 100.59 ;
      RECT MASK 1 13.983 99.54 14.043 100.59 ;
      RECT MASK 1 14.257 99.54 14.317 100.59 ;
      RECT MASK 1 14.531 99.54 14.591 100.59 ;
      RECT MASK 1 14.805 99.54 14.865 100.59 ;
      RECT MASK 1 15.079 99.54 15.139 100.59 ;
      RECT MASK 1 15.353 99.54 15.413 100.59 ;
      RECT MASK 1 15.627 99.54 15.687 100.59 ;
      RECT MASK 1 15.901 99.54 15.961 100.59 ;
      RECT MASK 1 16.175 99.54 16.235 100.59 ;
      RECT MASK 1 16.449 99.54 16.509 100.59 ;
      RECT MASK 1 16.723 99.54 16.783 100.59 ;
      RECT MASK 1 16.997 99.54 17.057 100.59 ;
      RECT MASK 1 17.271 99.54 17.331 100.59 ;
      RECT MASK 1 17.545 99.54 17.605 100.59 ;
      RECT MASK 1 17.819 99.54 17.879 100.59 ;
      RECT MASK 1 18.093 99.54 18.153 100.59 ;
      RECT MASK 1 18.367 99.54 18.427 100.59 ;
      RECT MASK 1 18.641 99.54 18.701 100.59 ;
      RECT MASK 1 18.915 99.54 18.975 100.59 ;
      RECT MASK 1 19.189 99.54 19.249 100.59 ;
      RECT MASK 1 19.463 99.54 19.523 100.59 ;
      RECT MASK 1 19.737 99.54 19.797 100.59 ;
      RECT MASK 1 20.011 99.54 20.071 100.59 ;
      RECT MASK 1 20.285 99.54 20.345 100.59 ;
      RECT MASK 1 20.559 99.54 20.619 100.59 ;
      RECT MASK 1 20.833 99.54 20.893 100.59 ;
      RECT MASK 1 21.107 99.54 21.167 100.59 ;
      RECT MASK 1 21.381 99.54 21.441 100.59 ;
      RECT MASK 1 21.655 99.54 21.715 100.59 ;
      RECT MASK 1 21.929 99.54 21.989 100.59 ;
      RECT MASK 1 22.203 99.54 22.263 100.59 ;
      RECT MASK 1 22.477 99.54 22.537 100.59 ;
      RECT MASK 1 22.751 99.54 22.811 100.59 ;
      RECT MASK 1 23.025 99.54 23.085 100.59 ;
      RECT MASK 1 23.299 99.54 23.359 100.59 ;
      RECT MASK 1 23.573 99.54 23.633 100.59 ;
      RECT MASK 1 23.847 99.54 23.907 100.59 ;
      RECT MASK 1 24.121 99.54 24.181 100.59 ;
      RECT MASK 1 24.395 99.54 24.455 100.59 ;
      RECT MASK 1 24.669 99.54 24.729 100.59 ;
      RECT MASK 1 24.943 99.54 25.003 100.59 ;
      RECT MASK 1 25.217 99.54 25.277 100.59 ;
      RECT MASK 1 25.491 99.54 25.551 100.59 ;
      RECT MASK 1 25.765 99.54 25.825 100.59 ;
      RECT MASK 1 26.039 99.54 26.099 100.59 ;
      RECT MASK 1 26.313 99.54 26.373 100.59 ;
      RECT MASK 1 26.587 99.54 26.647 100.59 ;
      RECT MASK 1 26.861 99.54 26.921 100.59 ;
      RECT MASK 1 27.135 99.54 27.195 100.59 ;
      RECT MASK 1 27.409 99.54 27.469 100.59 ;
      RECT MASK 1 27.683 99.54 27.743 100.59 ;
      RECT MASK 1 27.957 99.54 28.017 100.59 ;
      RECT MASK 1 28.231 99.54 28.291 100.59 ;
      RECT MASK 1 28.505 99.54 28.565 100.59 ;
      RECT MASK 1 28.779 99.54 28.839 100.59 ;
      RECT MASK 1 29.053 99.54 29.113 100.59 ;
      RECT MASK 1 29.327 99.54 29.387 100.59 ;
      RECT MASK 1 29.601 99.54 29.661 100.59 ;
      RECT MASK 1 29.875 99.54 29.935 100.59 ;
      RECT MASK 1 30.149 99.54 30.209 100.59 ;
      RECT MASK 1 30.423 99.54 30.483 100.59 ;
      RECT MASK 1 30.697 99.54 30.757 100.59 ;
      RECT MASK 1 30.971 99.54 31.031 100.59 ;
      RECT MASK 1 31.245 99.54 31.305 100.59 ;
      RECT MASK 1 31.519 99.54 31.579 100.59 ;
      RECT MASK 1 31.793 99.54 31.853 100.59 ;
      RECT MASK 1 32.067 99.54 32.127 100.59 ;
      RECT MASK 1 32.341 99.54 32.401 100.59 ;
      RECT MASK 1 32.615 99.54 32.675 100.59 ;
      RECT MASK 1 32.889 99.54 32.949 100.59 ;
      RECT MASK 1 33.163 99.54 33.223 100.59 ;
      RECT MASK 1 33.437 99.54 33.497 100.59 ;
      RECT MASK 1 33.711 99.54 33.771 100.59 ;
      RECT MASK 1 33.985 99.54 34.045 100.59 ;
      RECT MASK 1 34.259 99.54 34.319 100.59 ;
      RECT MASK 1 34.533 99.54 34.593 100.59 ;
      RECT MASK 1 34.807 99.54 34.867 100.59 ;
      RECT MASK 1 35.081 99.54 35.141 100.59 ;
      RECT MASK 1 35.355 99.54 35.415 100.59 ;
      RECT MASK 1 35.629 99.54 35.689 100.59 ;
      RECT MASK 1 35.903 99.54 35.963 100.59 ;
      RECT MASK 1 36.177 99.54 36.237 100.59 ;
      RECT MASK 1 36.451 99.54 36.511 100.59 ;
      RECT MASK 1 36.725 99.54 36.785 100.59 ;
      RECT MASK 1 36.999 99.54 37.059 100.59 ;
      RECT MASK 1 37.273 99.54 37.333 100.59 ;
      RECT MASK 1 37.547 99.54 37.607 100.59 ;
      RECT MASK 1 37.821 99.54 37.881 100.59 ;
      RECT MASK 1 38.095 99.54 38.155 100.59 ;
      RECT MASK 1 38.369 99.54 38.429 100.59 ;
      RECT MASK 1 38.643 99.54 38.703 100.59 ;
      RECT MASK 1 38.917 99.54 38.977 100.59 ;
      RECT MASK 1 39.191 99.54 39.251 100.59 ;
      RECT MASK 1 39.465 99.54 39.525 100.59 ;
      RECT MASK 1 39.739 99.54 39.799 100.59 ;
      RECT MASK 1 40.013 99.54 40.073 100.59 ;
      RECT MASK 1 40.287 99.54 40.347 100.59 ;
      RECT MASK 1 40.561 99.54 40.621 100.59 ;
      RECT MASK 1 40.835 99.54 40.895 100.59 ;
      RECT MASK 1 41.109 99.54 41.169 100.59 ;
      RECT MASK 1 41.383 99.54 41.443 100.59 ;
      RECT MASK 1 41.657 99.54 41.717 100.59 ;
      RECT MASK 1 41.931 99.54 41.991 100.59 ;
      RECT MASK 1 42.205 99.54 42.265 100.59 ;
      RECT MASK 1 42.479 99.54 42.539 100.59 ;
      RECT MASK 1 42.753 99.54 42.813 100.59 ;
      RECT MASK 1 43.027 99.54 43.087 100.59 ;
      RECT MASK 1 43.301 99.54 43.361 100.59 ;
      RECT MASK 1 43.575 99.54 43.635 100.59 ;
      RECT MASK 1 45.593 99.54 45.653 100.59 ;
      RECT MASK 1 45.867 99.54 45.927 100.59 ;
      RECT MASK 1 46.141 99.54 46.201 100.59 ;
      RECT MASK 1 46.415 99.54 46.475 100.59 ;
      RECT MASK 1 46.689 99.54 46.749 100.59 ;
      RECT MASK 1 46.963 99.54 47.023 100.59 ;
      RECT MASK 1 47.237 99.54 47.297 100.59 ;
      RECT MASK 1 47.511 99.54 47.571 100.59 ;
      RECT MASK 1 47.785 99.54 47.845 100.59 ;
      RECT MASK 1 48.059 99.54 48.119 100.59 ;
      RECT MASK 1 48.333 99.54 48.393 100.59 ;
      RECT MASK 1 48.607 99.54 48.667 100.59 ;
      RECT MASK 1 48.881 99.54 48.941 100.59 ;
      RECT MASK 1 49.155 99.54 49.215 100.59 ;
      RECT MASK 1 49.429 99.54 49.489 100.59 ;
      RECT MASK 1 49.703 99.54 49.763 100.59 ;
      RECT MASK 1 49.977 99.54 50.037 100.59 ;
      RECT MASK 1 50.251 99.54 50.311 100.59 ;
      RECT MASK 1 50.525 99.54 50.585 100.59 ;
      RECT MASK 1 50.799 99.54 50.859 100.59 ;
      RECT MASK 1 51.073 99.54 51.133 100.59 ;
      RECT MASK 1 51.347 99.54 51.407 100.59 ;
      RECT MASK 1 51.621 99.54 51.681 100.59 ;
      RECT MASK 1 51.895 99.54 51.955 100.59 ;
      RECT MASK 1 52.169 99.54 52.229 100.59 ;
      RECT MASK 1 52.443 99.54 52.503 100.59 ;
      RECT MASK 1 52.717 99.54 52.777 100.59 ;
      RECT MASK 1 52.991 99.54 53.051 100.59 ;
      RECT MASK 1 53.265 99.54 53.325 100.59 ;
      RECT MASK 1 53.539 99.54 53.599 100.59 ;
      RECT MASK 1 53.813 99.54 53.873 100.59 ;
      RECT MASK 1 54.087 99.54 54.147 100.59 ;
      RECT MASK 1 54.361 99.54 54.421 100.59 ;
      RECT MASK 1 54.635 99.54 54.695 100.59 ;
      RECT MASK 1 54.909 99.54 54.969 100.59 ;
      RECT MASK 1 55.183 99.54 55.243 100.59 ;
      RECT MASK 1 55.457 99.54 55.517 100.59 ;
      RECT MASK 1 55.731 99.54 55.791 100.59 ;
      RECT MASK 1 56.005 99.54 56.065 100.59 ;
      RECT MASK 1 56.279 99.54 56.339 100.59 ;
      RECT MASK 1 56.553 99.54 56.613 100.59 ;
      RECT MASK 1 56.827 99.54 56.887 100.59 ;
      RECT MASK 1 57.101 99.54 57.161 100.59 ;
      RECT MASK 1 57.375 99.54 57.435 100.59 ;
      RECT MASK 1 57.649 99.54 57.709 100.59 ;
      RECT MASK 1 57.923 99.54 57.983 100.59 ;
      RECT MASK 1 58.197 99.54 58.257 100.59 ;
      RECT MASK 1 58.471 99.54 58.531 100.59 ;
      RECT MASK 1 58.745 99.54 58.805 100.59 ;
      RECT MASK 1 59.019 99.54 59.079 100.59 ;
      RECT MASK 1 59.293 99.54 59.353 100.59 ;
      RECT MASK 1 59.567 99.54 59.627 100.59 ;
      RECT MASK 1 59.841 99.54 59.901 100.59 ;
      RECT MASK 1 60.115 99.54 60.175 100.59 ;
      RECT MASK 1 60.389 99.54 60.449 100.59 ;
      RECT MASK 1 60.663 99.54 60.723 100.59 ;
      RECT MASK 1 60.937 99.54 60.997 100.59 ;
      RECT MASK 1 61.211 99.54 61.271 100.59 ;
      RECT MASK 1 61.485 99.54 61.545 100.59 ;
      RECT MASK 1 61.759 99.54 61.819 100.59 ;
      RECT MASK 1 62.033 99.54 62.093 100.59 ;
      RECT MASK 1 62.307 99.54 62.367 100.59 ;
      RECT MASK 1 62.581 99.54 62.641 100.59 ;
      RECT MASK 1 62.855 99.54 62.915 100.59 ;
      RECT MASK 1 63.129 99.54 63.189 100.59 ;
      RECT MASK 1 63.403 99.54 63.463 100.59 ;
      RECT MASK 1 63.677 99.54 63.737 100.59 ;
      RECT MASK 1 63.951 99.54 64.011 100.59 ;
      RECT MASK 1 64.225 99.54 64.285 100.59 ;
      RECT MASK 1 64.499 99.54 64.559 100.59 ;
      RECT MASK 1 64.773 99.54 64.833 100.59 ;
      RECT MASK 1 65.047 99.54 65.107 100.59 ;
      RECT MASK 1 65.321 99.54 65.381 100.59 ;
      RECT MASK 1 65.595 99.54 65.655 100.59 ;
      RECT MASK 1 65.869 99.54 65.929 100.59 ;
      RECT MASK 1 66.143 99.54 66.203 100.59 ;
      RECT MASK 1 66.417 99.54 66.477 100.59 ;
      RECT MASK 1 66.691 99.54 66.751 100.59 ;
      RECT MASK 1 66.965 99.54 67.025 100.59 ;
      RECT MASK 1 67.239 99.54 67.299 100.59 ;
      RECT MASK 1 67.513 99.54 67.573 100.59 ;
      RECT MASK 1 67.787 99.54 67.847 100.59 ;
      RECT MASK 1 68.061 99.54 68.121 100.59 ;
      RECT MASK 1 68.335 99.54 68.395 100.59 ;
      RECT MASK 1 68.609 99.54 68.669 100.59 ;
      RECT MASK 1 68.883 99.54 68.943 100.59 ;
      RECT MASK 1 69.157 99.54 69.217 100.59 ;
      RECT MASK 1 69.431 99.54 69.491 100.59 ;
      RECT MASK 1 69.705 99.54 69.765 100.59 ;
      RECT MASK 1 69.979 99.54 70.039 100.59 ;
      RECT MASK 1 70.253 99.54 70.313 100.59 ;
      RECT MASK 1 70.527 99.54 70.587 100.59 ;
      RECT MASK 1 70.801 99.54 70.861 100.59 ;
      RECT MASK 1 71.075 99.54 71.135 100.59 ;
      RECT MASK 1 71.349 99.54 71.409 100.59 ;
      RECT MASK 1 71.623 99.54 71.683 100.59 ;
      RECT MASK 1 71.897 99.54 71.957 100.59 ;
      RECT MASK 1 72.171 99.54 72.231 100.59 ;
      RECT MASK 1 72.445 99.54 72.505 100.59 ;
      RECT MASK 1 72.719 99.54 72.779 100.59 ;
      RECT MASK 1 72.993 99.54 73.053 100.59 ;
      RECT MASK 1 73.267 99.54 73.327 100.59 ;
      RECT MASK 1 73.541 99.54 73.601 100.59 ;
      RECT MASK 1 73.815 99.54 73.875 100.59 ;
      RECT MASK 1 74.089 99.54 74.149 100.59 ;
      RECT MASK 1 74.363 99.54 74.423 100.59 ;
      RECT MASK 1 74.637 99.54 74.697 100.59 ;
      RECT MASK 1 74.911 99.54 74.971 100.59 ;
      RECT MASK 1 75.185 99.54 75.245 100.59 ;
      RECT MASK 1 75.459 99.54 75.519 100.59 ;
      RECT MASK 1 75.733 99.54 75.793 100.59 ;
      RECT MASK 1 76.007 99.54 76.067 100.59 ;
      RECT MASK 1 76.281 99.54 76.341 100.59 ;
      RECT MASK 1 76.555 99.54 76.615 100.59 ;
      RECT MASK 1 76.829 99.54 76.889 100.59 ;
      RECT MASK 1 77.103 99.54 77.163 100.59 ;
      RECT MASK 1 77.377 99.54 77.437 100.59 ;
      RECT MASK 1 77.651 99.54 77.711 100.59 ;
      RECT MASK 1 77.925 99.54 77.985 100.59 ;
      RECT MASK 1 78.199 99.54 78.259 100.59 ;
      RECT MASK 1 78.473 99.54 78.533 100.59 ;
      RECT MASK 1 78.747 99.54 78.807 100.59 ;
      RECT MASK 1 79.021 99.54 79.081 100.59 ;
      RECT MASK 1 79.295 99.54 79.355 100.59 ;
      RECT MASK 1 79.569 99.54 79.629 100.59 ;
      RECT MASK 1 79.843 99.54 79.903 100.59 ;
      RECT MASK 1 80.117 99.54 80.177 100.59 ;
      RECT MASK 1 80.391 99.54 80.451 100.59 ;
      RECT MASK 1 80.665 99.54 80.725 100.59 ;
      RECT MASK 1 80.939 99.54 80.999 100.59 ;
      RECT MASK 1 81.213 99.54 81.273 100.59 ;
      RECT MASK 1 81.487 99.54 81.547 100.59 ;
      RECT MASK 1 81.761 99.54 81.821 100.59 ;
      RECT MASK 1 82.035 99.54 82.095 100.59 ;
      RECT MASK 1 82.309 99.54 82.369 100.59 ;
      RECT MASK 1 82.583 99.54 82.643 100.59 ;
      RECT MASK 1 82.857 99.54 82.917 100.59 ;
      RECT MASK 1 83.131 99.54 83.191 100.59 ;
      RECT MASK 1 83.405 99.54 83.465 100.59 ;
      RECT MASK 1 83.679 99.54 83.739 100.59 ;
      RECT MASK 1 83.953 99.54 84.013 100.59 ;
      RECT MASK 1 84.227 99.54 84.287 100.59 ;
      RECT MASK 1 84.501 99.54 84.561 100.59 ;
      RECT MASK 1 84.775 99.54 84.835 100.59 ;
      RECT MASK 1 85.049 99.54 85.109 100.59 ;
      RECT MASK 1 85.323 99.54 85.383 100.59 ;
      RECT MASK 1 85.597 99.54 85.657 100.59 ;
      RECT MASK 1 85.871 99.54 85.931 100.59 ;
      RECT MASK 1 86.145 99.54 86.205 100.59 ;
      RECT MASK 1 86.419 99.54 86.479 100.59 ;
      RECT MASK 1 86.693 99.54 86.753 100.59 ;
      RECT MASK 1 86.967 99.54 87.027 100.59 ;
      RECT MASK 1 88.952 99.54 89.012 100.59 ;
      RECT MASK 1 89.226 99.54 89.286 100.59 ;
      RECT MASK 1 89.5 99.54 89.56 100.59 ;
      RECT MASK 1 89.774 99.54 89.834 100.59 ;
      RECT MASK 1 90.048 99.54 90.108 100.59 ;
      RECT MASK 1 90.322 99.54 90.382 100.59 ;
      RECT MASK 1 90.596 99.54 90.656 100.59 ;
      RECT MASK 1 90.87 99.54 90.93 100.59 ;
      RECT MASK 1 91.144 99.54 91.204 100.59 ;
      RECT MASK 1 91.418 99.54 91.478 100.59 ;
      RECT MASK 1 91.692 99.54 91.752 100.59 ;
      RECT MASK 1 91.966 99.54 92.026 100.59 ;
      RECT MASK 1 92.24 99.54 92.3 100.59 ;
      RECT MASK 1 92.514 99.54 92.574 100.59 ;
      RECT MASK 1 92.788 99.54 92.848 100.59 ;
      RECT MASK 1 93.062 99.54 93.122 100.59 ;
      RECT MASK 1 93.336 99.54 93.396 100.59 ;
      RECT MASK 1 93.61 99.54 93.67 100.59 ;
      RECT MASK 1 93.884 99.54 93.944 100.59 ;
      RECT MASK 1 94.158 99.54 94.218 100.59 ;
      RECT MASK 1 94.432 99.54 94.492 100.59 ;
      RECT MASK 1 94.706 99.54 94.766 100.59 ;
      RECT MASK 1 94.98 99.54 95.04 100.59 ;
      RECT MASK 1 95.254 99.54 95.314 100.59 ;
      RECT MASK 1 95.528 99.54 95.588 100.59 ;
      RECT MASK 1 95.802 99.54 95.862 100.59 ;
      RECT MASK 1 96.076 99.54 96.136 100.59 ;
      RECT MASK 1 96.35 99.54 96.41 100.59 ;
      RECT MASK 1 96.624 99.54 96.684 100.59 ;
      RECT MASK 1 96.898 99.54 96.958 100.59 ;
      RECT MASK 1 97.172 99.54 97.232 100.59 ;
      RECT MASK 1 97.446 99.54 97.506 100.59 ;
      RECT MASK 1 97.72 99.54 97.78 100.59 ;
      RECT MASK 1 97.994 99.54 98.054 100.59 ;
      RECT MASK 1 98.268 99.54 98.328 100.59 ;
      RECT MASK 1 98.542 99.54 98.602 100.59 ;
      RECT MASK 1 98.816 99.54 98.876 100.59 ;
      RECT MASK 1 99.09 99.54 99.15 100.59 ;
      RECT MASK 1 99.364 99.54 99.424 100.59 ;
      RECT MASK 1 99.638 99.54 99.698 100.59 ;
      RECT MASK 1 99.912 99.54 99.972 100.59 ;
      RECT MASK 1 100.186 99.54 100.246 100.59 ;
      RECT MASK 1 100.46 99.54 100.52 100.59 ;
      RECT MASK 1 100.734 99.54 100.794 100.59 ;
      RECT MASK 1 101.008 99.54 101.068 100.59 ;
      RECT MASK 1 101.282 99.54 101.342 100.59 ;
      RECT MASK 1 101.556 99.54 101.616 100.59 ;
      RECT MASK 1 101.83 99.54 101.89 100.59 ;
      RECT MASK 1 102.104 99.54 102.164 100.59 ;
      RECT MASK 1 102.378 99.54 102.438 100.59 ;
      RECT MASK 1 102.652 99.54 102.712 100.59 ;
      RECT MASK 1 102.926 99.54 102.986 100.59 ;
      RECT MASK 1 103.2 99.54 103.26 100.59 ;
      RECT MASK 1 103.474 99.54 103.534 100.59 ;
      RECT MASK 1 103.748 99.54 103.808 100.59 ;
      RECT MASK 1 104.022 99.54 104.082 100.59 ;
      RECT MASK 1 104.296 99.54 104.356 100.59 ;
      RECT MASK 1 104.57 99.54 104.63 100.59 ;
      RECT MASK 1 104.844 99.54 104.904 100.59 ;
      RECT MASK 1 105.118 99.54 105.178 100.59 ;
      RECT MASK 1 105.392 99.54 105.452 100.59 ;
      RECT MASK 1 105.666 99.54 105.726 100.59 ;
      RECT MASK 1 105.94 99.54 106 100.59 ;
      RECT MASK 1 106.214 99.54 106.274 100.59 ;
      RECT MASK 1 106.488 99.54 106.548 100.59 ;
      RECT MASK 1 106.762 99.54 106.822 100.59 ;
      RECT MASK 1 107.036 99.54 107.096 100.59 ;
      RECT MASK 1 107.31 99.54 107.37 100.59 ;
      RECT MASK 1 107.584 99.54 107.644 100.59 ;
      RECT MASK 1 107.858 99.54 107.918 100.59 ;
      RECT MASK 1 108.132 99.54 108.192 100.59 ;
      RECT MASK 1 108.406 99.54 108.466 100.59 ;
      RECT MASK 1 108.68 99.54 108.74 100.59 ;
      RECT MASK 1 108.954 99.54 109.014 100.59 ;
      RECT MASK 1 109.228 99.54 109.288 100.59 ;
      RECT MASK 1 109.502 99.54 109.562 100.59 ;
      RECT MASK 1 109.776 99.54 109.836 100.59 ;
      RECT MASK 1 110.05 99.54 110.11 100.59 ;
      RECT MASK 1 110.324 99.54 110.384 100.59 ;
      RECT MASK 1 110.598 99.54 110.658 100.59 ;
      RECT MASK 1 110.872 99.54 110.932 100.59 ;
      RECT MASK 1 111.146 99.54 111.206 100.59 ;
      RECT MASK 1 111.42 99.54 111.48 100.59 ;
      RECT MASK 1 111.694 99.54 111.754 100.59 ;
      RECT MASK 1 111.968 99.54 112.028 100.59 ;
      RECT MASK 1 112.242 99.54 112.302 100.59 ;
      RECT MASK 1 112.516 99.54 112.576 100.59 ;
      RECT MASK 1 112.79 99.54 112.85 100.59 ;
      RECT MASK 1 113.064 99.54 113.124 100.59 ;
      RECT MASK 1 113.338 99.54 113.398 100.59 ;
      RECT MASK 1 113.612 99.54 113.672 100.59 ;
      RECT MASK 1 113.886 99.54 113.946 100.59 ;
      RECT MASK 1 114.16 99.54 114.22 100.59 ;
      RECT MASK 1 114.434 99.54 114.494 100.59 ;
      RECT MASK 1 114.708 99.54 114.768 100.59 ;
      RECT MASK 1 114.982 99.54 115.042 100.59 ;
      RECT MASK 1 115.256 99.54 115.316 100.59 ;
      RECT MASK 1 115.53 99.54 115.59 100.59 ;
      RECT MASK 1 115.804 99.54 115.864 100.59 ;
      RECT MASK 1 116.078 99.54 116.138 100.59 ;
      RECT MASK 1 116.352 99.54 116.412 100.59 ;
      RECT MASK 1 116.626 99.54 116.686 100.59 ;
      RECT MASK 1 116.9 99.54 116.96 100.59 ;
      RECT MASK 1 117.174 99.54 117.234 100.59 ;
      RECT MASK 1 117.448 99.54 117.508 100.59 ;
      RECT MASK 1 117.722 99.54 117.782 100.59 ;
      RECT MASK 1 117.996 99.54 118.056 100.59 ;
      RECT MASK 1 118.27 99.54 118.33 100.59 ;
      RECT MASK 1 118.544 99.54 118.604 100.59 ;
      RECT MASK 1 118.818 99.54 118.878 100.59 ;
      RECT MASK 1 119.092 99.54 119.152 100.59 ;
      RECT MASK 1 119.366 99.54 119.426 100.59 ;
      RECT MASK 1 119.64 99.54 119.7 100.59 ;
      RECT MASK 1 119.914 99.54 119.974 100.59 ;
      RECT MASK 1 120.188 99.54 120.248 100.59 ;
      RECT MASK 1 120.462 99.54 120.522 100.59 ;
      RECT MASK 1 120.736 99.54 120.796 100.59 ;
      RECT MASK 1 121.01 99.54 121.07 100.59 ;
      RECT MASK 1 121.284 99.54 121.344 100.59 ;
      RECT MASK 1 121.558 99.54 121.618 100.59 ;
      RECT MASK 1 121.832 99.54 121.892 100.59 ;
      RECT MASK 1 122.106 99.54 122.166 100.59 ;
      RECT MASK 1 122.38 99.54 122.44 100.59 ;
      RECT MASK 1 122.654 99.54 122.714 100.59 ;
      RECT MASK 1 122.928 99.54 122.988 100.59 ;
      RECT MASK 1 123.202 99.54 123.262 100.59 ;
      RECT MASK 1 123.476 99.54 123.536 100.59 ;
      RECT MASK 1 123.75 99.54 123.81 100.59 ;
      RECT MASK 1 124.024 99.54 124.084 100.59 ;
      RECT MASK 1 124.298 99.54 124.358 100.59 ;
      RECT MASK 1 124.572 99.54 124.632 100.59 ;
      RECT MASK 1 124.846 99.54 124.906 100.59 ;
      RECT MASK 1 125.12 99.54 125.18 100.59 ;
      RECT MASK 1 125.394 99.54 125.454 100.59 ;
      RECT MASK 1 125.668 99.54 125.728 100.59 ;
      RECT MASK 1 125.942 99.54 126.002 100.59 ;
      RECT MASK 1 126.216 99.54 126.276 100.59 ;
      RECT MASK 1 126.49 99.54 126.55 100.59 ;
      RECT MASK 1 126.764 99.54 126.824 100.59 ;
      RECT MASK 1 127.038 99.54 127.098 100.59 ;
      RECT MASK 1 127.312 99.54 127.372 100.59 ;
      RECT MASK 1 127.586 99.54 127.646 100.59 ;
      RECT MASK 1 2.201 101.25 2.261 102.3 ;
      RECT MASK 1 2.475 101.25 2.535 102.3 ;
      RECT MASK 1 2.749 101.25 2.809 102.3 ;
      RECT MASK 1 3.023 101.25 3.083 102.3 ;
      RECT MASK 1 3.297 101.25 3.357 102.3 ;
      RECT MASK 1 3.571 101.25 3.631 102.3 ;
      RECT MASK 1 3.845 101.25 3.905 102.3 ;
      RECT MASK 1 4.119 101.25 4.179 102.3 ;
      RECT MASK 1 4.393 101.25 4.453 102.3 ;
      RECT MASK 1 4.667 101.25 4.727 102.3 ;
      RECT MASK 1 4.941 101.25 5.001 102.3 ;
      RECT MASK 1 5.215 101.25 5.275 102.3 ;
      RECT MASK 1 5.489 101.25 5.549 102.3 ;
      RECT MASK 1 5.763 101.25 5.823 102.3 ;
      RECT MASK 1 6.037 101.25 6.097 102.3 ;
      RECT MASK 1 6.311 101.25 6.371 102.3 ;
      RECT MASK 1 6.585 101.25 6.645 102.3 ;
      RECT MASK 1 6.859 101.25 6.919 102.3 ;
      RECT MASK 1 7.133 101.25 7.193 102.3 ;
      RECT MASK 1 7.407 101.25 7.467 102.3 ;
      RECT MASK 1 7.681 101.25 7.741 102.3 ;
      RECT MASK 1 7.955 101.25 8.015 102.3 ;
      RECT MASK 1 8.229 101.25 8.289 102.3 ;
      RECT MASK 1 8.503 101.25 8.563 102.3 ;
      RECT MASK 1 8.777 101.25 8.837 102.3 ;
      RECT MASK 1 9.051 101.25 9.111 102.3 ;
      RECT MASK 1 9.325 101.25 9.385 102.3 ;
      RECT MASK 1 9.599 101.25 9.659 102.3 ;
      RECT MASK 1 9.873 101.25 9.933 102.3 ;
      RECT MASK 1 10.147 101.25 10.207 102.3 ;
      RECT MASK 1 10.421 101.25 10.481 102.3 ;
      RECT MASK 1 10.695 101.25 10.755 102.3 ;
      RECT MASK 1 10.969 101.25 11.029 102.3 ;
      RECT MASK 1 11.243 101.25 11.303 102.3 ;
      RECT MASK 1 11.517 101.25 11.577 102.3 ;
      RECT MASK 1 11.791 101.25 11.851 102.3 ;
      RECT MASK 1 12.065 101.25 12.125 102.3 ;
      RECT MASK 1 12.339 101.25 12.399 102.3 ;
      RECT MASK 1 12.613 101.25 12.673 102.3 ;
      RECT MASK 1 12.887 101.25 12.947 102.3 ;
      RECT MASK 1 13.161 101.25 13.221 102.3 ;
      RECT MASK 1 13.435 101.25 13.495 102.3 ;
      RECT MASK 1 13.709 101.25 13.769 102.3 ;
      RECT MASK 1 13.983 101.25 14.043 102.3 ;
      RECT MASK 1 14.257 101.25 14.317 102.3 ;
      RECT MASK 1 14.531 101.25 14.591 102.3 ;
      RECT MASK 1 14.805 101.25 14.865 102.3 ;
      RECT MASK 1 15.079 101.25 15.139 102.3 ;
      RECT MASK 1 15.353 101.25 15.413 102.3 ;
      RECT MASK 1 15.627 101.25 15.687 102.3 ;
      RECT MASK 1 15.901 101.25 15.961 102.3 ;
      RECT MASK 1 16.175 101.25 16.235 102.3 ;
      RECT MASK 1 16.449 101.25 16.509 102.3 ;
      RECT MASK 1 16.723 101.25 16.783 102.3 ;
      RECT MASK 1 16.997 101.25 17.057 102.3 ;
      RECT MASK 1 17.271 101.25 17.331 102.3 ;
      RECT MASK 1 17.545 101.25 17.605 102.3 ;
      RECT MASK 1 17.819 101.25 17.879 102.3 ;
      RECT MASK 1 18.093 101.25 18.153 102.3 ;
      RECT MASK 1 18.367 101.25 18.427 102.3 ;
      RECT MASK 1 18.641 101.25 18.701 102.3 ;
      RECT MASK 1 18.915 101.25 18.975 102.3 ;
      RECT MASK 1 19.189 101.25 19.249 102.3 ;
      RECT MASK 1 19.463 101.25 19.523 102.3 ;
      RECT MASK 1 19.737 101.25 19.797 102.3 ;
      RECT MASK 1 20.011 101.25 20.071 102.3 ;
      RECT MASK 1 20.285 101.25 20.345 102.3 ;
      RECT MASK 1 20.559 101.25 20.619 102.3 ;
      RECT MASK 1 20.833 101.25 20.893 102.3 ;
      RECT MASK 1 21.107 101.25 21.167 102.3 ;
      RECT MASK 1 21.381 101.25 21.441 102.3 ;
      RECT MASK 1 21.655 101.25 21.715 102.3 ;
      RECT MASK 1 21.929 101.25 21.989 102.3 ;
      RECT MASK 1 22.203 101.25 22.263 102.3 ;
      RECT MASK 1 22.477 101.25 22.537 102.3 ;
      RECT MASK 1 22.751 101.25 22.811 102.3 ;
      RECT MASK 1 23.025 101.25 23.085 102.3 ;
      RECT MASK 1 23.299 101.25 23.359 102.3 ;
      RECT MASK 1 23.573 101.25 23.633 102.3 ;
      RECT MASK 1 23.847 101.25 23.907 102.3 ;
      RECT MASK 1 24.121 101.25 24.181 102.3 ;
      RECT MASK 1 24.395 101.25 24.455 102.3 ;
      RECT MASK 1 24.669 101.25 24.729 102.3 ;
      RECT MASK 1 24.943 101.25 25.003 102.3 ;
      RECT MASK 1 25.217 101.25 25.277 102.3 ;
      RECT MASK 1 25.491 101.25 25.551 102.3 ;
      RECT MASK 1 25.765 101.25 25.825 102.3 ;
      RECT MASK 1 26.039 101.25 26.099 102.3 ;
      RECT MASK 1 26.313 101.25 26.373 102.3 ;
      RECT MASK 1 26.587 101.25 26.647 102.3 ;
      RECT MASK 1 26.861 101.25 26.921 102.3 ;
      RECT MASK 1 27.135 101.25 27.195 102.3 ;
      RECT MASK 1 27.409 101.25 27.469 102.3 ;
      RECT MASK 1 27.683 101.25 27.743 102.3 ;
      RECT MASK 1 27.957 101.25 28.017 102.3 ;
      RECT MASK 1 28.231 101.25 28.291 102.3 ;
      RECT MASK 1 28.505 101.25 28.565 102.3 ;
      RECT MASK 1 28.779 101.25 28.839 102.3 ;
      RECT MASK 1 29.053 101.25 29.113 102.3 ;
      RECT MASK 1 29.327 101.25 29.387 102.3 ;
      RECT MASK 1 29.601 101.25 29.661 102.3 ;
      RECT MASK 1 29.875 101.25 29.935 102.3 ;
      RECT MASK 1 30.149 101.25 30.209 102.3 ;
      RECT MASK 1 30.423 101.25 30.483 102.3 ;
      RECT MASK 1 30.697 101.25 30.757 102.3 ;
      RECT MASK 1 30.971 101.25 31.031 102.3 ;
      RECT MASK 1 31.245 101.25 31.305 102.3 ;
      RECT MASK 1 31.519 101.25 31.579 102.3 ;
      RECT MASK 1 31.793 101.25 31.853 102.3 ;
      RECT MASK 1 32.067 101.25 32.127 102.3 ;
      RECT MASK 1 32.341 101.25 32.401 102.3 ;
      RECT MASK 1 32.615 101.25 32.675 102.3 ;
      RECT MASK 1 32.889 101.25 32.949 102.3 ;
      RECT MASK 1 33.163 101.25 33.223 102.3 ;
      RECT MASK 1 33.437 101.25 33.497 102.3 ;
      RECT MASK 1 33.711 101.25 33.771 102.3 ;
      RECT MASK 1 33.985 101.25 34.045 102.3 ;
      RECT MASK 1 34.259 101.25 34.319 102.3 ;
      RECT MASK 1 34.533 101.25 34.593 102.3 ;
      RECT MASK 1 34.807 101.25 34.867 102.3 ;
      RECT MASK 1 35.081 101.25 35.141 102.3 ;
      RECT MASK 1 35.355 101.25 35.415 102.3 ;
      RECT MASK 1 35.629 101.25 35.689 102.3 ;
      RECT MASK 1 35.903 101.25 35.963 102.3 ;
      RECT MASK 1 36.177 101.25 36.237 102.3 ;
      RECT MASK 1 36.451 101.25 36.511 102.3 ;
      RECT MASK 1 36.725 101.25 36.785 102.3 ;
      RECT MASK 1 36.999 101.25 37.059 102.3 ;
      RECT MASK 1 37.273 101.25 37.333 102.3 ;
      RECT MASK 1 37.547 101.25 37.607 102.3 ;
      RECT MASK 1 37.821 101.25 37.881 102.3 ;
      RECT MASK 1 38.095 101.25 38.155 102.3 ;
      RECT MASK 1 38.369 101.25 38.429 102.3 ;
      RECT MASK 1 38.643 101.25 38.703 102.3 ;
      RECT MASK 1 38.917 101.25 38.977 102.3 ;
      RECT MASK 1 39.191 101.25 39.251 102.3 ;
      RECT MASK 1 39.465 101.25 39.525 102.3 ;
      RECT MASK 1 39.739 101.25 39.799 102.3 ;
      RECT MASK 1 40.013 101.25 40.073 102.3 ;
      RECT MASK 1 40.287 101.25 40.347 102.3 ;
      RECT MASK 1 40.561 101.25 40.621 102.3 ;
      RECT MASK 1 40.835 101.25 40.895 102.3 ;
      RECT MASK 1 41.109 101.25 41.169 102.3 ;
      RECT MASK 1 41.383 101.25 41.443 102.3 ;
      RECT MASK 1 41.657 101.25 41.717 102.3 ;
      RECT MASK 1 41.931 101.25 41.991 102.3 ;
      RECT MASK 1 42.205 101.25 42.265 102.3 ;
      RECT MASK 1 42.479 101.25 42.539 102.3 ;
      RECT MASK 1 42.753 101.25 42.813 102.3 ;
      RECT MASK 1 43.027 101.25 43.087 102.3 ;
      RECT MASK 1 43.301 101.25 43.361 102.3 ;
      RECT MASK 1 43.575 101.25 43.635 102.3 ;
      RECT MASK 1 45.593 101.25 45.653 102.3 ;
      RECT MASK 1 45.867 101.25 45.927 102.3 ;
      RECT MASK 1 46.141 101.25 46.201 102.3 ;
      RECT MASK 1 46.415 101.25 46.475 102.3 ;
      RECT MASK 1 46.689 101.25 46.749 102.3 ;
      RECT MASK 1 46.963 101.25 47.023 102.3 ;
      RECT MASK 1 47.237 101.25 47.297 102.3 ;
      RECT MASK 1 47.511 101.25 47.571 102.3 ;
      RECT MASK 1 47.785 101.25 47.845 102.3 ;
      RECT MASK 1 48.059 101.25 48.119 102.3 ;
      RECT MASK 1 48.333 101.25 48.393 102.3 ;
      RECT MASK 1 48.607 101.25 48.667 102.3 ;
      RECT MASK 1 48.881 101.25 48.941 102.3 ;
      RECT MASK 1 49.155 101.25 49.215 102.3 ;
      RECT MASK 1 49.429 101.25 49.489 102.3 ;
      RECT MASK 1 49.703 101.25 49.763 102.3 ;
      RECT MASK 1 49.977 101.25 50.037 102.3 ;
      RECT MASK 1 50.251 101.25 50.311 102.3 ;
      RECT MASK 1 50.525 101.25 50.585 102.3 ;
      RECT MASK 1 50.799 101.25 50.859 102.3 ;
      RECT MASK 1 51.073 101.25 51.133 102.3 ;
      RECT MASK 1 51.347 101.25 51.407 102.3 ;
      RECT MASK 1 51.621 101.25 51.681 102.3 ;
      RECT MASK 1 51.895 101.25 51.955 102.3 ;
      RECT MASK 1 52.169 101.25 52.229 102.3 ;
      RECT MASK 1 52.443 101.25 52.503 102.3 ;
      RECT MASK 1 52.717 101.25 52.777 102.3 ;
      RECT MASK 1 52.991 101.25 53.051 102.3 ;
      RECT MASK 1 53.265 101.25 53.325 102.3 ;
      RECT MASK 1 53.539 101.25 53.599 102.3 ;
      RECT MASK 1 53.813 101.25 53.873 102.3 ;
      RECT MASK 1 54.087 101.25 54.147 102.3 ;
      RECT MASK 1 54.361 101.25 54.421 102.3 ;
      RECT MASK 1 54.635 101.25 54.695 102.3 ;
      RECT MASK 1 54.909 101.25 54.969 102.3 ;
      RECT MASK 1 55.183 101.25 55.243 102.3 ;
      RECT MASK 1 55.457 101.25 55.517 102.3 ;
      RECT MASK 1 55.731 101.25 55.791 102.3 ;
      RECT MASK 1 56.005 101.25 56.065 102.3 ;
      RECT MASK 1 56.279 101.25 56.339 102.3 ;
      RECT MASK 1 56.553 101.25 56.613 102.3 ;
      RECT MASK 1 56.827 101.25 56.887 102.3 ;
      RECT MASK 1 57.101 101.25 57.161 102.3 ;
      RECT MASK 1 57.375 101.25 57.435 102.3 ;
      RECT MASK 1 57.649 101.25 57.709 102.3 ;
      RECT MASK 1 57.923 101.25 57.983 102.3 ;
      RECT MASK 1 58.197 101.25 58.257 102.3 ;
      RECT MASK 1 58.471 101.25 58.531 102.3 ;
      RECT MASK 1 58.745 101.25 58.805 102.3 ;
      RECT MASK 1 59.019 101.25 59.079 102.3 ;
      RECT MASK 1 59.293 101.25 59.353 102.3 ;
      RECT MASK 1 59.567 101.25 59.627 102.3 ;
      RECT MASK 1 59.841 101.25 59.901 102.3 ;
      RECT MASK 1 60.115 101.25 60.175 102.3 ;
      RECT MASK 1 60.389 101.25 60.449 102.3 ;
      RECT MASK 1 60.663 101.25 60.723 102.3 ;
      RECT MASK 1 60.937 101.25 60.997 102.3 ;
      RECT MASK 1 61.211 101.25 61.271 102.3 ;
      RECT MASK 1 61.485 101.25 61.545 102.3 ;
      RECT MASK 1 61.759 101.25 61.819 102.3 ;
      RECT MASK 1 62.033 101.25 62.093 102.3 ;
      RECT MASK 1 62.307 101.25 62.367 102.3 ;
      RECT MASK 1 62.581 101.25 62.641 102.3 ;
      RECT MASK 1 62.855 101.25 62.915 102.3 ;
      RECT MASK 1 63.129 101.25 63.189 102.3 ;
      RECT MASK 1 63.403 101.25 63.463 102.3 ;
      RECT MASK 1 63.677 101.25 63.737 102.3 ;
      RECT MASK 1 63.951 101.25 64.011 102.3 ;
      RECT MASK 1 64.225 101.25 64.285 102.3 ;
      RECT MASK 1 64.499 101.25 64.559 102.3 ;
      RECT MASK 1 64.773 101.25 64.833 102.3 ;
      RECT MASK 1 65.047 101.25 65.107 102.3 ;
      RECT MASK 1 65.321 101.25 65.381 102.3 ;
      RECT MASK 1 65.595 101.25 65.655 102.3 ;
      RECT MASK 1 65.869 101.25 65.929 102.3 ;
      RECT MASK 1 66.143 101.25 66.203 102.3 ;
      RECT MASK 1 66.417 101.25 66.477 102.3 ;
      RECT MASK 1 66.691 101.25 66.751 102.3 ;
      RECT MASK 1 66.965 101.25 67.025 102.3 ;
      RECT MASK 1 67.239 101.25 67.299 102.3 ;
      RECT MASK 1 67.513 101.25 67.573 102.3 ;
      RECT MASK 1 67.787 101.25 67.847 102.3 ;
      RECT MASK 1 68.061 101.25 68.121 102.3 ;
      RECT MASK 1 68.335 101.25 68.395 102.3 ;
      RECT MASK 1 68.609 101.25 68.669 102.3 ;
      RECT MASK 1 68.883 101.25 68.943 102.3 ;
      RECT MASK 1 69.157 101.25 69.217 102.3 ;
      RECT MASK 1 69.431 101.25 69.491 102.3 ;
      RECT MASK 1 69.705 101.25 69.765 102.3 ;
      RECT MASK 1 69.979 101.25 70.039 102.3 ;
      RECT MASK 1 70.253 101.25 70.313 102.3 ;
      RECT MASK 1 70.527 101.25 70.587 102.3 ;
      RECT MASK 1 70.801 101.25 70.861 102.3 ;
      RECT MASK 1 71.075 101.25 71.135 102.3 ;
      RECT MASK 1 71.349 101.25 71.409 102.3 ;
      RECT MASK 1 71.623 101.25 71.683 102.3 ;
      RECT MASK 1 71.897 101.25 71.957 102.3 ;
      RECT MASK 1 72.171 101.25 72.231 102.3 ;
      RECT MASK 1 72.445 101.25 72.505 102.3 ;
      RECT MASK 1 72.719 101.25 72.779 102.3 ;
      RECT MASK 1 72.993 101.25 73.053 102.3 ;
      RECT MASK 1 73.267 101.25 73.327 102.3 ;
      RECT MASK 1 73.541 101.25 73.601 102.3 ;
      RECT MASK 1 73.815 101.25 73.875 102.3 ;
      RECT MASK 1 74.089 101.25 74.149 102.3 ;
      RECT MASK 1 74.363 101.25 74.423 102.3 ;
      RECT MASK 1 74.637 101.25 74.697 102.3 ;
      RECT MASK 1 74.911 101.25 74.971 102.3 ;
      RECT MASK 1 75.185 101.25 75.245 102.3 ;
      RECT MASK 1 75.459 101.25 75.519 102.3 ;
      RECT MASK 1 75.733 101.25 75.793 102.3 ;
      RECT MASK 1 76.007 101.25 76.067 102.3 ;
      RECT MASK 1 76.281 101.25 76.341 102.3 ;
      RECT MASK 1 76.555 101.25 76.615 102.3 ;
      RECT MASK 1 76.829 101.25 76.889 102.3 ;
      RECT MASK 1 77.103 101.25 77.163 102.3 ;
      RECT MASK 1 77.377 101.25 77.437 102.3 ;
      RECT MASK 1 77.651 101.25 77.711 102.3 ;
      RECT MASK 1 77.925 101.25 77.985 102.3 ;
      RECT MASK 1 78.199 101.25 78.259 102.3 ;
      RECT MASK 1 78.473 101.25 78.533 102.3 ;
      RECT MASK 1 78.747 101.25 78.807 102.3 ;
      RECT MASK 1 79.021 101.25 79.081 102.3 ;
      RECT MASK 1 79.295 101.25 79.355 102.3 ;
      RECT MASK 1 79.569 101.25 79.629 102.3 ;
      RECT MASK 1 79.843 101.25 79.903 102.3 ;
      RECT MASK 1 80.117 101.25 80.177 102.3 ;
      RECT MASK 1 80.391 101.25 80.451 102.3 ;
      RECT MASK 1 80.665 101.25 80.725 102.3 ;
      RECT MASK 1 80.939 101.25 80.999 102.3 ;
      RECT MASK 1 81.213 101.25 81.273 102.3 ;
      RECT MASK 1 81.487 101.25 81.547 102.3 ;
      RECT MASK 1 81.761 101.25 81.821 102.3 ;
      RECT MASK 1 82.035 101.25 82.095 102.3 ;
      RECT MASK 1 82.309 101.25 82.369 102.3 ;
      RECT MASK 1 82.583 101.25 82.643 102.3 ;
      RECT MASK 1 82.857 101.25 82.917 102.3 ;
      RECT MASK 1 83.131 101.25 83.191 102.3 ;
      RECT MASK 1 83.405 101.25 83.465 102.3 ;
      RECT MASK 1 83.679 101.25 83.739 102.3 ;
      RECT MASK 1 83.953 101.25 84.013 102.3 ;
      RECT MASK 1 84.227 101.25 84.287 102.3 ;
      RECT MASK 1 84.501 101.25 84.561 102.3 ;
      RECT MASK 1 84.775 101.25 84.835 102.3 ;
      RECT MASK 1 85.049 101.25 85.109 102.3 ;
      RECT MASK 1 85.323 101.25 85.383 102.3 ;
      RECT MASK 1 85.597 101.25 85.657 102.3 ;
      RECT MASK 1 85.871 101.25 85.931 102.3 ;
      RECT MASK 1 86.145 101.25 86.205 102.3 ;
      RECT MASK 1 86.419 101.25 86.479 102.3 ;
      RECT MASK 1 86.693 101.25 86.753 102.3 ;
      RECT MASK 1 86.967 101.25 87.027 102.3 ;
      RECT MASK 1 88.952 101.25 89.012 102.3 ;
      RECT MASK 1 89.226 101.25 89.286 102.3 ;
      RECT MASK 1 89.5 101.25 89.56 102.3 ;
      RECT MASK 1 89.774 101.25 89.834 102.3 ;
      RECT MASK 1 90.048 101.25 90.108 102.3 ;
      RECT MASK 1 90.322 101.25 90.382 102.3 ;
      RECT MASK 1 90.596 101.25 90.656 102.3 ;
      RECT MASK 1 90.87 101.25 90.93 102.3 ;
      RECT MASK 1 91.144 101.25 91.204 102.3 ;
      RECT MASK 1 91.418 101.25 91.478 102.3 ;
      RECT MASK 1 91.692 101.25 91.752 102.3 ;
      RECT MASK 1 91.966 101.25 92.026 102.3 ;
      RECT MASK 1 92.24 101.25 92.3 102.3 ;
      RECT MASK 1 92.514 101.25 92.574 102.3 ;
      RECT MASK 1 92.788 101.25 92.848 102.3 ;
      RECT MASK 1 93.062 101.25 93.122 102.3 ;
      RECT MASK 1 93.336 101.25 93.396 102.3 ;
      RECT MASK 1 93.61 101.25 93.67 102.3 ;
      RECT MASK 1 93.884 101.25 93.944 102.3 ;
      RECT MASK 1 94.158 101.25 94.218 102.3 ;
      RECT MASK 1 94.432 101.25 94.492 102.3 ;
      RECT MASK 1 94.706 101.25 94.766 102.3 ;
      RECT MASK 1 94.98 101.25 95.04 102.3 ;
      RECT MASK 1 95.254 101.25 95.314 102.3 ;
      RECT MASK 1 95.528 101.25 95.588 102.3 ;
      RECT MASK 1 95.802 101.25 95.862 102.3 ;
      RECT MASK 1 96.076 101.25 96.136 102.3 ;
      RECT MASK 1 96.35 101.25 96.41 102.3 ;
      RECT MASK 1 96.624 101.25 96.684 102.3 ;
      RECT MASK 1 96.898 101.25 96.958 102.3 ;
      RECT MASK 1 97.172 101.25 97.232 102.3 ;
      RECT MASK 1 97.446 101.25 97.506 102.3 ;
      RECT MASK 1 97.72 101.25 97.78 102.3 ;
      RECT MASK 1 97.994 101.25 98.054 102.3 ;
      RECT MASK 1 98.268 101.25 98.328 102.3 ;
      RECT MASK 1 98.542 101.25 98.602 102.3 ;
      RECT MASK 1 98.816 101.25 98.876 102.3 ;
      RECT MASK 1 99.09 101.25 99.15 102.3 ;
      RECT MASK 1 99.364 101.25 99.424 102.3 ;
      RECT MASK 1 99.638 101.25 99.698 102.3 ;
      RECT MASK 1 99.912 101.25 99.972 102.3 ;
      RECT MASK 1 100.186 101.25 100.246 102.3 ;
      RECT MASK 1 100.46 101.25 100.52 102.3 ;
      RECT MASK 1 100.734 101.25 100.794 102.3 ;
      RECT MASK 1 101.008 101.25 101.068 102.3 ;
      RECT MASK 1 101.282 101.25 101.342 102.3 ;
      RECT MASK 1 101.556 101.25 101.616 102.3 ;
      RECT MASK 1 101.83 101.25 101.89 102.3 ;
      RECT MASK 1 102.104 101.25 102.164 102.3 ;
      RECT MASK 1 102.378 101.25 102.438 102.3 ;
      RECT MASK 1 102.652 101.25 102.712 102.3 ;
      RECT MASK 1 102.926 101.25 102.986 102.3 ;
      RECT MASK 1 103.2 101.25 103.26 102.3 ;
      RECT MASK 1 103.474 101.25 103.534 102.3 ;
      RECT MASK 1 103.748 101.25 103.808 102.3 ;
      RECT MASK 1 104.022 101.25 104.082 102.3 ;
      RECT MASK 1 104.296 101.25 104.356 102.3 ;
      RECT MASK 1 104.57 101.25 104.63 102.3 ;
      RECT MASK 1 104.844 101.25 104.904 102.3 ;
      RECT MASK 1 105.118 101.25 105.178 102.3 ;
      RECT MASK 1 105.392 101.25 105.452 102.3 ;
      RECT MASK 1 105.666 101.25 105.726 102.3 ;
      RECT MASK 1 105.94 101.25 106 102.3 ;
      RECT MASK 1 106.214 101.25 106.274 102.3 ;
      RECT MASK 1 106.488 101.25 106.548 102.3 ;
      RECT MASK 1 106.762 101.25 106.822 102.3 ;
      RECT MASK 1 107.036 101.25 107.096 102.3 ;
      RECT MASK 1 107.31 101.25 107.37 102.3 ;
      RECT MASK 1 107.584 101.25 107.644 102.3 ;
      RECT MASK 1 107.858 101.25 107.918 102.3 ;
      RECT MASK 1 108.132 101.25 108.192 102.3 ;
      RECT MASK 1 108.406 101.25 108.466 102.3 ;
      RECT MASK 1 108.68 101.25 108.74 102.3 ;
      RECT MASK 1 108.954 101.25 109.014 102.3 ;
      RECT MASK 1 109.228 101.25 109.288 102.3 ;
      RECT MASK 1 109.502 101.25 109.562 102.3 ;
      RECT MASK 1 109.776 101.25 109.836 102.3 ;
      RECT MASK 1 110.05 101.25 110.11 102.3 ;
      RECT MASK 1 110.324 101.25 110.384 102.3 ;
      RECT MASK 1 110.598 101.25 110.658 102.3 ;
      RECT MASK 1 110.872 101.25 110.932 102.3 ;
      RECT MASK 1 111.146 101.25 111.206 102.3 ;
      RECT MASK 1 111.42 101.25 111.48 102.3 ;
      RECT MASK 1 111.694 101.25 111.754 102.3 ;
      RECT MASK 1 111.968 101.25 112.028 102.3 ;
      RECT MASK 1 112.242 101.25 112.302 102.3 ;
      RECT MASK 1 112.516 101.25 112.576 102.3 ;
      RECT MASK 1 112.79 101.25 112.85 102.3 ;
      RECT MASK 1 113.064 101.25 113.124 102.3 ;
      RECT MASK 1 113.338 101.25 113.398 102.3 ;
      RECT MASK 1 113.612 101.25 113.672 102.3 ;
      RECT MASK 1 113.886 101.25 113.946 102.3 ;
      RECT MASK 1 114.16 101.25 114.22 102.3 ;
      RECT MASK 1 114.434 101.25 114.494 102.3 ;
      RECT MASK 1 114.708 101.25 114.768 102.3 ;
      RECT MASK 1 114.982 101.25 115.042 102.3 ;
      RECT MASK 1 115.256 101.25 115.316 102.3 ;
      RECT MASK 1 115.53 101.25 115.59 102.3 ;
      RECT MASK 1 115.804 101.25 115.864 102.3 ;
      RECT MASK 1 116.078 101.25 116.138 102.3 ;
      RECT MASK 1 116.352 101.25 116.412 102.3 ;
      RECT MASK 1 116.626 101.25 116.686 102.3 ;
      RECT MASK 1 116.9 101.25 116.96 102.3 ;
      RECT MASK 1 117.174 101.25 117.234 102.3 ;
      RECT MASK 1 117.448 101.25 117.508 102.3 ;
      RECT MASK 1 117.722 101.25 117.782 102.3 ;
      RECT MASK 1 117.996 101.25 118.056 102.3 ;
      RECT MASK 1 118.27 101.25 118.33 102.3 ;
      RECT MASK 1 118.544 101.25 118.604 102.3 ;
      RECT MASK 1 118.818 101.25 118.878 102.3 ;
      RECT MASK 1 119.092 101.25 119.152 102.3 ;
      RECT MASK 1 119.366 101.25 119.426 102.3 ;
      RECT MASK 1 119.64 101.25 119.7 102.3 ;
      RECT MASK 1 119.914 101.25 119.974 102.3 ;
      RECT MASK 1 120.188 101.25 120.248 102.3 ;
      RECT MASK 1 120.462 101.25 120.522 102.3 ;
      RECT MASK 1 120.736 101.25 120.796 102.3 ;
      RECT MASK 1 121.01 101.25 121.07 102.3 ;
      RECT MASK 1 121.284 101.25 121.344 102.3 ;
      RECT MASK 1 121.558 101.25 121.618 102.3 ;
      RECT MASK 1 121.832 101.25 121.892 102.3 ;
      RECT MASK 1 122.106 101.25 122.166 102.3 ;
      RECT MASK 1 122.38 101.25 122.44 102.3 ;
      RECT MASK 1 122.654 101.25 122.714 102.3 ;
      RECT MASK 1 122.928 101.25 122.988 102.3 ;
      RECT MASK 1 123.202 101.25 123.262 102.3 ;
      RECT MASK 1 123.476 101.25 123.536 102.3 ;
      RECT MASK 1 123.75 101.25 123.81 102.3 ;
      RECT MASK 1 124.024 101.25 124.084 102.3 ;
      RECT MASK 1 124.298 101.25 124.358 102.3 ;
      RECT MASK 1 124.572 101.25 124.632 102.3 ;
      RECT MASK 1 124.846 101.25 124.906 102.3 ;
      RECT MASK 1 125.12 101.25 125.18 102.3 ;
      RECT MASK 1 125.394 101.25 125.454 102.3 ;
      RECT MASK 1 125.668 101.25 125.728 102.3 ;
      RECT MASK 1 125.942 101.25 126.002 102.3 ;
      RECT MASK 1 126.216 101.25 126.276 102.3 ;
      RECT MASK 1 126.49 101.25 126.55 102.3 ;
      RECT MASK 1 126.764 101.25 126.824 102.3 ;
      RECT MASK 1 127.038 101.25 127.098 102.3 ;
      RECT MASK 1 127.312 101.25 127.372 102.3 ;
      RECT MASK 1 127.586 101.25 127.646 102.3 ;
      RECT MASK 1 2.201 102.96 2.261 104.01 ;
      RECT MASK 1 2.475 102.96 2.535 104.01 ;
      RECT MASK 1 2.749 102.96 2.809 104.01 ;
      RECT MASK 1 3.023 102.96 3.083 104.01 ;
      RECT MASK 1 3.297 102.96 3.357 104.01 ;
      RECT MASK 1 3.571 102.96 3.631 104.01 ;
      RECT MASK 1 3.845 102.96 3.905 104.01 ;
      RECT MASK 1 4.119 102.96 4.179 104.01 ;
      RECT MASK 1 4.393 102.96 4.453 104.01 ;
      RECT MASK 1 4.667 102.96 4.727 104.01 ;
      RECT MASK 1 4.941 102.96 5.001 104.01 ;
      RECT MASK 1 5.215 102.96 5.275 104.01 ;
      RECT MASK 1 5.489 102.96 5.549 104.01 ;
      RECT MASK 1 5.763 102.96 5.823 104.01 ;
      RECT MASK 1 6.037 102.96 6.097 104.01 ;
      RECT MASK 1 6.311 102.96 6.371 104.01 ;
      RECT MASK 1 6.585 102.96 6.645 104.01 ;
      RECT MASK 1 6.859 102.96 6.919 104.01 ;
      RECT MASK 1 7.133 102.96 7.193 104.01 ;
      RECT MASK 1 7.407 102.96 7.467 104.01 ;
      RECT MASK 1 7.681 102.96 7.741 104.01 ;
      RECT MASK 1 7.955 102.96 8.015 104.01 ;
      RECT MASK 1 8.229 102.96 8.289 104.01 ;
      RECT MASK 1 8.503 102.96 8.563 104.01 ;
      RECT MASK 1 8.777 102.96 8.837 104.01 ;
      RECT MASK 1 9.051 102.96 9.111 104.01 ;
      RECT MASK 1 9.325 102.96 9.385 104.01 ;
      RECT MASK 1 9.599 102.96 9.659 104.01 ;
      RECT MASK 1 9.873 102.96 9.933 104.01 ;
      RECT MASK 1 10.147 102.96 10.207 104.01 ;
      RECT MASK 1 10.421 102.96 10.481 104.01 ;
      RECT MASK 1 10.695 102.96 10.755 104.01 ;
      RECT MASK 1 10.969 102.96 11.029 104.01 ;
      RECT MASK 1 11.243 102.96 11.303 104.01 ;
      RECT MASK 1 11.517 102.96 11.577 104.01 ;
      RECT MASK 1 11.791 102.96 11.851 104.01 ;
      RECT MASK 1 12.065 102.96 12.125 104.01 ;
      RECT MASK 1 12.339 102.96 12.399 104.01 ;
      RECT MASK 1 12.613 102.96 12.673 104.01 ;
      RECT MASK 1 12.887 102.96 12.947 104.01 ;
      RECT MASK 1 13.161 102.96 13.221 104.01 ;
      RECT MASK 1 13.435 102.96 13.495 104.01 ;
      RECT MASK 1 13.709 102.96 13.769 104.01 ;
      RECT MASK 1 13.983 102.96 14.043 104.01 ;
      RECT MASK 1 14.257 102.96 14.317 104.01 ;
      RECT MASK 1 14.531 102.96 14.591 104.01 ;
      RECT MASK 1 14.805 102.96 14.865 104.01 ;
      RECT MASK 1 15.079 102.96 15.139 104.01 ;
      RECT MASK 1 15.353 102.96 15.413 104.01 ;
      RECT MASK 1 15.627 102.96 15.687 104.01 ;
      RECT MASK 1 15.901 102.96 15.961 104.01 ;
      RECT MASK 1 16.175 102.96 16.235 104.01 ;
      RECT MASK 1 16.449 102.96 16.509 104.01 ;
      RECT MASK 1 16.723 102.96 16.783 104.01 ;
      RECT MASK 1 16.997 102.96 17.057 104.01 ;
      RECT MASK 1 17.271 102.96 17.331 104.01 ;
      RECT MASK 1 17.545 102.96 17.605 104.01 ;
      RECT MASK 1 17.819 102.96 17.879 104.01 ;
      RECT MASK 1 18.093 102.96 18.153 104.01 ;
      RECT MASK 1 18.367 102.96 18.427 104.01 ;
      RECT MASK 1 18.641 102.96 18.701 104.01 ;
      RECT MASK 1 18.915 102.96 18.975 104.01 ;
      RECT MASK 1 19.189 102.96 19.249 104.01 ;
      RECT MASK 1 19.463 102.96 19.523 104.01 ;
      RECT MASK 1 19.737 102.96 19.797 104.01 ;
      RECT MASK 1 20.011 102.96 20.071 104.01 ;
      RECT MASK 1 20.285 102.96 20.345 104.01 ;
      RECT MASK 1 20.559 102.96 20.619 104.01 ;
      RECT MASK 1 20.833 102.96 20.893 104.01 ;
      RECT MASK 1 21.107 102.96 21.167 104.01 ;
      RECT MASK 1 21.381 102.96 21.441 104.01 ;
      RECT MASK 1 21.655 102.96 21.715 104.01 ;
      RECT MASK 1 21.929 102.96 21.989 104.01 ;
      RECT MASK 1 22.203 102.96 22.263 104.01 ;
      RECT MASK 1 22.477 102.96 22.537 104.01 ;
      RECT MASK 1 22.751 102.96 22.811 104.01 ;
      RECT MASK 1 23.025 102.96 23.085 104.01 ;
      RECT MASK 1 23.299 102.96 23.359 104.01 ;
      RECT MASK 1 23.573 102.96 23.633 104.01 ;
      RECT MASK 1 23.847 102.96 23.907 104.01 ;
      RECT MASK 1 24.121 102.96 24.181 104.01 ;
      RECT MASK 1 24.395 102.96 24.455 104.01 ;
      RECT MASK 1 24.669 102.96 24.729 104.01 ;
      RECT MASK 1 24.943 102.96 25.003 104.01 ;
      RECT MASK 1 25.217 102.96 25.277 104.01 ;
      RECT MASK 1 25.491 102.96 25.551 104.01 ;
      RECT MASK 1 25.765 102.96 25.825 104.01 ;
      RECT MASK 1 26.039 102.96 26.099 104.01 ;
      RECT MASK 1 26.313 102.96 26.373 104.01 ;
      RECT MASK 1 26.587 102.96 26.647 104.01 ;
      RECT MASK 1 26.861 102.96 26.921 104.01 ;
      RECT MASK 1 27.135 102.96 27.195 104.01 ;
      RECT MASK 1 27.409 102.96 27.469 104.01 ;
      RECT MASK 1 27.683 102.96 27.743 104.01 ;
      RECT MASK 1 27.957 102.96 28.017 104.01 ;
      RECT MASK 1 28.231 102.96 28.291 104.01 ;
      RECT MASK 1 28.505 102.96 28.565 104.01 ;
      RECT MASK 1 28.779 102.96 28.839 104.01 ;
      RECT MASK 1 29.053 102.96 29.113 104.01 ;
      RECT MASK 1 29.327 102.96 29.387 104.01 ;
      RECT MASK 1 29.601 102.96 29.661 104.01 ;
      RECT MASK 1 29.875 102.96 29.935 104.01 ;
      RECT MASK 1 30.149 102.96 30.209 104.01 ;
      RECT MASK 1 30.423 102.96 30.483 104.01 ;
      RECT MASK 1 30.697 102.96 30.757 104.01 ;
      RECT MASK 1 30.971 102.96 31.031 104.01 ;
      RECT MASK 1 31.245 102.96 31.305 104.01 ;
      RECT MASK 1 31.519 102.96 31.579 104.01 ;
      RECT MASK 1 31.793 102.96 31.853 104.01 ;
      RECT MASK 1 32.067 102.96 32.127 104.01 ;
      RECT MASK 1 32.341 102.96 32.401 104.01 ;
      RECT MASK 1 32.615 102.96 32.675 104.01 ;
      RECT MASK 1 32.889 102.96 32.949 104.01 ;
      RECT MASK 1 33.163 102.96 33.223 104.01 ;
      RECT MASK 1 33.437 102.96 33.497 104.01 ;
      RECT MASK 1 33.711 102.96 33.771 104.01 ;
      RECT MASK 1 33.985 102.96 34.045 104.01 ;
      RECT MASK 1 34.259 102.96 34.319 104.01 ;
      RECT MASK 1 34.533 102.96 34.593 104.01 ;
      RECT MASK 1 34.807 102.96 34.867 104.01 ;
      RECT MASK 1 35.081 102.96 35.141 104.01 ;
      RECT MASK 1 35.355 102.96 35.415 104.01 ;
      RECT MASK 1 35.629 102.96 35.689 104.01 ;
      RECT MASK 1 35.903 102.96 35.963 104.01 ;
      RECT MASK 1 36.177 102.96 36.237 104.01 ;
      RECT MASK 1 36.451 102.96 36.511 104.01 ;
      RECT MASK 1 36.725 102.96 36.785 104.01 ;
      RECT MASK 1 36.999 102.96 37.059 104.01 ;
      RECT MASK 1 37.273 102.96 37.333 104.01 ;
      RECT MASK 1 37.547 102.96 37.607 104.01 ;
      RECT MASK 1 37.821 102.96 37.881 104.01 ;
      RECT MASK 1 38.095 102.96 38.155 104.01 ;
      RECT MASK 1 38.369 102.96 38.429 104.01 ;
      RECT MASK 1 38.643 102.96 38.703 104.01 ;
      RECT MASK 1 38.917 102.96 38.977 104.01 ;
      RECT MASK 1 39.191 102.96 39.251 104.01 ;
      RECT MASK 1 39.465 102.96 39.525 104.01 ;
      RECT MASK 1 39.739 102.96 39.799 104.01 ;
      RECT MASK 1 40.013 102.96 40.073 104.01 ;
      RECT MASK 1 40.287 102.96 40.347 104.01 ;
      RECT MASK 1 40.561 102.96 40.621 104.01 ;
      RECT MASK 1 40.835 102.96 40.895 104.01 ;
      RECT MASK 1 41.109 102.96 41.169 104.01 ;
      RECT MASK 1 41.383 102.96 41.443 104.01 ;
      RECT MASK 1 41.657 102.96 41.717 104.01 ;
      RECT MASK 1 41.931 102.96 41.991 104.01 ;
      RECT MASK 1 42.205 102.96 42.265 104.01 ;
      RECT MASK 1 42.479 102.96 42.539 104.01 ;
      RECT MASK 1 42.753 102.96 42.813 104.01 ;
      RECT MASK 1 43.027 102.96 43.087 104.01 ;
      RECT MASK 1 43.301 102.96 43.361 104.01 ;
      RECT MASK 1 43.575 102.96 43.635 104.01 ;
      RECT MASK 1 45.593 102.96 45.653 104.01 ;
      RECT MASK 1 45.867 102.96 45.927 104.01 ;
      RECT MASK 1 46.141 102.96 46.201 104.01 ;
      RECT MASK 1 46.415 102.96 46.475 104.01 ;
      RECT MASK 1 46.689 102.96 46.749 104.01 ;
      RECT MASK 1 46.963 102.96 47.023 104.01 ;
      RECT MASK 1 47.237 102.96 47.297 104.01 ;
      RECT MASK 1 47.511 102.96 47.571 104.01 ;
      RECT MASK 1 47.785 102.96 47.845 104.01 ;
      RECT MASK 1 48.059 102.96 48.119 104.01 ;
      RECT MASK 1 48.333 102.96 48.393 104.01 ;
      RECT MASK 1 48.607 102.96 48.667 104.01 ;
      RECT MASK 1 48.881 102.96 48.941 104.01 ;
      RECT MASK 1 49.155 102.96 49.215 104.01 ;
      RECT MASK 1 49.429 102.96 49.489 104.01 ;
      RECT MASK 1 49.703 102.96 49.763 104.01 ;
      RECT MASK 1 49.977 102.96 50.037 104.01 ;
      RECT MASK 1 50.251 102.96 50.311 104.01 ;
      RECT MASK 1 50.525 102.96 50.585 104.01 ;
      RECT MASK 1 50.799 102.96 50.859 104.01 ;
      RECT MASK 1 51.073 102.96 51.133 104.01 ;
      RECT MASK 1 51.347 102.96 51.407 104.01 ;
      RECT MASK 1 51.621 102.96 51.681 104.01 ;
      RECT MASK 1 51.895 102.96 51.955 104.01 ;
      RECT MASK 1 52.169 102.96 52.229 104.01 ;
      RECT MASK 1 52.443 102.96 52.503 104.01 ;
      RECT MASK 1 52.717 102.96 52.777 104.01 ;
      RECT MASK 1 52.991 102.96 53.051 104.01 ;
      RECT MASK 1 53.265 102.96 53.325 104.01 ;
      RECT MASK 1 53.539 102.96 53.599 104.01 ;
      RECT MASK 1 53.813 102.96 53.873 104.01 ;
      RECT MASK 1 54.087 102.96 54.147 104.01 ;
      RECT MASK 1 54.361 102.96 54.421 104.01 ;
      RECT MASK 1 54.635 102.96 54.695 104.01 ;
      RECT MASK 1 54.909 102.96 54.969 104.01 ;
      RECT MASK 1 55.183 102.96 55.243 104.01 ;
      RECT MASK 1 55.457 102.96 55.517 104.01 ;
      RECT MASK 1 55.731 102.96 55.791 104.01 ;
      RECT MASK 1 56.005 102.96 56.065 104.01 ;
      RECT MASK 1 56.279 102.96 56.339 104.01 ;
      RECT MASK 1 56.553 102.96 56.613 104.01 ;
      RECT MASK 1 56.827 102.96 56.887 104.01 ;
      RECT MASK 1 57.101 102.96 57.161 104.01 ;
      RECT MASK 1 57.375 102.96 57.435 104.01 ;
      RECT MASK 1 57.649 102.96 57.709 104.01 ;
      RECT MASK 1 57.923 102.96 57.983 104.01 ;
      RECT MASK 1 58.197 102.96 58.257 104.01 ;
      RECT MASK 1 58.471 102.96 58.531 104.01 ;
      RECT MASK 1 58.745 102.96 58.805 104.01 ;
      RECT MASK 1 59.019 102.96 59.079 104.01 ;
      RECT MASK 1 59.293 102.96 59.353 104.01 ;
      RECT MASK 1 59.567 102.96 59.627 104.01 ;
      RECT MASK 1 59.841 102.96 59.901 104.01 ;
      RECT MASK 1 60.115 102.96 60.175 104.01 ;
      RECT MASK 1 60.389 102.96 60.449 104.01 ;
      RECT MASK 1 60.663 102.96 60.723 104.01 ;
      RECT MASK 1 60.937 102.96 60.997 104.01 ;
      RECT MASK 1 61.211 102.96 61.271 104.01 ;
      RECT MASK 1 61.485 102.96 61.545 104.01 ;
      RECT MASK 1 61.759 102.96 61.819 104.01 ;
      RECT MASK 1 62.033 102.96 62.093 104.01 ;
      RECT MASK 1 62.307 102.96 62.367 104.01 ;
      RECT MASK 1 62.581 102.96 62.641 104.01 ;
      RECT MASK 1 62.855 102.96 62.915 104.01 ;
      RECT MASK 1 63.129 102.96 63.189 104.01 ;
      RECT MASK 1 63.403 102.96 63.463 104.01 ;
      RECT MASK 1 63.677 102.96 63.737 104.01 ;
      RECT MASK 1 63.951 102.96 64.011 104.01 ;
      RECT MASK 1 64.225 102.96 64.285 104.01 ;
      RECT MASK 1 64.499 102.96 64.559 104.01 ;
      RECT MASK 1 64.773 102.96 64.833 104.01 ;
      RECT MASK 1 65.047 102.96 65.107 104.01 ;
      RECT MASK 1 65.321 102.96 65.381 104.01 ;
      RECT MASK 1 65.595 102.96 65.655 104.01 ;
      RECT MASK 1 65.869 102.96 65.929 104.01 ;
      RECT MASK 1 66.143 102.96 66.203 104.01 ;
      RECT MASK 1 66.417 102.96 66.477 104.01 ;
      RECT MASK 1 66.691 102.96 66.751 104.01 ;
      RECT MASK 1 66.965 102.96 67.025 104.01 ;
      RECT MASK 1 67.239 102.96 67.299 104.01 ;
      RECT MASK 1 67.513 102.96 67.573 104.01 ;
      RECT MASK 1 67.787 102.96 67.847 104.01 ;
      RECT MASK 1 68.061 102.96 68.121 104.01 ;
      RECT MASK 1 68.335 102.96 68.395 104.01 ;
      RECT MASK 1 68.609 102.96 68.669 104.01 ;
      RECT MASK 1 68.883 102.96 68.943 104.01 ;
      RECT MASK 1 69.157 102.96 69.217 104.01 ;
      RECT MASK 1 69.431 102.96 69.491 104.01 ;
      RECT MASK 1 69.705 102.96 69.765 104.01 ;
      RECT MASK 1 69.979 102.96 70.039 104.01 ;
      RECT MASK 1 70.253 102.96 70.313 104.01 ;
      RECT MASK 1 70.527 102.96 70.587 104.01 ;
      RECT MASK 1 70.801 102.96 70.861 104.01 ;
      RECT MASK 1 71.075 102.96 71.135 104.01 ;
      RECT MASK 1 71.349 102.96 71.409 104.01 ;
      RECT MASK 1 71.623 102.96 71.683 104.01 ;
      RECT MASK 1 71.897 102.96 71.957 104.01 ;
      RECT MASK 1 72.171 102.96 72.231 104.01 ;
      RECT MASK 1 72.445 102.96 72.505 104.01 ;
      RECT MASK 1 72.719 102.96 72.779 104.01 ;
      RECT MASK 1 72.993 102.96 73.053 104.01 ;
      RECT MASK 1 73.267 102.96 73.327 104.01 ;
      RECT MASK 1 73.541 102.96 73.601 104.01 ;
      RECT MASK 1 73.815 102.96 73.875 104.01 ;
      RECT MASK 1 74.089 102.96 74.149 104.01 ;
      RECT MASK 1 74.363 102.96 74.423 104.01 ;
      RECT MASK 1 74.637 102.96 74.697 104.01 ;
      RECT MASK 1 74.911 102.96 74.971 104.01 ;
      RECT MASK 1 75.185 102.96 75.245 104.01 ;
      RECT MASK 1 75.459 102.96 75.519 104.01 ;
      RECT MASK 1 75.733 102.96 75.793 104.01 ;
      RECT MASK 1 76.007 102.96 76.067 104.01 ;
      RECT MASK 1 76.281 102.96 76.341 104.01 ;
      RECT MASK 1 76.555 102.96 76.615 104.01 ;
      RECT MASK 1 76.829 102.96 76.889 104.01 ;
      RECT MASK 1 77.103 102.96 77.163 104.01 ;
      RECT MASK 1 77.377 102.96 77.437 104.01 ;
      RECT MASK 1 77.651 102.96 77.711 104.01 ;
      RECT MASK 1 77.925 102.96 77.985 104.01 ;
      RECT MASK 1 78.199 102.96 78.259 104.01 ;
      RECT MASK 1 78.473 102.96 78.533 104.01 ;
      RECT MASK 1 78.747 102.96 78.807 104.01 ;
      RECT MASK 1 79.021 102.96 79.081 104.01 ;
      RECT MASK 1 79.295 102.96 79.355 104.01 ;
      RECT MASK 1 79.569 102.96 79.629 104.01 ;
      RECT MASK 1 79.843 102.96 79.903 104.01 ;
      RECT MASK 1 80.117 102.96 80.177 104.01 ;
      RECT MASK 1 80.391 102.96 80.451 104.01 ;
      RECT MASK 1 80.665 102.96 80.725 104.01 ;
      RECT MASK 1 80.939 102.96 80.999 104.01 ;
      RECT MASK 1 81.213 102.96 81.273 104.01 ;
      RECT MASK 1 81.487 102.96 81.547 104.01 ;
      RECT MASK 1 81.761 102.96 81.821 104.01 ;
      RECT MASK 1 82.035 102.96 82.095 104.01 ;
      RECT MASK 1 82.309 102.96 82.369 104.01 ;
      RECT MASK 1 82.583 102.96 82.643 104.01 ;
      RECT MASK 1 82.857 102.96 82.917 104.01 ;
      RECT MASK 1 83.131 102.96 83.191 104.01 ;
      RECT MASK 1 83.405 102.96 83.465 104.01 ;
      RECT MASK 1 83.679 102.96 83.739 104.01 ;
      RECT MASK 1 83.953 102.96 84.013 104.01 ;
      RECT MASK 1 84.227 102.96 84.287 104.01 ;
      RECT MASK 1 84.501 102.96 84.561 104.01 ;
      RECT MASK 1 84.775 102.96 84.835 104.01 ;
      RECT MASK 1 85.049 102.96 85.109 104.01 ;
      RECT MASK 1 85.323 102.96 85.383 104.01 ;
      RECT MASK 1 85.597 102.96 85.657 104.01 ;
      RECT MASK 1 85.871 102.96 85.931 104.01 ;
      RECT MASK 1 86.145 102.96 86.205 104.01 ;
      RECT MASK 1 86.419 102.96 86.479 104.01 ;
      RECT MASK 1 86.693 102.96 86.753 104.01 ;
      RECT MASK 1 86.967 102.96 87.027 104.01 ;
      RECT MASK 1 88.952 102.96 89.012 104.01 ;
      RECT MASK 1 89.226 102.96 89.286 104.01 ;
      RECT MASK 1 89.5 102.96 89.56 104.01 ;
      RECT MASK 1 89.774 102.96 89.834 104.01 ;
      RECT MASK 1 90.048 102.96 90.108 104.01 ;
      RECT MASK 1 90.322 102.96 90.382 104.01 ;
      RECT MASK 1 90.596 102.96 90.656 104.01 ;
      RECT MASK 1 90.87 102.96 90.93 104.01 ;
      RECT MASK 1 91.144 102.96 91.204 104.01 ;
      RECT MASK 1 91.418 102.96 91.478 104.01 ;
      RECT MASK 1 91.692 102.96 91.752 104.01 ;
      RECT MASK 1 91.966 102.96 92.026 104.01 ;
      RECT MASK 1 92.24 102.96 92.3 104.01 ;
      RECT MASK 1 92.514 102.96 92.574 104.01 ;
      RECT MASK 1 92.788 102.96 92.848 104.01 ;
      RECT MASK 1 93.062 102.96 93.122 104.01 ;
      RECT MASK 1 93.336 102.96 93.396 104.01 ;
      RECT MASK 1 93.61 102.96 93.67 104.01 ;
      RECT MASK 1 93.884 102.96 93.944 104.01 ;
      RECT MASK 1 94.158 102.96 94.218 104.01 ;
      RECT MASK 1 94.432 102.96 94.492 104.01 ;
      RECT MASK 1 94.706 102.96 94.766 104.01 ;
      RECT MASK 1 94.98 102.96 95.04 104.01 ;
      RECT MASK 1 95.254 102.96 95.314 104.01 ;
      RECT MASK 1 95.528 102.96 95.588 104.01 ;
      RECT MASK 1 95.802 102.96 95.862 104.01 ;
      RECT MASK 1 96.076 102.96 96.136 104.01 ;
      RECT MASK 1 96.35 102.96 96.41 104.01 ;
      RECT MASK 1 96.624 102.96 96.684 104.01 ;
      RECT MASK 1 96.898 102.96 96.958 104.01 ;
      RECT MASK 1 97.172 102.96 97.232 104.01 ;
      RECT MASK 1 97.446 102.96 97.506 104.01 ;
      RECT MASK 1 97.72 102.96 97.78 104.01 ;
      RECT MASK 1 97.994 102.96 98.054 104.01 ;
      RECT MASK 1 98.268 102.96 98.328 104.01 ;
      RECT MASK 1 98.542 102.96 98.602 104.01 ;
      RECT MASK 1 98.816 102.96 98.876 104.01 ;
      RECT MASK 1 99.09 102.96 99.15 104.01 ;
      RECT MASK 1 99.364 102.96 99.424 104.01 ;
      RECT MASK 1 99.638 102.96 99.698 104.01 ;
      RECT MASK 1 99.912 102.96 99.972 104.01 ;
      RECT MASK 1 100.186 102.96 100.246 104.01 ;
      RECT MASK 1 100.46 102.96 100.52 104.01 ;
      RECT MASK 1 100.734 102.96 100.794 104.01 ;
      RECT MASK 1 101.008 102.96 101.068 104.01 ;
      RECT MASK 1 101.282 102.96 101.342 104.01 ;
      RECT MASK 1 101.556 102.96 101.616 104.01 ;
      RECT MASK 1 101.83 102.96 101.89 104.01 ;
      RECT MASK 1 102.104 102.96 102.164 104.01 ;
      RECT MASK 1 102.378 102.96 102.438 104.01 ;
      RECT MASK 1 102.652 102.96 102.712 104.01 ;
      RECT MASK 1 102.926 102.96 102.986 104.01 ;
      RECT MASK 1 103.2 102.96 103.26 104.01 ;
      RECT MASK 1 103.474 102.96 103.534 104.01 ;
      RECT MASK 1 103.748 102.96 103.808 104.01 ;
      RECT MASK 1 104.022 102.96 104.082 104.01 ;
      RECT MASK 1 104.296 102.96 104.356 104.01 ;
      RECT MASK 1 104.57 102.96 104.63 104.01 ;
      RECT MASK 1 104.844 102.96 104.904 104.01 ;
      RECT MASK 1 105.118 102.96 105.178 104.01 ;
      RECT MASK 1 105.392 102.96 105.452 104.01 ;
      RECT MASK 1 105.666 102.96 105.726 104.01 ;
      RECT MASK 1 105.94 102.96 106 104.01 ;
      RECT MASK 1 106.214 102.96 106.274 104.01 ;
      RECT MASK 1 106.488 102.96 106.548 104.01 ;
      RECT MASK 1 106.762 102.96 106.822 104.01 ;
      RECT MASK 1 107.036 102.96 107.096 104.01 ;
      RECT MASK 1 107.31 102.96 107.37 104.01 ;
      RECT MASK 1 107.584 102.96 107.644 104.01 ;
      RECT MASK 1 107.858 102.96 107.918 104.01 ;
      RECT MASK 1 108.132 102.96 108.192 104.01 ;
      RECT MASK 1 108.406 102.96 108.466 104.01 ;
      RECT MASK 1 108.68 102.96 108.74 104.01 ;
      RECT MASK 1 108.954 102.96 109.014 104.01 ;
      RECT MASK 1 109.228 102.96 109.288 104.01 ;
      RECT MASK 1 109.502 102.96 109.562 104.01 ;
      RECT MASK 1 109.776 102.96 109.836 104.01 ;
      RECT MASK 1 110.05 102.96 110.11 104.01 ;
      RECT MASK 1 110.324 102.96 110.384 104.01 ;
      RECT MASK 1 110.598 102.96 110.658 104.01 ;
      RECT MASK 1 110.872 102.96 110.932 104.01 ;
      RECT MASK 1 111.146 102.96 111.206 104.01 ;
      RECT MASK 1 111.42 102.96 111.48 104.01 ;
      RECT MASK 1 111.694 102.96 111.754 104.01 ;
      RECT MASK 1 111.968 102.96 112.028 104.01 ;
      RECT MASK 1 112.242 102.96 112.302 104.01 ;
      RECT MASK 1 112.516 102.96 112.576 104.01 ;
      RECT MASK 1 112.79 102.96 112.85 104.01 ;
      RECT MASK 1 113.064 102.96 113.124 104.01 ;
      RECT MASK 1 113.338 102.96 113.398 104.01 ;
      RECT MASK 1 113.612 102.96 113.672 104.01 ;
      RECT MASK 1 113.886 102.96 113.946 104.01 ;
      RECT MASK 1 114.16 102.96 114.22 104.01 ;
      RECT MASK 1 114.434 102.96 114.494 104.01 ;
      RECT MASK 1 114.708 102.96 114.768 104.01 ;
      RECT MASK 1 114.982 102.96 115.042 104.01 ;
      RECT MASK 1 115.256 102.96 115.316 104.01 ;
      RECT MASK 1 115.53 102.96 115.59 104.01 ;
      RECT MASK 1 115.804 102.96 115.864 104.01 ;
      RECT MASK 1 116.078 102.96 116.138 104.01 ;
      RECT MASK 1 116.352 102.96 116.412 104.01 ;
      RECT MASK 1 116.626 102.96 116.686 104.01 ;
      RECT MASK 1 116.9 102.96 116.96 104.01 ;
      RECT MASK 1 117.174 102.96 117.234 104.01 ;
      RECT MASK 1 117.448 102.96 117.508 104.01 ;
      RECT MASK 1 117.722 102.96 117.782 104.01 ;
      RECT MASK 1 117.996 102.96 118.056 104.01 ;
      RECT MASK 1 118.27 102.96 118.33 104.01 ;
      RECT MASK 1 118.544 102.96 118.604 104.01 ;
      RECT MASK 1 118.818 102.96 118.878 104.01 ;
      RECT MASK 1 119.092 102.96 119.152 104.01 ;
      RECT MASK 1 119.366 102.96 119.426 104.01 ;
      RECT MASK 1 119.64 102.96 119.7 104.01 ;
      RECT MASK 1 119.914 102.96 119.974 104.01 ;
      RECT MASK 1 120.188 102.96 120.248 104.01 ;
      RECT MASK 1 120.462 102.96 120.522 104.01 ;
      RECT MASK 1 120.736 102.96 120.796 104.01 ;
      RECT MASK 1 121.01 102.96 121.07 104.01 ;
      RECT MASK 1 121.284 102.96 121.344 104.01 ;
      RECT MASK 1 121.558 102.96 121.618 104.01 ;
      RECT MASK 1 121.832 102.96 121.892 104.01 ;
      RECT MASK 1 122.106 102.96 122.166 104.01 ;
      RECT MASK 1 122.38 102.96 122.44 104.01 ;
      RECT MASK 1 122.654 102.96 122.714 104.01 ;
      RECT MASK 1 122.928 102.96 122.988 104.01 ;
      RECT MASK 1 123.202 102.96 123.262 104.01 ;
      RECT MASK 1 123.476 102.96 123.536 104.01 ;
      RECT MASK 1 123.75 102.96 123.81 104.01 ;
      RECT MASK 1 124.024 102.96 124.084 104.01 ;
      RECT MASK 1 124.298 102.96 124.358 104.01 ;
      RECT MASK 1 124.572 102.96 124.632 104.01 ;
      RECT MASK 1 124.846 102.96 124.906 104.01 ;
      RECT MASK 1 125.12 102.96 125.18 104.01 ;
      RECT MASK 1 125.394 102.96 125.454 104.01 ;
      RECT MASK 1 125.668 102.96 125.728 104.01 ;
      RECT MASK 1 125.942 102.96 126.002 104.01 ;
      RECT MASK 1 126.216 102.96 126.276 104.01 ;
      RECT MASK 1 126.49 102.96 126.55 104.01 ;
      RECT MASK 1 126.764 102.96 126.824 104.01 ;
      RECT MASK 1 127.038 102.96 127.098 104.01 ;
      RECT MASK 1 127.312 102.96 127.372 104.01 ;
      RECT MASK 1 127.586 102.96 127.646 104.01 ;
      RECT MASK 1 2.201 104.67 2.261 105.72 ;
      RECT MASK 1 2.475 104.67 2.535 105.72 ;
      RECT MASK 1 2.749 104.67 2.809 105.72 ;
      RECT MASK 1 3.023 104.67 3.083 105.72 ;
      RECT MASK 1 3.297 104.67 3.357 105.72 ;
      RECT MASK 1 3.571 104.67 3.631 105.72 ;
      RECT MASK 1 3.845 104.67 3.905 105.72 ;
      RECT MASK 1 4.119 104.67 4.179 105.72 ;
      RECT MASK 1 4.393 104.67 4.453 105.72 ;
      RECT MASK 1 4.667 104.67 4.727 105.72 ;
      RECT MASK 1 4.941 104.67 5.001 105.72 ;
      RECT MASK 1 5.215 104.67 5.275 105.72 ;
      RECT MASK 1 5.489 104.67 5.549 105.72 ;
      RECT MASK 1 5.763 104.67 5.823 105.72 ;
      RECT MASK 1 6.037 104.67 6.097 105.72 ;
      RECT MASK 1 6.311 104.67 6.371 105.72 ;
      RECT MASK 1 6.585 104.67 6.645 105.72 ;
      RECT MASK 1 6.859 104.67 6.919 105.72 ;
      RECT MASK 1 7.133 104.67 7.193 105.72 ;
      RECT MASK 1 7.407 104.67 7.467 105.72 ;
      RECT MASK 1 7.681 104.67 7.741 105.72 ;
      RECT MASK 1 7.955 104.67 8.015 105.72 ;
      RECT MASK 1 8.229 104.67 8.289 105.72 ;
      RECT MASK 1 8.503 104.67 8.563 105.72 ;
      RECT MASK 1 8.777 104.67 8.837 105.72 ;
      RECT MASK 1 9.051 104.67 9.111 105.72 ;
      RECT MASK 1 9.325 104.67 9.385 105.72 ;
      RECT MASK 1 9.599 104.67 9.659 105.72 ;
      RECT MASK 1 9.873 104.67 9.933 105.72 ;
      RECT MASK 1 10.147 104.67 10.207 105.72 ;
      RECT MASK 1 10.421 104.67 10.481 105.72 ;
      RECT MASK 1 10.695 104.67 10.755 105.72 ;
      RECT MASK 1 10.969 104.67 11.029 105.72 ;
      RECT MASK 1 11.243 104.67 11.303 105.72 ;
      RECT MASK 1 11.517 104.67 11.577 105.72 ;
      RECT MASK 1 11.791 104.67 11.851 105.72 ;
      RECT MASK 1 12.065 104.67 12.125 105.72 ;
      RECT MASK 1 12.339 104.67 12.399 105.72 ;
      RECT MASK 1 12.613 104.67 12.673 105.72 ;
      RECT MASK 1 12.887 104.67 12.947 105.72 ;
      RECT MASK 1 13.161 104.67 13.221 105.72 ;
      RECT MASK 1 13.435 104.67 13.495 105.72 ;
      RECT MASK 1 13.709 104.67 13.769 105.72 ;
      RECT MASK 1 13.983 104.67 14.043 105.72 ;
      RECT MASK 1 14.257 104.67 14.317 105.72 ;
      RECT MASK 1 14.531 104.67 14.591 105.72 ;
      RECT MASK 1 14.805 104.67 14.865 105.72 ;
      RECT MASK 1 15.079 104.67 15.139 105.72 ;
      RECT MASK 1 15.353 104.67 15.413 105.72 ;
      RECT MASK 1 15.627 104.67 15.687 105.72 ;
      RECT MASK 1 15.901 104.67 15.961 105.72 ;
      RECT MASK 1 16.175 104.67 16.235 105.72 ;
      RECT MASK 1 16.449 104.67 16.509 105.72 ;
      RECT MASK 1 16.723 104.67 16.783 105.72 ;
      RECT MASK 1 16.997 104.67 17.057 105.72 ;
      RECT MASK 1 17.271 104.67 17.331 105.72 ;
      RECT MASK 1 17.545 104.67 17.605 105.72 ;
      RECT MASK 1 17.819 104.67 17.879 105.72 ;
      RECT MASK 1 18.093 104.67 18.153 105.72 ;
      RECT MASK 1 18.367 104.67 18.427 105.72 ;
      RECT MASK 1 18.641 104.67 18.701 105.72 ;
      RECT MASK 1 18.915 104.67 18.975 105.72 ;
      RECT MASK 1 19.189 104.67 19.249 105.72 ;
      RECT MASK 1 19.463 104.67 19.523 105.72 ;
      RECT MASK 1 19.737 104.67 19.797 105.72 ;
      RECT MASK 1 20.011 104.67 20.071 105.72 ;
      RECT MASK 1 20.285 104.67 20.345 105.72 ;
      RECT MASK 1 20.559 104.67 20.619 105.72 ;
      RECT MASK 1 20.833 104.67 20.893 105.72 ;
      RECT MASK 1 21.107 104.67 21.167 105.72 ;
      RECT MASK 1 21.381 104.67 21.441 105.72 ;
      RECT MASK 1 21.655 104.67 21.715 105.72 ;
      RECT MASK 1 21.929 104.67 21.989 105.72 ;
      RECT MASK 1 22.203 104.67 22.263 105.72 ;
      RECT MASK 1 22.477 104.67 22.537 105.72 ;
      RECT MASK 1 22.751 104.67 22.811 105.72 ;
      RECT MASK 1 23.025 104.67 23.085 105.72 ;
      RECT MASK 1 23.299 104.67 23.359 105.72 ;
      RECT MASK 1 23.573 104.67 23.633 105.72 ;
      RECT MASK 1 23.847 104.67 23.907 105.72 ;
      RECT MASK 1 24.121 104.67 24.181 105.72 ;
      RECT MASK 1 24.395 104.67 24.455 105.72 ;
      RECT MASK 1 24.669 104.67 24.729 105.72 ;
      RECT MASK 1 24.943 104.67 25.003 105.72 ;
      RECT MASK 1 25.217 104.67 25.277 105.72 ;
      RECT MASK 1 25.491 104.67 25.551 105.72 ;
      RECT MASK 1 25.765 104.67 25.825 105.72 ;
      RECT MASK 1 26.039 104.67 26.099 105.72 ;
      RECT MASK 1 26.313 104.67 26.373 105.72 ;
      RECT MASK 1 26.587 104.67 26.647 105.72 ;
      RECT MASK 1 26.861 104.67 26.921 105.72 ;
      RECT MASK 1 27.135 104.67 27.195 105.72 ;
      RECT MASK 1 27.409 104.67 27.469 105.72 ;
      RECT MASK 1 27.683 104.67 27.743 105.72 ;
      RECT MASK 1 27.957 104.67 28.017 105.72 ;
      RECT MASK 1 28.231 104.67 28.291 105.72 ;
      RECT MASK 1 28.505 104.67 28.565 105.72 ;
      RECT MASK 1 28.779 104.67 28.839 105.72 ;
      RECT MASK 1 29.053 104.67 29.113 105.72 ;
      RECT MASK 1 29.327 104.67 29.387 105.72 ;
      RECT MASK 1 29.601 104.67 29.661 105.72 ;
      RECT MASK 1 29.875 104.67 29.935 105.72 ;
      RECT MASK 1 30.149 104.67 30.209 105.72 ;
      RECT MASK 1 30.423 104.67 30.483 105.72 ;
      RECT MASK 1 30.697 104.67 30.757 105.72 ;
      RECT MASK 1 30.971 104.67 31.031 105.72 ;
      RECT MASK 1 31.245 104.67 31.305 105.72 ;
      RECT MASK 1 31.519 104.67 31.579 105.72 ;
      RECT MASK 1 31.793 104.67 31.853 105.72 ;
      RECT MASK 1 32.067 104.67 32.127 105.72 ;
      RECT MASK 1 32.341 104.67 32.401 105.72 ;
      RECT MASK 1 32.615 104.67 32.675 105.72 ;
      RECT MASK 1 32.889 104.67 32.949 105.72 ;
      RECT MASK 1 33.163 104.67 33.223 105.72 ;
      RECT MASK 1 33.437 104.67 33.497 105.72 ;
      RECT MASK 1 33.711 104.67 33.771 105.72 ;
      RECT MASK 1 33.985 104.67 34.045 105.72 ;
      RECT MASK 1 34.259 104.67 34.319 105.72 ;
      RECT MASK 1 34.533 104.67 34.593 105.72 ;
      RECT MASK 1 34.807 104.67 34.867 105.72 ;
      RECT MASK 1 35.081 104.67 35.141 105.72 ;
      RECT MASK 1 35.355 104.67 35.415 105.72 ;
      RECT MASK 1 35.629 104.67 35.689 105.72 ;
      RECT MASK 1 35.903 104.67 35.963 105.72 ;
      RECT MASK 1 36.177 104.67 36.237 105.72 ;
      RECT MASK 1 36.451 104.67 36.511 105.72 ;
      RECT MASK 1 36.725 104.67 36.785 105.72 ;
      RECT MASK 1 36.999 104.67 37.059 105.72 ;
      RECT MASK 1 37.273 104.67 37.333 105.72 ;
      RECT MASK 1 37.547 104.67 37.607 105.72 ;
      RECT MASK 1 37.821 104.67 37.881 105.72 ;
      RECT MASK 1 38.095 104.67 38.155 105.72 ;
      RECT MASK 1 38.369 104.67 38.429 105.72 ;
      RECT MASK 1 38.643 104.67 38.703 105.72 ;
      RECT MASK 1 38.917 104.67 38.977 105.72 ;
      RECT MASK 1 39.191 104.67 39.251 105.72 ;
      RECT MASK 1 39.465 104.67 39.525 105.72 ;
      RECT MASK 1 39.739 104.67 39.799 105.72 ;
      RECT MASK 1 40.013 104.67 40.073 105.72 ;
      RECT MASK 1 40.287 104.67 40.347 105.72 ;
      RECT MASK 1 40.561 104.67 40.621 105.72 ;
      RECT MASK 1 40.835 104.67 40.895 105.72 ;
      RECT MASK 1 41.109 104.67 41.169 105.72 ;
      RECT MASK 1 41.383 104.67 41.443 105.72 ;
      RECT MASK 1 41.657 104.67 41.717 105.72 ;
      RECT MASK 1 41.931 104.67 41.991 105.72 ;
      RECT MASK 1 42.205 104.67 42.265 105.72 ;
      RECT MASK 1 42.479 104.67 42.539 105.72 ;
      RECT MASK 1 42.753 104.67 42.813 105.72 ;
      RECT MASK 1 43.027 104.67 43.087 105.72 ;
      RECT MASK 1 43.301 104.67 43.361 105.72 ;
      RECT MASK 1 43.575 104.67 43.635 105.72 ;
      RECT MASK 1 45.593 104.67 45.653 105.72 ;
      RECT MASK 1 45.867 104.67 45.927 105.72 ;
      RECT MASK 1 46.141 104.67 46.201 105.72 ;
      RECT MASK 1 46.415 104.67 46.475 105.72 ;
      RECT MASK 1 46.689 104.67 46.749 105.72 ;
      RECT MASK 1 46.963 104.67 47.023 105.72 ;
      RECT MASK 1 47.237 104.67 47.297 105.72 ;
      RECT MASK 1 47.511 104.67 47.571 105.72 ;
      RECT MASK 1 47.785 104.67 47.845 105.72 ;
      RECT MASK 1 48.059 104.67 48.119 105.72 ;
      RECT MASK 1 48.333 104.67 48.393 105.72 ;
      RECT MASK 1 48.607 104.67 48.667 105.72 ;
      RECT MASK 1 48.881 104.67 48.941 105.72 ;
      RECT MASK 1 49.155 104.67 49.215 105.72 ;
      RECT MASK 1 49.429 104.67 49.489 105.72 ;
      RECT MASK 1 49.703 104.67 49.763 105.72 ;
      RECT MASK 1 49.977 104.67 50.037 105.72 ;
      RECT MASK 1 50.251 104.67 50.311 105.72 ;
      RECT MASK 1 50.525 104.67 50.585 105.72 ;
      RECT MASK 1 50.799 104.67 50.859 105.72 ;
      RECT MASK 1 51.073 104.67 51.133 105.72 ;
      RECT MASK 1 51.347 104.67 51.407 105.72 ;
      RECT MASK 1 51.621 104.67 51.681 105.72 ;
      RECT MASK 1 51.895 104.67 51.955 105.72 ;
      RECT MASK 1 52.169 104.67 52.229 105.72 ;
      RECT MASK 1 52.443 104.67 52.503 105.72 ;
      RECT MASK 1 52.717 104.67 52.777 105.72 ;
      RECT MASK 1 52.991 104.67 53.051 105.72 ;
      RECT MASK 1 53.265 104.67 53.325 105.72 ;
      RECT MASK 1 53.539 104.67 53.599 105.72 ;
      RECT MASK 1 53.813 104.67 53.873 105.72 ;
      RECT MASK 1 54.087 104.67 54.147 105.72 ;
      RECT MASK 1 54.361 104.67 54.421 105.72 ;
      RECT MASK 1 54.635 104.67 54.695 105.72 ;
      RECT MASK 1 54.909 104.67 54.969 105.72 ;
      RECT MASK 1 55.183 104.67 55.243 105.72 ;
      RECT MASK 1 55.457 104.67 55.517 105.72 ;
      RECT MASK 1 55.731 104.67 55.791 105.72 ;
      RECT MASK 1 56.005 104.67 56.065 105.72 ;
      RECT MASK 1 56.279 104.67 56.339 105.72 ;
      RECT MASK 1 56.553 104.67 56.613 105.72 ;
      RECT MASK 1 56.827 104.67 56.887 105.72 ;
      RECT MASK 1 57.101 104.67 57.161 105.72 ;
      RECT MASK 1 57.375 104.67 57.435 105.72 ;
      RECT MASK 1 57.649 104.67 57.709 105.72 ;
      RECT MASK 1 57.923 104.67 57.983 105.72 ;
      RECT MASK 1 58.197 104.67 58.257 105.72 ;
      RECT MASK 1 58.471 104.67 58.531 105.72 ;
      RECT MASK 1 58.745 104.67 58.805 105.72 ;
      RECT MASK 1 59.019 104.67 59.079 105.72 ;
      RECT MASK 1 59.293 104.67 59.353 105.72 ;
      RECT MASK 1 59.567 104.67 59.627 105.72 ;
      RECT MASK 1 59.841 104.67 59.901 105.72 ;
      RECT MASK 1 60.115 104.67 60.175 105.72 ;
      RECT MASK 1 60.389 104.67 60.449 105.72 ;
      RECT MASK 1 60.663 104.67 60.723 105.72 ;
      RECT MASK 1 60.937 104.67 60.997 105.72 ;
      RECT MASK 1 61.211 104.67 61.271 105.72 ;
      RECT MASK 1 61.485 104.67 61.545 105.72 ;
      RECT MASK 1 61.759 104.67 61.819 105.72 ;
      RECT MASK 1 62.033 104.67 62.093 105.72 ;
      RECT MASK 1 62.307 104.67 62.367 105.72 ;
      RECT MASK 1 62.581 104.67 62.641 105.72 ;
      RECT MASK 1 62.855 104.67 62.915 105.72 ;
      RECT MASK 1 63.129 104.67 63.189 105.72 ;
      RECT MASK 1 63.403 104.67 63.463 105.72 ;
      RECT MASK 1 63.677 104.67 63.737 105.72 ;
      RECT MASK 1 63.951 104.67 64.011 105.72 ;
      RECT MASK 1 64.225 104.67 64.285 105.72 ;
      RECT MASK 1 64.499 104.67 64.559 105.72 ;
      RECT MASK 1 64.773 104.67 64.833 105.72 ;
      RECT MASK 1 65.047 104.67 65.107 105.72 ;
      RECT MASK 1 65.321 104.67 65.381 105.72 ;
      RECT MASK 1 65.595 104.67 65.655 105.72 ;
      RECT MASK 1 65.869 104.67 65.929 105.72 ;
      RECT MASK 1 66.143 104.67 66.203 105.72 ;
      RECT MASK 1 66.417 104.67 66.477 105.72 ;
      RECT MASK 1 66.691 104.67 66.751 105.72 ;
      RECT MASK 1 66.965 104.67 67.025 105.72 ;
      RECT MASK 1 67.239 104.67 67.299 105.72 ;
      RECT MASK 1 67.513 104.67 67.573 105.72 ;
      RECT MASK 1 67.787 104.67 67.847 105.72 ;
      RECT MASK 1 68.061 104.67 68.121 105.72 ;
      RECT MASK 1 68.335 104.67 68.395 105.72 ;
      RECT MASK 1 68.609 104.67 68.669 105.72 ;
      RECT MASK 1 68.883 104.67 68.943 105.72 ;
      RECT MASK 1 69.157 104.67 69.217 105.72 ;
      RECT MASK 1 69.431 104.67 69.491 105.72 ;
      RECT MASK 1 69.705 104.67 69.765 105.72 ;
      RECT MASK 1 69.979 104.67 70.039 105.72 ;
      RECT MASK 1 70.253 104.67 70.313 105.72 ;
      RECT MASK 1 70.527 104.67 70.587 105.72 ;
      RECT MASK 1 70.801 104.67 70.861 105.72 ;
      RECT MASK 1 71.075 104.67 71.135 105.72 ;
      RECT MASK 1 71.349 104.67 71.409 105.72 ;
      RECT MASK 1 71.623 104.67 71.683 105.72 ;
      RECT MASK 1 71.897 104.67 71.957 105.72 ;
      RECT MASK 1 72.171 104.67 72.231 105.72 ;
      RECT MASK 1 72.445 104.67 72.505 105.72 ;
      RECT MASK 1 72.719 104.67 72.779 105.72 ;
      RECT MASK 1 72.993 104.67 73.053 105.72 ;
      RECT MASK 1 73.267 104.67 73.327 105.72 ;
      RECT MASK 1 73.541 104.67 73.601 105.72 ;
      RECT MASK 1 73.815 104.67 73.875 105.72 ;
      RECT MASK 1 74.089 104.67 74.149 105.72 ;
      RECT MASK 1 74.363 104.67 74.423 105.72 ;
      RECT MASK 1 74.637 104.67 74.697 105.72 ;
      RECT MASK 1 74.911 104.67 74.971 105.72 ;
      RECT MASK 1 75.185 104.67 75.245 105.72 ;
      RECT MASK 1 75.459 104.67 75.519 105.72 ;
      RECT MASK 1 75.733 104.67 75.793 105.72 ;
      RECT MASK 1 76.007 104.67 76.067 105.72 ;
      RECT MASK 1 76.281 104.67 76.341 105.72 ;
      RECT MASK 1 76.555 104.67 76.615 105.72 ;
      RECT MASK 1 76.829 104.67 76.889 105.72 ;
      RECT MASK 1 77.103 104.67 77.163 105.72 ;
      RECT MASK 1 77.377 104.67 77.437 105.72 ;
      RECT MASK 1 77.651 104.67 77.711 105.72 ;
      RECT MASK 1 77.925 104.67 77.985 105.72 ;
      RECT MASK 1 78.199 104.67 78.259 105.72 ;
      RECT MASK 1 78.473 104.67 78.533 105.72 ;
      RECT MASK 1 78.747 104.67 78.807 105.72 ;
      RECT MASK 1 79.021 104.67 79.081 105.72 ;
      RECT MASK 1 79.295 104.67 79.355 105.72 ;
      RECT MASK 1 79.569 104.67 79.629 105.72 ;
      RECT MASK 1 79.843 104.67 79.903 105.72 ;
      RECT MASK 1 80.117 104.67 80.177 105.72 ;
      RECT MASK 1 80.391 104.67 80.451 105.72 ;
      RECT MASK 1 80.665 104.67 80.725 105.72 ;
      RECT MASK 1 80.939 104.67 80.999 105.72 ;
      RECT MASK 1 81.213 104.67 81.273 105.72 ;
      RECT MASK 1 81.487 104.67 81.547 105.72 ;
      RECT MASK 1 81.761 104.67 81.821 105.72 ;
      RECT MASK 1 82.035 104.67 82.095 105.72 ;
      RECT MASK 1 82.309 104.67 82.369 105.72 ;
      RECT MASK 1 82.583 104.67 82.643 105.72 ;
      RECT MASK 1 82.857 104.67 82.917 105.72 ;
      RECT MASK 1 83.131 104.67 83.191 105.72 ;
      RECT MASK 1 83.405 104.67 83.465 105.72 ;
      RECT MASK 1 83.679 104.67 83.739 105.72 ;
      RECT MASK 1 83.953 104.67 84.013 105.72 ;
      RECT MASK 1 84.227 104.67 84.287 105.72 ;
      RECT MASK 1 84.501 104.67 84.561 105.72 ;
      RECT MASK 1 84.775 104.67 84.835 105.72 ;
      RECT MASK 1 85.049 104.67 85.109 105.72 ;
      RECT MASK 1 85.323 104.67 85.383 105.72 ;
      RECT MASK 1 85.597 104.67 85.657 105.72 ;
      RECT MASK 1 85.871 104.67 85.931 105.72 ;
      RECT MASK 1 86.145 104.67 86.205 105.72 ;
      RECT MASK 1 86.419 104.67 86.479 105.72 ;
      RECT MASK 1 86.693 104.67 86.753 105.72 ;
      RECT MASK 1 86.967 104.67 87.027 105.72 ;
      RECT MASK 1 88.952 104.67 89.012 105.72 ;
      RECT MASK 1 89.226 104.67 89.286 105.72 ;
      RECT MASK 1 89.5 104.67 89.56 105.72 ;
      RECT MASK 1 89.774 104.67 89.834 105.72 ;
      RECT MASK 1 90.048 104.67 90.108 105.72 ;
      RECT MASK 1 90.322 104.67 90.382 105.72 ;
      RECT MASK 1 90.596 104.67 90.656 105.72 ;
      RECT MASK 1 90.87 104.67 90.93 105.72 ;
      RECT MASK 1 91.144 104.67 91.204 105.72 ;
      RECT MASK 1 91.418 104.67 91.478 105.72 ;
      RECT MASK 1 91.692 104.67 91.752 105.72 ;
      RECT MASK 1 91.966 104.67 92.026 105.72 ;
      RECT MASK 1 92.24 104.67 92.3 105.72 ;
      RECT MASK 1 92.514 104.67 92.574 105.72 ;
      RECT MASK 1 92.788 104.67 92.848 105.72 ;
      RECT MASK 1 93.062 104.67 93.122 105.72 ;
      RECT MASK 1 93.336 104.67 93.396 105.72 ;
      RECT MASK 1 93.61 104.67 93.67 105.72 ;
      RECT MASK 1 93.884 104.67 93.944 105.72 ;
      RECT MASK 1 94.158 104.67 94.218 105.72 ;
      RECT MASK 1 94.432 104.67 94.492 105.72 ;
      RECT MASK 1 94.706 104.67 94.766 105.72 ;
      RECT MASK 1 94.98 104.67 95.04 105.72 ;
      RECT MASK 1 95.254 104.67 95.314 105.72 ;
      RECT MASK 1 95.528 104.67 95.588 105.72 ;
      RECT MASK 1 95.802 104.67 95.862 105.72 ;
      RECT MASK 1 96.076 104.67 96.136 105.72 ;
      RECT MASK 1 96.35 104.67 96.41 105.72 ;
      RECT MASK 1 96.624 104.67 96.684 105.72 ;
      RECT MASK 1 96.898 104.67 96.958 105.72 ;
      RECT MASK 1 97.172 104.67 97.232 105.72 ;
      RECT MASK 1 97.446 104.67 97.506 105.72 ;
      RECT MASK 1 97.72 104.67 97.78 105.72 ;
      RECT MASK 1 97.994 104.67 98.054 105.72 ;
      RECT MASK 1 98.268 104.67 98.328 105.72 ;
      RECT MASK 1 98.542 104.67 98.602 105.72 ;
      RECT MASK 1 98.816 104.67 98.876 105.72 ;
      RECT MASK 1 99.09 104.67 99.15 105.72 ;
      RECT MASK 1 99.364 104.67 99.424 105.72 ;
      RECT MASK 1 99.638 104.67 99.698 105.72 ;
      RECT MASK 1 99.912 104.67 99.972 105.72 ;
      RECT MASK 1 100.186 104.67 100.246 105.72 ;
      RECT MASK 1 100.46 104.67 100.52 105.72 ;
      RECT MASK 1 100.734 104.67 100.794 105.72 ;
      RECT MASK 1 101.008 104.67 101.068 105.72 ;
      RECT MASK 1 101.282 104.67 101.342 105.72 ;
      RECT MASK 1 101.556 104.67 101.616 105.72 ;
      RECT MASK 1 101.83 104.67 101.89 105.72 ;
      RECT MASK 1 102.104 104.67 102.164 105.72 ;
      RECT MASK 1 102.378 104.67 102.438 105.72 ;
      RECT MASK 1 102.652 104.67 102.712 105.72 ;
      RECT MASK 1 102.926 104.67 102.986 105.72 ;
      RECT MASK 1 103.2 104.67 103.26 105.72 ;
      RECT MASK 1 103.474 104.67 103.534 105.72 ;
      RECT MASK 1 103.748 104.67 103.808 105.72 ;
      RECT MASK 1 104.022 104.67 104.082 105.72 ;
      RECT MASK 1 104.296 104.67 104.356 105.72 ;
      RECT MASK 1 104.57 104.67 104.63 105.72 ;
      RECT MASK 1 104.844 104.67 104.904 105.72 ;
      RECT MASK 1 105.118 104.67 105.178 105.72 ;
      RECT MASK 1 105.392 104.67 105.452 105.72 ;
      RECT MASK 1 105.666 104.67 105.726 105.72 ;
      RECT MASK 1 105.94 104.67 106 105.72 ;
      RECT MASK 1 106.214 104.67 106.274 105.72 ;
      RECT MASK 1 106.488 104.67 106.548 105.72 ;
      RECT MASK 1 106.762 104.67 106.822 105.72 ;
      RECT MASK 1 107.036 104.67 107.096 105.72 ;
      RECT MASK 1 107.31 104.67 107.37 105.72 ;
      RECT MASK 1 107.584 104.67 107.644 105.72 ;
      RECT MASK 1 107.858 104.67 107.918 105.72 ;
      RECT MASK 1 108.132 104.67 108.192 105.72 ;
      RECT MASK 1 108.406 104.67 108.466 105.72 ;
      RECT MASK 1 108.68 104.67 108.74 105.72 ;
      RECT MASK 1 108.954 104.67 109.014 105.72 ;
      RECT MASK 1 109.228 104.67 109.288 105.72 ;
      RECT MASK 1 109.502 104.67 109.562 105.72 ;
      RECT MASK 1 109.776 104.67 109.836 105.72 ;
      RECT MASK 1 110.05 104.67 110.11 105.72 ;
      RECT MASK 1 110.324 104.67 110.384 105.72 ;
      RECT MASK 1 110.598 104.67 110.658 105.72 ;
      RECT MASK 1 110.872 104.67 110.932 105.72 ;
      RECT MASK 1 111.146 104.67 111.206 105.72 ;
      RECT MASK 1 111.42 104.67 111.48 105.72 ;
      RECT MASK 1 111.694 104.67 111.754 105.72 ;
      RECT MASK 1 111.968 104.67 112.028 105.72 ;
      RECT MASK 1 112.242 104.67 112.302 105.72 ;
      RECT MASK 1 112.516 104.67 112.576 105.72 ;
      RECT MASK 1 112.79 104.67 112.85 105.72 ;
      RECT MASK 1 113.064 104.67 113.124 105.72 ;
      RECT MASK 1 113.338 104.67 113.398 105.72 ;
      RECT MASK 1 113.612 104.67 113.672 105.72 ;
      RECT MASK 1 113.886 104.67 113.946 105.72 ;
      RECT MASK 1 114.16 104.67 114.22 105.72 ;
      RECT MASK 1 114.434 104.67 114.494 105.72 ;
      RECT MASK 1 114.708 104.67 114.768 105.72 ;
      RECT MASK 1 114.982 104.67 115.042 105.72 ;
      RECT MASK 1 115.256 104.67 115.316 105.72 ;
      RECT MASK 1 115.53 104.67 115.59 105.72 ;
      RECT MASK 1 115.804 104.67 115.864 105.72 ;
      RECT MASK 1 116.078 104.67 116.138 105.72 ;
      RECT MASK 1 116.352 104.67 116.412 105.72 ;
      RECT MASK 1 116.626 104.67 116.686 105.72 ;
      RECT MASK 1 116.9 104.67 116.96 105.72 ;
      RECT MASK 1 117.174 104.67 117.234 105.72 ;
      RECT MASK 1 117.448 104.67 117.508 105.72 ;
      RECT MASK 1 117.722 104.67 117.782 105.72 ;
      RECT MASK 1 117.996 104.67 118.056 105.72 ;
      RECT MASK 1 118.27 104.67 118.33 105.72 ;
      RECT MASK 1 118.544 104.67 118.604 105.72 ;
      RECT MASK 1 118.818 104.67 118.878 105.72 ;
      RECT MASK 1 119.092 104.67 119.152 105.72 ;
      RECT MASK 1 119.366 104.67 119.426 105.72 ;
      RECT MASK 1 119.64 104.67 119.7 105.72 ;
      RECT MASK 1 119.914 104.67 119.974 105.72 ;
      RECT MASK 1 120.188 104.67 120.248 105.72 ;
      RECT MASK 1 120.462 104.67 120.522 105.72 ;
      RECT MASK 1 120.736 104.67 120.796 105.72 ;
      RECT MASK 1 121.01 104.67 121.07 105.72 ;
      RECT MASK 1 121.284 104.67 121.344 105.72 ;
      RECT MASK 1 121.558 104.67 121.618 105.72 ;
      RECT MASK 1 121.832 104.67 121.892 105.72 ;
      RECT MASK 1 122.106 104.67 122.166 105.72 ;
      RECT MASK 1 122.38 104.67 122.44 105.72 ;
      RECT MASK 1 122.654 104.67 122.714 105.72 ;
      RECT MASK 1 122.928 104.67 122.988 105.72 ;
      RECT MASK 1 123.202 104.67 123.262 105.72 ;
      RECT MASK 1 123.476 104.67 123.536 105.72 ;
      RECT MASK 1 123.75 104.67 123.81 105.72 ;
      RECT MASK 1 124.024 104.67 124.084 105.72 ;
      RECT MASK 1 124.298 104.67 124.358 105.72 ;
      RECT MASK 1 124.572 104.67 124.632 105.72 ;
      RECT MASK 1 124.846 104.67 124.906 105.72 ;
      RECT MASK 1 125.12 104.67 125.18 105.72 ;
      RECT MASK 1 125.394 104.67 125.454 105.72 ;
      RECT MASK 1 125.668 104.67 125.728 105.72 ;
      RECT MASK 1 125.942 104.67 126.002 105.72 ;
      RECT MASK 1 126.216 104.67 126.276 105.72 ;
      RECT MASK 1 126.49 104.67 126.55 105.72 ;
      RECT MASK 1 126.764 104.67 126.824 105.72 ;
      RECT MASK 1 127.038 104.67 127.098 105.72 ;
      RECT MASK 1 127.312 104.67 127.372 105.72 ;
      RECT MASK 1 127.586 104.67 127.646 105.72 ;
      RECT MASK 1 2.201 106.38 2.261 107.43 ;
      RECT MASK 1 2.475 106.38 2.535 107.43 ;
      RECT MASK 1 2.749 106.38 2.809 107.43 ;
      RECT MASK 1 3.023 106.38 3.083 107.43 ;
      RECT MASK 1 3.297 106.38 3.357 107.43 ;
      RECT MASK 1 3.571 106.38 3.631 107.43 ;
      RECT MASK 1 3.845 106.38 3.905 107.43 ;
      RECT MASK 1 4.119 106.38 4.179 107.43 ;
      RECT MASK 1 4.393 106.38 4.453 107.43 ;
      RECT MASK 1 4.667 106.38 4.727 107.43 ;
      RECT MASK 1 4.941 106.38 5.001 107.43 ;
      RECT MASK 1 5.215 106.38 5.275 107.43 ;
      RECT MASK 1 5.489 106.38 5.549 107.43 ;
      RECT MASK 1 5.763 106.38 5.823 107.43 ;
      RECT MASK 1 6.037 106.38 6.097 107.43 ;
      RECT MASK 1 6.311 106.38 6.371 107.43 ;
      RECT MASK 1 6.585 106.38 6.645 107.43 ;
      RECT MASK 1 6.859 106.38 6.919 107.43 ;
      RECT MASK 1 7.133 106.38 7.193 107.43 ;
      RECT MASK 1 7.407 106.38 7.467 107.43 ;
      RECT MASK 1 7.681 106.38 7.741 107.43 ;
      RECT MASK 1 7.955 106.38 8.015 107.43 ;
      RECT MASK 1 8.229 106.38 8.289 107.43 ;
      RECT MASK 1 8.503 106.38 8.563 107.43 ;
      RECT MASK 1 8.777 106.38 8.837 107.43 ;
      RECT MASK 1 9.051 106.38 9.111 107.43 ;
      RECT MASK 1 9.325 106.38 9.385 107.43 ;
      RECT MASK 1 9.599 106.38 9.659 107.43 ;
      RECT MASK 1 9.873 106.38 9.933 107.43 ;
      RECT MASK 1 10.147 106.38 10.207 107.43 ;
      RECT MASK 1 10.421 106.38 10.481 107.43 ;
      RECT MASK 1 10.695 106.38 10.755 107.43 ;
      RECT MASK 1 10.969 106.38 11.029 107.43 ;
      RECT MASK 1 11.243 106.38 11.303 107.43 ;
      RECT MASK 1 11.517 106.38 11.577 107.43 ;
      RECT MASK 1 11.791 106.38 11.851 107.43 ;
      RECT MASK 1 12.065 106.38 12.125 107.43 ;
      RECT MASK 1 12.339 106.38 12.399 107.43 ;
      RECT MASK 1 12.613 106.38 12.673 107.43 ;
      RECT MASK 1 12.887 106.38 12.947 107.43 ;
      RECT MASK 1 13.161 106.38 13.221 107.43 ;
      RECT MASK 1 13.435 106.38 13.495 107.43 ;
      RECT MASK 1 13.709 106.38 13.769 107.43 ;
      RECT MASK 1 13.983 106.38 14.043 107.43 ;
      RECT MASK 1 14.257 106.38 14.317 107.43 ;
      RECT MASK 1 14.531 106.38 14.591 107.43 ;
      RECT MASK 1 14.805 106.38 14.865 107.43 ;
      RECT MASK 1 15.079 106.38 15.139 107.43 ;
      RECT MASK 1 15.353 106.38 15.413 107.43 ;
      RECT MASK 1 15.627 106.38 15.687 107.43 ;
      RECT MASK 1 15.901 106.38 15.961 107.43 ;
      RECT MASK 1 16.175 106.38 16.235 107.43 ;
      RECT MASK 1 16.449 106.38 16.509 107.43 ;
      RECT MASK 1 16.723 106.38 16.783 107.43 ;
      RECT MASK 1 16.997 106.38 17.057 107.43 ;
      RECT MASK 1 17.271 106.38 17.331 107.43 ;
      RECT MASK 1 17.545 106.38 17.605 107.43 ;
      RECT MASK 1 17.819 106.38 17.879 107.43 ;
      RECT MASK 1 18.093 106.38 18.153 107.43 ;
      RECT MASK 1 18.367 106.38 18.427 107.43 ;
      RECT MASK 1 18.641 106.38 18.701 107.43 ;
      RECT MASK 1 18.915 106.38 18.975 107.43 ;
      RECT MASK 1 19.189 106.38 19.249 107.43 ;
      RECT MASK 1 19.463 106.38 19.523 107.43 ;
      RECT MASK 1 19.737 106.38 19.797 107.43 ;
      RECT MASK 1 20.011 106.38 20.071 107.43 ;
      RECT MASK 1 20.285 106.38 20.345 107.43 ;
      RECT MASK 1 20.559 106.38 20.619 107.43 ;
      RECT MASK 1 20.833 106.38 20.893 107.43 ;
      RECT MASK 1 21.107 106.38 21.167 107.43 ;
      RECT MASK 1 21.381 106.38 21.441 107.43 ;
      RECT MASK 1 21.655 106.38 21.715 107.43 ;
      RECT MASK 1 21.929 106.38 21.989 107.43 ;
      RECT MASK 1 22.203 106.38 22.263 107.43 ;
      RECT MASK 1 22.477 106.38 22.537 107.43 ;
      RECT MASK 1 22.751 106.38 22.811 107.43 ;
      RECT MASK 1 23.025 106.38 23.085 107.43 ;
      RECT MASK 1 23.299 106.38 23.359 107.43 ;
      RECT MASK 1 23.573 106.38 23.633 107.43 ;
      RECT MASK 1 23.847 106.38 23.907 107.43 ;
      RECT MASK 1 24.121 106.38 24.181 107.43 ;
      RECT MASK 1 24.395 106.38 24.455 107.43 ;
      RECT MASK 1 24.669 106.38 24.729 107.43 ;
      RECT MASK 1 24.943 106.38 25.003 107.43 ;
      RECT MASK 1 25.217 106.38 25.277 107.43 ;
      RECT MASK 1 25.491 106.38 25.551 107.43 ;
      RECT MASK 1 25.765 106.38 25.825 107.43 ;
      RECT MASK 1 26.039 106.38 26.099 107.43 ;
      RECT MASK 1 26.313 106.38 26.373 107.43 ;
      RECT MASK 1 26.587 106.38 26.647 107.43 ;
      RECT MASK 1 26.861 106.38 26.921 107.43 ;
      RECT MASK 1 27.135 106.38 27.195 107.43 ;
      RECT MASK 1 27.409 106.38 27.469 107.43 ;
      RECT MASK 1 27.683 106.38 27.743 107.43 ;
      RECT MASK 1 27.957 106.38 28.017 107.43 ;
      RECT MASK 1 28.231 106.38 28.291 107.43 ;
      RECT MASK 1 28.505 106.38 28.565 107.43 ;
      RECT MASK 1 28.779 106.38 28.839 107.43 ;
      RECT MASK 1 29.053 106.38 29.113 107.43 ;
      RECT MASK 1 29.327 106.38 29.387 107.43 ;
      RECT MASK 1 29.601 106.38 29.661 107.43 ;
      RECT MASK 1 29.875 106.38 29.935 107.43 ;
      RECT MASK 1 30.149 106.38 30.209 107.43 ;
      RECT MASK 1 30.423 106.38 30.483 107.43 ;
      RECT MASK 1 30.697 106.38 30.757 107.43 ;
      RECT MASK 1 30.971 106.38 31.031 107.43 ;
      RECT MASK 1 31.245 106.38 31.305 107.43 ;
      RECT MASK 1 31.519 106.38 31.579 107.43 ;
      RECT MASK 1 31.793 106.38 31.853 107.43 ;
      RECT MASK 1 32.067 106.38 32.127 107.43 ;
      RECT MASK 1 32.341 106.38 32.401 107.43 ;
      RECT MASK 1 32.615 106.38 32.675 107.43 ;
      RECT MASK 1 32.889 106.38 32.949 107.43 ;
      RECT MASK 1 33.163 106.38 33.223 107.43 ;
      RECT MASK 1 33.437 106.38 33.497 107.43 ;
      RECT MASK 1 33.711 106.38 33.771 107.43 ;
      RECT MASK 1 33.985 106.38 34.045 107.43 ;
      RECT MASK 1 34.259 106.38 34.319 107.43 ;
      RECT MASK 1 34.533 106.38 34.593 107.43 ;
      RECT MASK 1 34.807 106.38 34.867 107.43 ;
      RECT MASK 1 35.081 106.38 35.141 107.43 ;
      RECT MASK 1 35.355 106.38 35.415 107.43 ;
      RECT MASK 1 35.629 106.38 35.689 107.43 ;
      RECT MASK 1 35.903 106.38 35.963 107.43 ;
      RECT MASK 1 36.177 106.38 36.237 107.43 ;
      RECT MASK 1 36.451 106.38 36.511 107.43 ;
      RECT MASK 1 36.725 106.38 36.785 107.43 ;
      RECT MASK 1 36.999 106.38 37.059 107.43 ;
      RECT MASK 1 37.273 106.38 37.333 107.43 ;
      RECT MASK 1 37.547 106.38 37.607 107.43 ;
      RECT MASK 1 37.821 106.38 37.881 107.43 ;
      RECT MASK 1 38.095 106.38 38.155 107.43 ;
      RECT MASK 1 38.369 106.38 38.429 107.43 ;
      RECT MASK 1 38.643 106.38 38.703 107.43 ;
      RECT MASK 1 38.917 106.38 38.977 107.43 ;
      RECT MASK 1 39.191 106.38 39.251 107.43 ;
      RECT MASK 1 39.465 106.38 39.525 107.43 ;
      RECT MASK 1 39.739 106.38 39.799 107.43 ;
      RECT MASK 1 40.013 106.38 40.073 107.43 ;
      RECT MASK 1 40.287 106.38 40.347 107.43 ;
      RECT MASK 1 40.561 106.38 40.621 107.43 ;
      RECT MASK 1 40.835 106.38 40.895 107.43 ;
      RECT MASK 1 41.109 106.38 41.169 107.43 ;
      RECT MASK 1 41.383 106.38 41.443 107.43 ;
      RECT MASK 1 41.657 106.38 41.717 107.43 ;
      RECT MASK 1 41.931 106.38 41.991 107.43 ;
      RECT MASK 1 42.205 106.38 42.265 107.43 ;
      RECT MASK 1 42.479 106.38 42.539 107.43 ;
      RECT MASK 1 42.753 106.38 42.813 107.43 ;
      RECT MASK 1 43.027 106.38 43.087 107.43 ;
      RECT MASK 1 43.301 106.38 43.361 107.43 ;
      RECT MASK 1 43.575 106.38 43.635 107.43 ;
      RECT MASK 1 45.593 106.38 45.653 107.43 ;
      RECT MASK 1 45.867 106.38 45.927 107.43 ;
      RECT MASK 1 46.141 106.38 46.201 107.43 ;
      RECT MASK 1 46.415 106.38 46.475 107.43 ;
      RECT MASK 1 46.689 106.38 46.749 107.43 ;
      RECT MASK 1 46.963 106.38 47.023 107.43 ;
      RECT MASK 1 47.237 106.38 47.297 107.43 ;
      RECT MASK 1 47.511 106.38 47.571 107.43 ;
      RECT MASK 1 47.785 106.38 47.845 107.43 ;
      RECT MASK 1 48.059 106.38 48.119 107.43 ;
      RECT MASK 1 48.333 106.38 48.393 107.43 ;
      RECT MASK 1 48.607 106.38 48.667 107.43 ;
      RECT MASK 1 48.881 106.38 48.941 107.43 ;
      RECT MASK 1 49.155 106.38 49.215 107.43 ;
      RECT MASK 1 49.429 106.38 49.489 107.43 ;
      RECT MASK 1 49.703 106.38 49.763 107.43 ;
      RECT MASK 1 49.977 106.38 50.037 107.43 ;
      RECT MASK 1 50.251 106.38 50.311 107.43 ;
      RECT MASK 1 50.525 106.38 50.585 107.43 ;
      RECT MASK 1 50.799 106.38 50.859 107.43 ;
      RECT MASK 1 51.073 106.38 51.133 107.43 ;
      RECT MASK 1 51.347 106.38 51.407 107.43 ;
      RECT MASK 1 51.621 106.38 51.681 107.43 ;
      RECT MASK 1 51.895 106.38 51.955 107.43 ;
      RECT MASK 1 52.169 106.38 52.229 107.43 ;
      RECT MASK 1 52.443 106.38 52.503 107.43 ;
      RECT MASK 1 52.717 106.38 52.777 107.43 ;
      RECT MASK 1 52.991 106.38 53.051 107.43 ;
      RECT MASK 1 53.265 106.38 53.325 107.43 ;
      RECT MASK 1 53.539 106.38 53.599 107.43 ;
      RECT MASK 1 53.813 106.38 53.873 107.43 ;
      RECT MASK 1 54.087 106.38 54.147 107.43 ;
      RECT MASK 1 54.361 106.38 54.421 107.43 ;
      RECT MASK 1 54.635 106.38 54.695 107.43 ;
      RECT MASK 1 54.909 106.38 54.969 107.43 ;
      RECT MASK 1 55.183 106.38 55.243 107.43 ;
      RECT MASK 1 55.457 106.38 55.517 107.43 ;
      RECT MASK 1 55.731 106.38 55.791 107.43 ;
      RECT MASK 1 56.005 106.38 56.065 107.43 ;
      RECT MASK 1 56.279 106.38 56.339 107.43 ;
      RECT MASK 1 56.553 106.38 56.613 107.43 ;
      RECT MASK 1 56.827 106.38 56.887 107.43 ;
      RECT MASK 1 57.101 106.38 57.161 107.43 ;
      RECT MASK 1 57.375 106.38 57.435 107.43 ;
      RECT MASK 1 57.649 106.38 57.709 107.43 ;
      RECT MASK 1 57.923 106.38 57.983 107.43 ;
      RECT MASK 1 58.197 106.38 58.257 107.43 ;
      RECT MASK 1 58.471 106.38 58.531 107.43 ;
      RECT MASK 1 58.745 106.38 58.805 107.43 ;
      RECT MASK 1 59.019 106.38 59.079 107.43 ;
      RECT MASK 1 59.293 106.38 59.353 107.43 ;
      RECT MASK 1 59.567 106.38 59.627 107.43 ;
      RECT MASK 1 59.841 106.38 59.901 107.43 ;
      RECT MASK 1 60.115 106.38 60.175 107.43 ;
      RECT MASK 1 60.389 106.38 60.449 107.43 ;
      RECT MASK 1 60.663 106.38 60.723 107.43 ;
      RECT MASK 1 60.937 106.38 60.997 107.43 ;
      RECT MASK 1 61.211 106.38 61.271 107.43 ;
      RECT MASK 1 61.485 106.38 61.545 107.43 ;
      RECT MASK 1 61.759 106.38 61.819 107.43 ;
      RECT MASK 1 62.033 106.38 62.093 107.43 ;
      RECT MASK 1 62.307 106.38 62.367 107.43 ;
      RECT MASK 1 62.581 106.38 62.641 107.43 ;
      RECT MASK 1 62.855 106.38 62.915 107.43 ;
      RECT MASK 1 63.129 106.38 63.189 107.43 ;
      RECT MASK 1 63.403 106.38 63.463 107.43 ;
      RECT MASK 1 63.677 106.38 63.737 107.43 ;
      RECT MASK 1 63.951 106.38 64.011 107.43 ;
      RECT MASK 1 64.225 106.38 64.285 107.43 ;
      RECT MASK 1 64.499 106.38 64.559 107.43 ;
      RECT MASK 1 64.773 106.38 64.833 107.43 ;
      RECT MASK 1 65.047 106.38 65.107 107.43 ;
      RECT MASK 1 65.321 106.38 65.381 107.43 ;
      RECT MASK 1 65.595 106.38 65.655 107.43 ;
      RECT MASK 1 65.869 106.38 65.929 107.43 ;
      RECT MASK 1 66.143 106.38 66.203 107.43 ;
      RECT MASK 1 66.417 106.38 66.477 107.43 ;
      RECT MASK 1 66.691 106.38 66.751 107.43 ;
      RECT MASK 1 66.965 106.38 67.025 107.43 ;
      RECT MASK 1 67.239 106.38 67.299 107.43 ;
      RECT MASK 1 67.513 106.38 67.573 107.43 ;
      RECT MASK 1 67.787 106.38 67.847 107.43 ;
      RECT MASK 1 68.061 106.38 68.121 107.43 ;
      RECT MASK 1 68.335 106.38 68.395 107.43 ;
      RECT MASK 1 68.609 106.38 68.669 107.43 ;
      RECT MASK 1 68.883 106.38 68.943 107.43 ;
      RECT MASK 1 69.157 106.38 69.217 107.43 ;
      RECT MASK 1 69.431 106.38 69.491 107.43 ;
      RECT MASK 1 69.705 106.38 69.765 107.43 ;
      RECT MASK 1 69.979 106.38 70.039 107.43 ;
      RECT MASK 1 70.253 106.38 70.313 107.43 ;
      RECT MASK 1 70.527 106.38 70.587 107.43 ;
      RECT MASK 1 70.801 106.38 70.861 107.43 ;
      RECT MASK 1 71.075 106.38 71.135 107.43 ;
      RECT MASK 1 71.349 106.38 71.409 107.43 ;
      RECT MASK 1 71.623 106.38 71.683 107.43 ;
      RECT MASK 1 71.897 106.38 71.957 107.43 ;
      RECT MASK 1 72.171 106.38 72.231 107.43 ;
      RECT MASK 1 72.445 106.38 72.505 107.43 ;
      RECT MASK 1 72.719 106.38 72.779 107.43 ;
      RECT MASK 1 72.993 106.38 73.053 107.43 ;
      RECT MASK 1 73.267 106.38 73.327 107.43 ;
      RECT MASK 1 73.541 106.38 73.601 107.43 ;
      RECT MASK 1 73.815 106.38 73.875 107.43 ;
      RECT MASK 1 74.089 106.38 74.149 107.43 ;
      RECT MASK 1 74.363 106.38 74.423 107.43 ;
      RECT MASK 1 74.637 106.38 74.697 107.43 ;
      RECT MASK 1 74.911 106.38 74.971 107.43 ;
      RECT MASK 1 75.185 106.38 75.245 107.43 ;
      RECT MASK 1 75.459 106.38 75.519 107.43 ;
      RECT MASK 1 75.733 106.38 75.793 107.43 ;
      RECT MASK 1 76.007 106.38 76.067 107.43 ;
      RECT MASK 1 76.281 106.38 76.341 107.43 ;
      RECT MASK 1 76.555 106.38 76.615 107.43 ;
      RECT MASK 1 76.829 106.38 76.889 107.43 ;
      RECT MASK 1 77.103 106.38 77.163 107.43 ;
      RECT MASK 1 77.377 106.38 77.437 107.43 ;
      RECT MASK 1 77.651 106.38 77.711 107.43 ;
      RECT MASK 1 77.925 106.38 77.985 107.43 ;
      RECT MASK 1 78.199 106.38 78.259 107.43 ;
      RECT MASK 1 78.473 106.38 78.533 107.43 ;
      RECT MASK 1 78.747 106.38 78.807 107.43 ;
      RECT MASK 1 79.021 106.38 79.081 107.43 ;
      RECT MASK 1 79.295 106.38 79.355 107.43 ;
      RECT MASK 1 79.569 106.38 79.629 107.43 ;
      RECT MASK 1 79.843 106.38 79.903 107.43 ;
      RECT MASK 1 80.117 106.38 80.177 107.43 ;
      RECT MASK 1 80.391 106.38 80.451 107.43 ;
      RECT MASK 1 80.665 106.38 80.725 107.43 ;
      RECT MASK 1 80.939 106.38 80.999 107.43 ;
      RECT MASK 1 81.213 106.38 81.273 107.43 ;
      RECT MASK 1 81.487 106.38 81.547 107.43 ;
      RECT MASK 1 81.761 106.38 81.821 107.43 ;
      RECT MASK 1 82.035 106.38 82.095 107.43 ;
      RECT MASK 1 82.309 106.38 82.369 107.43 ;
      RECT MASK 1 82.583 106.38 82.643 107.43 ;
      RECT MASK 1 82.857 106.38 82.917 107.43 ;
      RECT MASK 1 83.131 106.38 83.191 107.43 ;
      RECT MASK 1 83.405 106.38 83.465 107.43 ;
      RECT MASK 1 83.679 106.38 83.739 107.43 ;
      RECT MASK 1 83.953 106.38 84.013 107.43 ;
      RECT MASK 1 84.227 106.38 84.287 107.43 ;
      RECT MASK 1 84.501 106.38 84.561 107.43 ;
      RECT MASK 1 84.775 106.38 84.835 107.43 ;
      RECT MASK 1 85.049 106.38 85.109 107.43 ;
      RECT MASK 1 85.323 106.38 85.383 107.43 ;
      RECT MASK 1 85.597 106.38 85.657 107.43 ;
      RECT MASK 1 85.871 106.38 85.931 107.43 ;
      RECT MASK 1 86.145 106.38 86.205 107.43 ;
      RECT MASK 1 86.419 106.38 86.479 107.43 ;
      RECT MASK 1 86.693 106.38 86.753 107.43 ;
      RECT MASK 1 86.967 106.38 87.027 107.43 ;
      RECT MASK 1 88.952 106.38 89.012 107.43 ;
      RECT MASK 1 89.226 106.38 89.286 107.43 ;
      RECT MASK 1 89.5 106.38 89.56 107.43 ;
      RECT MASK 1 89.774 106.38 89.834 107.43 ;
      RECT MASK 1 90.048 106.38 90.108 107.43 ;
      RECT MASK 1 90.322 106.38 90.382 107.43 ;
      RECT MASK 1 90.596 106.38 90.656 107.43 ;
      RECT MASK 1 90.87 106.38 90.93 107.43 ;
      RECT MASK 1 91.144 106.38 91.204 107.43 ;
      RECT MASK 1 91.418 106.38 91.478 107.43 ;
      RECT MASK 1 91.692 106.38 91.752 107.43 ;
      RECT MASK 1 91.966 106.38 92.026 107.43 ;
      RECT MASK 1 92.24 106.38 92.3 107.43 ;
      RECT MASK 1 92.514 106.38 92.574 107.43 ;
      RECT MASK 1 92.788 106.38 92.848 107.43 ;
      RECT MASK 1 93.062 106.38 93.122 107.43 ;
      RECT MASK 1 93.336 106.38 93.396 107.43 ;
      RECT MASK 1 93.61 106.38 93.67 107.43 ;
      RECT MASK 1 93.884 106.38 93.944 107.43 ;
      RECT MASK 1 94.158 106.38 94.218 107.43 ;
      RECT MASK 1 94.432 106.38 94.492 107.43 ;
      RECT MASK 1 94.706 106.38 94.766 107.43 ;
      RECT MASK 1 94.98 106.38 95.04 107.43 ;
      RECT MASK 1 95.254 106.38 95.314 107.43 ;
      RECT MASK 1 95.528 106.38 95.588 107.43 ;
      RECT MASK 1 95.802 106.38 95.862 107.43 ;
      RECT MASK 1 96.076 106.38 96.136 107.43 ;
      RECT MASK 1 96.35 106.38 96.41 107.43 ;
      RECT MASK 1 96.624 106.38 96.684 107.43 ;
      RECT MASK 1 96.898 106.38 96.958 107.43 ;
      RECT MASK 1 97.172 106.38 97.232 107.43 ;
      RECT MASK 1 97.446 106.38 97.506 107.43 ;
      RECT MASK 1 97.72 106.38 97.78 107.43 ;
      RECT MASK 1 97.994 106.38 98.054 107.43 ;
      RECT MASK 1 98.268 106.38 98.328 107.43 ;
      RECT MASK 1 98.542 106.38 98.602 107.43 ;
      RECT MASK 1 98.816 106.38 98.876 107.43 ;
      RECT MASK 1 99.09 106.38 99.15 107.43 ;
      RECT MASK 1 99.364 106.38 99.424 107.43 ;
      RECT MASK 1 99.638 106.38 99.698 107.43 ;
      RECT MASK 1 99.912 106.38 99.972 107.43 ;
      RECT MASK 1 100.186 106.38 100.246 107.43 ;
      RECT MASK 1 100.46 106.38 100.52 107.43 ;
      RECT MASK 1 100.734 106.38 100.794 107.43 ;
      RECT MASK 1 101.008 106.38 101.068 107.43 ;
      RECT MASK 1 101.282 106.38 101.342 107.43 ;
      RECT MASK 1 101.556 106.38 101.616 107.43 ;
      RECT MASK 1 101.83 106.38 101.89 107.43 ;
      RECT MASK 1 102.104 106.38 102.164 107.43 ;
      RECT MASK 1 102.378 106.38 102.438 107.43 ;
      RECT MASK 1 102.652 106.38 102.712 107.43 ;
      RECT MASK 1 102.926 106.38 102.986 107.43 ;
      RECT MASK 1 103.2 106.38 103.26 107.43 ;
      RECT MASK 1 103.474 106.38 103.534 107.43 ;
      RECT MASK 1 103.748 106.38 103.808 107.43 ;
      RECT MASK 1 104.022 106.38 104.082 107.43 ;
      RECT MASK 1 104.296 106.38 104.356 107.43 ;
      RECT MASK 1 104.57 106.38 104.63 107.43 ;
      RECT MASK 1 104.844 106.38 104.904 107.43 ;
      RECT MASK 1 105.118 106.38 105.178 107.43 ;
      RECT MASK 1 105.392 106.38 105.452 107.43 ;
      RECT MASK 1 105.666 106.38 105.726 107.43 ;
      RECT MASK 1 105.94 106.38 106 107.43 ;
      RECT MASK 1 106.214 106.38 106.274 107.43 ;
      RECT MASK 1 106.488 106.38 106.548 107.43 ;
      RECT MASK 1 106.762 106.38 106.822 107.43 ;
      RECT MASK 1 107.036 106.38 107.096 107.43 ;
      RECT MASK 1 107.31 106.38 107.37 107.43 ;
      RECT MASK 1 107.584 106.38 107.644 107.43 ;
      RECT MASK 1 107.858 106.38 107.918 107.43 ;
      RECT MASK 1 108.132 106.38 108.192 107.43 ;
      RECT MASK 1 108.406 106.38 108.466 107.43 ;
      RECT MASK 1 108.68 106.38 108.74 107.43 ;
      RECT MASK 1 108.954 106.38 109.014 107.43 ;
      RECT MASK 1 109.228 106.38 109.288 107.43 ;
      RECT MASK 1 109.502 106.38 109.562 107.43 ;
      RECT MASK 1 109.776 106.38 109.836 107.43 ;
      RECT MASK 1 110.05 106.38 110.11 107.43 ;
      RECT MASK 1 110.324 106.38 110.384 107.43 ;
      RECT MASK 1 110.598 106.38 110.658 107.43 ;
      RECT MASK 1 110.872 106.38 110.932 107.43 ;
      RECT MASK 1 111.146 106.38 111.206 107.43 ;
      RECT MASK 1 111.42 106.38 111.48 107.43 ;
      RECT MASK 1 111.694 106.38 111.754 107.43 ;
      RECT MASK 1 111.968 106.38 112.028 107.43 ;
      RECT MASK 1 112.242 106.38 112.302 107.43 ;
      RECT MASK 1 112.516 106.38 112.576 107.43 ;
      RECT MASK 1 112.79 106.38 112.85 107.43 ;
      RECT MASK 1 113.064 106.38 113.124 107.43 ;
      RECT MASK 1 113.338 106.38 113.398 107.43 ;
      RECT MASK 1 113.612 106.38 113.672 107.43 ;
      RECT MASK 1 113.886 106.38 113.946 107.43 ;
      RECT MASK 1 114.16 106.38 114.22 107.43 ;
      RECT MASK 1 114.434 106.38 114.494 107.43 ;
      RECT MASK 1 114.708 106.38 114.768 107.43 ;
      RECT MASK 1 114.982 106.38 115.042 107.43 ;
      RECT MASK 1 115.256 106.38 115.316 107.43 ;
      RECT MASK 1 115.53 106.38 115.59 107.43 ;
      RECT MASK 1 115.804 106.38 115.864 107.43 ;
      RECT MASK 1 116.078 106.38 116.138 107.43 ;
      RECT MASK 1 116.352 106.38 116.412 107.43 ;
      RECT MASK 1 116.626 106.38 116.686 107.43 ;
      RECT MASK 1 116.9 106.38 116.96 107.43 ;
      RECT MASK 1 117.174 106.38 117.234 107.43 ;
      RECT MASK 1 117.448 106.38 117.508 107.43 ;
      RECT MASK 1 117.722 106.38 117.782 107.43 ;
      RECT MASK 1 117.996 106.38 118.056 107.43 ;
      RECT MASK 1 118.27 106.38 118.33 107.43 ;
      RECT MASK 1 118.544 106.38 118.604 107.43 ;
      RECT MASK 1 118.818 106.38 118.878 107.43 ;
      RECT MASK 1 119.092 106.38 119.152 107.43 ;
      RECT MASK 1 119.366 106.38 119.426 107.43 ;
      RECT MASK 1 119.64 106.38 119.7 107.43 ;
      RECT MASK 1 119.914 106.38 119.974 107.43 ;
      RECT MASK 1 120.188 106.38 120.248 107.43 ;
      RECT MASK 1 120.462 106.38 120.522 107.43 ;
      RECT MASK 1 120.736 106.38 120.796 107.43 ;
      RECT MASK 1 121.01 106.38 121.07 107.43 ;
      RECT MASK 1 121.284 106.38 121.344 107.43 ;
      RECT MASK 1 121.558 106.38 121.618 107.43 ;
      RECT MASK 1 121.832 106.38 121.892 107.43 ;
      RECT MASK 1 122.106 106.38 122.166 107.43 ;
      RECT MASK 1 122.38 106.38 122.44 107.43 ;
      RECT MASK 1 122.654 106.38 122.714 107.43 ;
      RECT MASK 1 122.928 106.38 122.988 107.43 ;
      RECT MASK 1 123.202 106.38 123.262 107.43 ;
      RECT MASK 1 123.476 106.38 123.536 107.43 ;
      RECT MASK 1 123.75 106.38 123.81 107.43 ;
      RECT MASK 1 124.024 106.38 124.084 107.43 ;
      RECT MASK 1 124.298 106.38 124.358 107.43 ;
      RECT MASK 1 124.572 106.38 124.632 107.43 ;
      RECT MASK 1 124.846 106.38 124.906 107.43 ;
      RECT MASK 1 125.12 106.38 125.18 107.43 ;
      RECT MASK 1 125.394 106.38 125.454 107.43 ;
      RECT MASK 1 125.668 106.38 125.728 107.43 ;
      RECT MASK 1 125.942 106.38 126.002 107.43 ;
      RECT MASK 1 126.216 106.38 126.276 107.43 ;
      RECT MASK 1 126.49 106.38 126.55 107.43 ;
      RECT MASK 1 126.764 106.38 126.824 107.43 ;
      RECT MASK 1 127.038 106.38 127.098 107.43 ;
      RECT MASK 1 127.312 106.38 127.372 107.43 ;
      RECT MASK 1 127.586 106.38 127.646 107.43 ;
      RECT MASK 1 1.454 107.845 44.382 107.885 ;
      RECT MASK 1 44.846 107.845 87.774 107.885 ;
      RECT MASK 1 88.238 107.845 128.51 107.885 ;
      RECT MASK 2 57.7415 0.62 65.984 0.66 ;
      RECT MASK 2 57.7415 0.78 65.984 0.82 ;
      RECT MASK 2 49.9395 1.04 52.6895 1.08 ;
      RECT MASK 2 58.6465 1.05 58.85 1.078 ;
      RECT MASK 2 59.656 1.05 60.775 1.078 ;
      RECT MASK 2 63.2265 1.05 63.888 1.078 ;
      RECT MASK 2 58.994 1.198 59.054 1.378 ;
      RECT MASK 2 59.452 1.198 59.512 1.378 ;
      RECT MASK 2 61.055 1.198 61.115 1.378 ;
      RECT MASK 2 61.513 1.198 61.573 1.378 ;
      RECT MASK 2 61.971 1.198 62.031 1.378 ;
      RECT MASK 2 62.429 1.198 62.489 1.378 ;
      RECT MASK 2 62.887 1.198 62.947 1.378 ;
      RECT MASK 2 64.032 1.198 64.092 1.378 ;
      RECT MASK 2 64.49 1.198 64.55 1.378 ;
      RECT MASK 2 64.948 1.198 65.008 1.378 ;
      RECT MASK 2 49.9395 1.2 52.6895 1.24 ;
      RECT MASK 2 115.425 1.34 129.001 1.38 ;
      RECT MASK 2 57.789 1.3825 57.969 1.4225 ;
      RECT MASK 2 60.1675 1.3825 60.3475 1.4225 ;
      RECT MASK 2 65.575 1.3825 65.984 1.4225 ;
      RECT MASK 2 115.425 1.53 129.001 1.57 ;
      RECT MASK 2 49.9465 1.54 52.6925 1.58 ;
      RECT MASK 2 1.6805 1.55 10.7245 1.59 ;
      RECT MASK 2 11.1705 1.55 12.9295 1.59 ;
      RECT MASK 2 13.4005 1.55 21.7575 1.59 ;
      RECT MASK 2 25.1795 1.55 33.5365 1.59 ;
      RECT MASK 2 34.0075 1.55 35.7665 1.59 ;
      RECT MASK 2 36.2125 1.55 45.2565 1.59 ;
      RECT MASK 2 58.74 1.619 59.766 1.659 ;
      RECT MASK 2 60.9255 1.619 63.0765 1.659 ;
      RECT MASK 2 63.778 1.619 64.9085 1.659 ;
      RECT MASK 2 49.9465 1.7 52.6825 1.74 ;
      RECT MASK 2 1.6805 1.71 10.7245 1.75 ;
      RECT MASK 2 11.1705 1.71 12.9295 1.75 ;
      RECT MASK 2 13.4005 1.71 21.7575 1.75 ;
      RECT MASK 2 25.1795 1.71 33.5365 1.75 ;
      RECT MASK 2 34.0075 1.71 35.7665 1.75 ;
      RECT MASK 2 36.2125 1.71 45.2565 1.75 ;
      RECT MASK 2 58.74 1.821 59.766 1.861 ;
      RECT MASK 2 60.9255 1.821 63.0765 1.861 ;
      RECT MASK 2 63.778 1.821 64.9085 1.861 ;
      RECT MASK 2 116.291 1.89 116.351 2.94 ;
      RECT MASK 2 116.565 1.89 116.625 2.94 ;
      RECT MASK 2 116.839 1.89 116.899 2.94 ;
      RECT MASK 2 117.113 1.89 117.173 2.94 ;
      RECT MASK 2 117.387 1.89 117.447 2.94 ;
      RECT MASK 2 117.661 1.89 117.721 2.94 ;
      RECT MASK 2 117.935 1.89 117.995 2.94 ;
      RECT MASK 2 118.209 1.89 118.269 2.94 ;
      RECT MASK 2 118.483 1.89 118.543 2.94 ;
      RECT MASK 2 118.757 1.89 118.817 2.94 ;
      RECT MASK 2 119.031 1.89 119.091 2.94 ;
      RECT MASK 2 119.305 1.89 119.365 2.94 ;
      RECT MASK 2 119.579 1.89 119.639 2.94 ;
      RECT MASK 2 119.853 1.89 119.913 2.94 ;
      RECT MASK 2 120.127 1.89 120.187 2.94 ;
      RECT MASK 2 120.401 1.89 120.461 2.94 ;
      RECT MASK 2 120.675 1.89 120.735 2.94 ;
      RECT MASK 2 120.949 1.89 121.009 2.94 ;
      RECT MASK 2 121.223 1.89 121.283 2.94 ;
      RECT MASK 2 121.497 1.89 121.557 2.94 ;
      RECT MASK 2 121.771 1.89 121.831 2.94 ;
      RECT MASK 2 122.045 1.89 122.105 2.94 ;
      RECT MASK 2 122.319 1.89 122.379 2.94 ;
      RECT MASK 2 122.593 1.89 122.653 2.94 ;
      RECT MASK 2 122.867 1.89 122.927 2.94 ;
      RECT MASK 2 123.141 1.89 123.201 2.94 ;
      RECT MASK 2 123.415 1.89 123.475 2.94 ;
      RECT MASK 2 123.689 1.89 123.749 2.94 ;
      RECT MASK 2 123.963 1.89 124.023 2.94 ;
      RECT MASK 2 124.237 1.89 124.297 2.94 ;
      RECT MASK 2 124.511 1.89 124.571 2.94 ;
      RECT MASK 2 124.785 1.89 124.845 2.94 ;
      RECT MASK 2 125.059 1.89 125.119 2.94 ;
      RECT MASK 2 125.333 1.89 125.393 2.94 ;
      RECT MASK 2 125.607 1.89 125.667 2.94 ;
      RECT MASK 2 125.881 1.89 125.941 2.94 ;
      RECT MASK 2 126.155 1.89 126.215 2.94 ;
      RECT MASK 2 126.429 1.89 126.489 2.94 ;
      RECT MASK 2 126.703 1.89 126.763 2.94 ;
      RECT MASK 2 126.977 1.89 127.037 2.94 ;
      RECT MASK 2 127.251 1.89 127.311 2.94 ;
      RECT MASK 2 127.525 1.89 127.585 2.94 ;
      RECT MASK 2 127.799 1.89 127.859 2.94 ;
      RECT MASK 2 128.073 1.89 128.133 2.94 ;
      RECT MASK 2 49.9465 1.975 52.6825 2.015 ;
      RECT MASK 2 2.2045 1.992 2.4335 2.02 ;
      RECT MASK 2 2.961 1.992 3.28 2.02 ;
      RECT MASK 2 5.251 1.992 5.57 2.02 ;
      RECT MASK 2 8.457 1.992 8.776 2.02 ;
      RECT MASK 2 9.831 1.992 10.0455 2.02 ;
      RECT MASK 2 11.1705 1.992 11.3505 2.02 ;
      RECT MASK 2 11.903 1.992 12.222 2.02 ;
      RECT MASK 2 12.7735 1.992 12.9535 2.02 ;
      RECT MASK 2 14.3195 1.992 14.534 2.02 ;
      RECT MASK 2 21.543 1.992 21.7575 2.02 ;
      RECT MASK 2 25.1795 1.992 25.394 2.02 ;
      RECT MASK 2 32.403 1.992 32.6175 2.02 ;
      RECT MASK 2 33.9835 1.992 34.1635 2.02 ;
      RECT MASK 2 34.715 1.992 35.034 2.02 ;
      RECT MASK 2 35.5865 1.992 35.7665 2.02 ;
      RECT MASK 2 36.8915 1.992 37.106 2.02 ;
      RECT MASK 2 38.161 1.992 38.48 2.02 ;
      RECT MASK 2 41.367 1.992 41.686 2.02 ;
      RECT MASK 2 43.657 1.992 43.976 2.02 ;
      RECT MASK 2 44.5035 1.992 44.7325 2.02 ;
      RECT MASK 2 57.789 2.0575 57.969 2.0975 ;
      RECT MASK 2 58.994 2.102 59.054 2.282 ;
      RECT MASK 2 59.452 2.102 59.512 2.282 ;
      RECT MASK 2 61.055 2.102 61.115 2.282 ;
      RECT MASK 2 61.513 2.102 61.573 2.282 ;
      RECT MASK 2 61.971 2.102 62.031 2.282 ;
      RECT MASK 2 62.429 2.102 62.489 2.282 ;
      RECT MASK 2 62.887 2.102 62.947 2.282 ;
      RECT MASK 2 64.032 2.102 64.092 2.282 ;
      RECT MASK 2 64.49 2.102 64.55 2.282 ;
      RECT MASK 2 64.948 2.102 65.008 2.282 ;
      RECT MASK 2 2.6325 2.128 2.6925 2.308 ;
      RECT MASK 2 11.5745 2.128 11.6345 2.308 ;
      RECT MASK 2 12.4905 2.128 12.5505 2.308 ;
      RECT MASK 2 14.8025 2.128 14.8625 2.308 ;
      RECT MASK 2 15.2605 2.128 15.3205 2.308 ;
      RECT MASK 2 15.7185 2.128 15.7785 2.308 ;
      RECT MASK 2 16.1765 2.128 16.2365 2.308 ;
      RECT MASK 2 16.6345 2.128 16.6945 2.308 ;
      RECT MASK 2 17.0925 2.128 17.1525 2.308 ;
      RECT MASK 2 17.5505 2.128 17.6105 2.308 ;
      RECT MASK 2 18.0085 2.128 18.0685 2.308 ;
      RECT MASK 2 18.4665 2.128 18.5265 2.308 ;
      RECT MASK 2 18.9245 2.128 18.9845 2.308 ;
      RECT MASK 2 19.3825 2.128 19.4425 2.308 ;
      RECT MASK 2 19.8405 2.128 19.9005 2.308 ;
      RECT MASK 2 20.2985 2.128 20.3585 2.308 ;
      RECT MASK 2 20.7565 2.128 20.8165 2.308 ;
      RECT MASK 2 21.2145 2.128 21.2745 2.308 ;
      RECT MASK 2 25.6625 2.128 25.7225 2.308 ;
      RECT MASK 2 26.1205 2.128 26.1805 2.308 ;
      RECT MASK 2 26.5785 2.128 26.6385 2.308 ;
      RECT MASK 2 27.0365 2.128 27.0965 2.308 ;
      RECT MASK 2 27.4945 2.128 27.5545 2.308 ;
      RECT MASK 2 27.9525 2.128 28.0125 2.308 ;
      RECT MASK 2 28.4105 2.128 28.4705 2.308 ;
      RECT MASK 2 28.8685 2.128 28.9285 2.308 ;
      RECT MASK 2 29.3265 2.128 29.3865 2.308 ;
      RECT MASK 2 29.7845 2.128 29.8445 2.308 ;
      RECT MASK 2 30.2425 2.128 30.3025 2.308 ;
      RECT MASK 2 30.7005 2.128 30.7605 2.308 ;
      RECT MASK 2 31.1585 2.128 31.2185 2.308 ;
      RECT MASK 2 31.6165 2.128 31.6765 2.308 ;
      RECT MASK 2 32.0745 2.128 32.1345 2.308 ;
      RECT MASK 2 34.3865 2.128 34.4465 2.308 ;
      RECT MASK 2 35.3025 2.128 35.3625 2.308 ;
      RECT MASK 2 44.2445 2.128 44.3045 2.308 ;
      RECT MASK 2 50.1885 2.135 50.4485 2.175 ;
      RECT MASK 2 50.8525 2.135 51.1125 2.175 ;
      RECT MASK 2 51.5165 2.135 51.7765 2.175 ;
      RECT MASK 2 52.1805 2.135 52.4405 2.175 ;
      RECT MASK 2 46.6605 2.16 49.2605 2.18 ;
      RECT MASK 2 60.1675 2.1775 60.3475 2.2175 ;
      RECT MASK 2 65.575 2.1775 65.984 2.2175 ;
      RECT MASK 2 22.2135 2.193 23.3235 2.217 ;
      RECT MASK 2 23.6135 2.193 24.7235 2.217 ;
      RECT MASK 2 46.6605 2.24 49.2605 2.26 ;
      RECT MASK 2 22.2135 2.283 23.3235 2.307 ;
      RECT MASK 2 23.6135 2.283 24.7235 2.307 ;
      RECT MASK 2 10.3585 2.3125 10.5385 2.3525 ;
      RECT MASK 2 13.5865 2.3125 13.7665 2.3525 ;
      RECT MASK 2 33.1705 2.3125 33.3505 2.3525 ;
      RECT MASK 2 36.3985 2.3125 36.5785 2.3525 ;
      RECT MASK 2 46.6605 2.32 49.2605 2.34 ;
      RECT MASK 2 1.6135 2.3725 1.8575 2.4125 ;
      RECT MASK 2 45.0795 2.3725 45.3235 2.4125 ;
      RECT MASK 2 22.2135 2.373 23.3235 2.397 ;
      RECT MASK 2 23.6135 2.373 24.7235 2.397 ;
      RECT MASK 2 46.6605 2.4 49.2605 2.42 ;
      RECT MASK 2 58.6465 2.402 58.85 2.43 ;
      RECT MASK 2 59.656 2.402 60.775 2.43 ;
      RECT MASK 2 63.2265 2.402 63.888 2.43 ;
      RECT MASK 2 2.3785 2.448 2.8505 2.488 ;
      RECT MASK 2 3.3985 2.448 3.738 2.488 ;
      RECT MASK 2 4.3185 2.448 5.4655 2.488 ;
      RECT MASK 2 5.938 2.448 6.3815 2.488 ;
      RECT MASK 2 6.854 2.448 7.2975 2.488 ;
      RECT MASK 2 7.77 2.448 8.6715 2.488 ;
      RECT MASK 2 8.915 2.448 10.1875 2.488 ;
      RECT MASK 2 36.7495 2.448 38.022 2.488 ;
      RECT MASK 2 38.2655 2.448 39.167 2.488 ;
      RECT MASK 2 39.6395 2.448 40.083 2.488 ;
      RECT MASK 2 40.5555 2.448 40.999 2.488 ;
      RECT MASK 2 41.4715 2.448 42.6185 2.488 ;
      RECT MASK 2 43.199 2.448 43.5385 2.488 ;
      RECT MASK 2 44.0865 2.448 44.5585 2.488 ;
      RECT MASK 2 46.6605 2.48 49.2605 2.5 ;
      RECT MASK 2 49.9395 2.51 52.6895 2.55 ;
      RECT MASK 2 46.6605 2.56 49.2605 2.58 ;
      RECT MASK 2 58.4175 2.61 58.621 2.638 ;
      RECT MASK 2 60.343 2.61 60.546 2.638 ;
      RECT MASK 2 49.9395 2.67 52.6895 2.71 ;
      RECT MASK 2 22.3735 2.733 22.7635 2.757 ;
      RECT MASK 2 24.1735 2.733 24.5635 2.757 ;
      RECT MASK 2 58.765 2.758 58.825 2.938 ;
      RECT MASK 2 59.223 2.758 59.283 2.938 ;
      RECT MASK 2 59.681 2.758 59.741 2.938 ;
      RECT MASK 2 60.139 2.758 60.199 2.938 ;
      RECT MASK 2 62.658 2.758 62.718 2.938 ;
      RECT MASK 2 63.116 2.758 63.176 2.938 ;
      RECT MASK 2 63.574 2.758 63.634 2.938 ;
      RECT MASK 2 64.032 2.758 64.092 2.938 ;
      RECT MASK 2 64.49 2.758 64.55 2.938 ;
      RECT MASK 2 64.948 2.758 65.008 2.938 ;
      RECT MASK 2 65.406 2.758 65.466 2.938 ;
      RECT MASK 2 65.864 2.758 65.924 2.938 ;
      RECT MASK 2 60.995 2.8225 61.404 2.8625 ;
      RECT MASK 2 61.911 2.8225 62.091 2.8625 ;
      RECT MASK 2 22.2135 2.823 23.3235 2.847 ;
      RECT MASK 2 23.6135 2.823 24.7235 2.847 ;
      RECT MASK 2 2.3785 2.852 2.8505 2.892 ;
      RECT MASK 2 3.3985 2.852 3.738 2.892 ;
      RECT MASK 2 4.3185 2.852 5.4655 2.892 ;
      RECT MASK 2 5.938 2.852 6.3815 2.892 ;
      RECT MASK 2 6.854 2.852 7.2975 2.892 ;
      RECT MASK 2 7.77 2.852 8.6715 2.892 ;
      RECT MASK 2 12.361 2.852 13.0765 2.892 ;
      RECT MASK 2 33.8605 2.852 34.576 2.892 ;
      RECT MASK 2 38.2655 2.852 39.167 2.892 ;
      RECT MASK 2 39.6395 2.852 40.083 2.892 ;
      RECT MASK 2 40.5555 2.852 40.999 2.892 ;
      RECT MASK 2 41.4715 2.852 42.6185 2.892 ;
      RECT MASK 2 43.199 2.852 43.5385 2.892 ;
      RECT MASK 2 44.0865 2.852 44.5585 2.892 ;
      RECT MASK 2 46.6605 2.88 49.2605 2.9 ;
      RECT MASK 2 22.4135 2.913 22.7135 2.937 ;
      RECT MASK 2 22.8235 2.913 23.1235 2.937 ;
      RECT MASK 2 23.8135 2.913 24.1135 2.937 ;
      RECT MASK 2 24.2235 2.913 24.5235 2.937 ;
      RECT MASK 2 1.6135 2.9275 1.8575 2.9675 ;
      RECT MASK 2 45.0795 2.9275 45.3235 2.9675 ;
      RECT MASK 2 49.9395 2.93 52.6895 2.97 ;
      RECT MASK 2 57.789 2.9425 57.969 2.9825 ;
      RECT MASK 2 46.6605 2.96 49.2605 2.98 ;
      RECT MASK 2 10.107 2.9875 10.7505 3.0275 ;
      RECT MASK 2 13.5865 2.9875 13.7665 3.0275 ;
      RECT MASK 2 33.1705 2.9875 33.3505 3.0275 ;
      RECT MASK 2 36.3985 2.9875 36.5785 3.0275 ;
      RECT MASK 2 22.4135 3.003 22.7135 3.027 ;
      RECT MASK 2 22.8235 3.003 23.1235 3.027 ;
      RECT MASK 2 23.8135 3.003 24.1135 3.027 ;
      RECT MASK 2 24.2235 3.003 24.5235 3.027 ;
      RECT MASK 2 2.6325 3.032 2.6925 3.212 ;
      RECT MASK 2 11.5745 3.032 11.6345 3.212 ;
      RECT MASK 2 12.4905 3.032 12.5505 3.212 ;
      RECT MASK 2 14.8025 3.032 14.8625 3.212 ;
      RECT MASK 2 15.2605 3.032 15.3205 3.212 ;
      RECT MASK 2 15.7185 3.032 15.7785 3.212 ;
      RECT MASK 2 16.1765 3.032 16.2365 3.212 ;
      RECT MASK 2 16.6345 3.032 16.6945 3.212 ;
      RECT MASK 2 17.0925 3.032 17.1525 3.212 ;
      RECT MASK 2 17.5505 3.032 17.6105 3.212 ;
      RECT MASK 2 18.0085 3.032 18.0685 3.212 ;
      RECT MASK 2 18.4665 3.032 18.5265 3.212 ;
      RECT MASK 2 18.9245 3.032 18.9845 3.212 ;
      RECT MASK 2 19.3825 3.032 19.4425 3.212 ;
      RECT MASK 2 19.8405 3.032 19.9005 3.212 ;
      RECT MASK 2 20.2985 3.032 20.3585 3.212 ;
      RECT MASK 2 20.7565 3.032 20.8165 3.212 ;
      RECT MASK 2 21.2145 3.032 21.2745 3.212 ;
      RECT MASK 2 25.6625 3.032 25.7225 3.212 ;
      RECT MASK 2 26.1205 3.032 26.1805 3.212 ;
      RECT MASK 2 26.5785 3.032 26.6385 3.212 ;
      RECT MASK 2 27.0365 3.032 27.0965 3.212 ;
      RECT MASK 2 27.4945 3.032 27.5545 3.212 ;
      RECT MASK 2 27.9525 3.032 28.0125 3.212 ;
      RECT MASK 2 28.4105 3.032 28.4705 3.212 ;
      RECT MASK 2 28.8685 3.032 28.9285 3.212 ;
      RECT MASK 2 29.3265 3.032 29.3865 3.212 ;
      RECT MASK 2 29.7845 3.032 29.8445 3.212 ;
      RECT MASK 2 30.2425 3.032 30.3025 3.212 ;
      RECT MASK 2 30.7005 3.032 30.7605 3.212 ;
      RECT MASK 2 31.1585 3.032 31.2185 3.212 ;
      RECT MASK 2 31.6165 3.032 31.6765 3.212 ;
      RECT MASK 2 32.0745 3.032 32.1345 3.212 ;
      RECT MASK 2 34.3865 3.032 34.4465 3.212 ;
      RECT MASK 2 35.3025 3.032 35.3625 3.212 ;
      RECT MASK 2 44.2445 3.032 44.3045 3.212 ;
      RECT MASK 2 46.6605 3.04 49.2605 3.06 ;
      RECT MASK 2 49.9395 3.09 52.6895 3.13 ;
      RECT MASK 2 22.4135 3.093 22.7135 3.117 ;
      RECT MASK 2 22.8235 3.093 23.1235 3.117 ;
      RECT MASK 2 23.8135 3.093 24.1135 3.117 ;
      RECT MASK 2 24.2235 3.093 24.5235 3.117 ;
      RECT MASK 2 46.6605 3.12 49.2605 3.14 ;
      RECT MASK 2 58.6355 3.179 59.4225 3.219 ;
      RECT MASK 2 59.5415 3.179 60.3285 3.219 ;
      RECT MASK 2 62.862 3.179 64.4505 3.219 ;
      RECT MASK 2 64.5795 3.179 64.9085 3.219 ;
      RECT MASK 2 46.6605 3.2 49.2605 3.22 ;
      RECT MASK 2 46.6605 3.28 49.2605 3.3 ;
      RECT MASK 2 2.2045 3.32 2.4335 3.348 ;
      RECT MASK 2 2.961 3.32 3.28 3.348 ;
      RECT MASK 2 5.251 3.32 5.57 3.348 ;
      RECT MASK 2 8.457 3.32 8.776 3.348 ;
      RECT MASK 2 9.831 3.32 10.0455 3.348 ;
      RECT MASK 2 11.1705 3.32 11.3505 3.348 ;
      RECT MASK 2 11.903 3.32 12.222 3.348 ;
      RECT MASK 2 12.7735 3.32 12.9535 3.348 ;
      RECT MASK 2 14.3195 3.32 14.534 3.348 ;
      RECT MASK 2 21.543 3.32 21.7575 3.348 ;
      RECT MASK 2 25.1795 3.32 25.394 3.348 ;
      RECT MASK 2 32.403 3.32 32.6175 3.348 ;
      RECT MASK 2 33.9835 3.32 34.1635 3.348 ;
      RECT MASK 2 34.715 3.32 35.034 3.348 ;
      RECT MASK 2 35.5865 3.32 35.7665 3.348 ;
      RECT MASK 2 36.8915 3.32 37.106 3.348 ;
      RECT MASK 2 38.161 3.32 38.48 3.348 ;
      RECT MASK 2 41.367 3.32 41.686 3.348 ;
      RECT MASK 2 43.657 3.32 43.976 3.348 ;
      RECT MASK 2 44.5035 3.32 44.7325 3.348 ;
      RECT MASK 2 58.4065 3.381 58.9545 3.421 ;
      RECT MASK 2 59.0935 3.381 59.4225 3.421 ;
      RECT MASK 2 59.5415 3.381 59.8705 3.421 ;
      RECT MASK 2 60.0095 3.381 60.5575 3.421 ;
      RECT MASK 2 62.862 3.381 63.557 3.421 ;
      RECT MASK 2 63.6735 3.381 64.473 3.421 ;
      RECT MASK 2 64.8185 3.381 65.491 3.421 ;
      RECT MASK 2 22.2235 3.438 23.3135 3.462 ;
      RECT MASK 2 23.6235 3.438 24.7135 3.462 ;
      RECT MASK 2 49.9415 3.45 52.6875 3.51 ;
      RECT MASK 2 72.7245 3.56 76.9845 3.6 ;
      RECT MASK 2 77.4385 3.56 82.3625 3.6 ;
      RECT MASK 2 104.3425 3.56 109.2665 3.6 ;
      RECT MASK 2 109.7205 3.56 113.9805 3.6 ;
      RECT MASK 2 1.6805 3.59 13.9525 3.63 ;
      RECT MASK 2 14.3195 3.59 21.7575 3.63 ;
      RECT MASK 2 25.1795 3.59 32.6175 3.63 ;
      RECT MASK 2 32.9845 3.59 45.2565 3.63 ;
      RECT MASK 2 46.6605 3.6 49.2605 3.62 ;
      RECT MASK 2 116.291 3.6 116.351 4.65 ;
      RECT MASK 2 116.565 3.6 116.625 4.65 ;
      RECT MASK 2 116.839 3.6 116.899 4.65 ;
      RECT MASK 2 117.113 3.6 117.173 4.65 ;
      RECT MASK 2 117.387 3.6 117.447 4.65 ;
      RECT MASK 2 117.661 3.6 117.721 4.65 ;
      RECT MASK 2 117.935 3.6 117.995 4.65 ;
      RECT MASK 2 118.209 3.6 118.269 4.65 ;
      RECT MASK 2 118.483 3.6 118.543 4.65 ;
      RECT MASK 2 118.757 3.6 118.817 4.65 ;
      RECT MASK 2 119.031 3.6 119.091 4.65 ;
      RECT MASK 2 119.305 3.6 119.365 4.65 ;
      RECT MASK 2 119.579 3.6 119.639 4.65 ;
      RECT MASK 2 119.853 3.6 119.913 4.65 ;
      RECT MASK 2 120.127 3.6 120.187 4.65 ;
      RECT MASK 2 120.401 3.6 120.461 4.65 ;
      RECT MASK 2 120.675 3.6 120.735 4.65 ;
      RECT MASK 2 120.949 3.6 121.009 4.65 ;
      RECT MASK 2 121.223 3.6 121.283 4.65 ;
      RECT MASK 2 121.497 3.6 121.557 4.65 ;
      RECT MASK 2 121.771 3.6 121.831 4.65 ;
      RECT MASK 2 122.045 3.6 122.105 4.65 ;
      RECT MASK 2 122.319 3.6 122.379 4.65 ;
      RECT MASK 2 122.593 3.6 122.653 4.65 ;
      RECT MASK 2 122.867 3.6 122.927 4.65 ;
      RECT MASK 2 123.141 3.6 123.201 4.65 ;
      RECT MASK 2 123.415 3.6 123.475 4.65 ;
      RECT MASK 2 123.689 3.6 123.749 4.65 ;
      RECT MASK 2 123.963 3.6 124.023 4.65 ;
      RECT MASK 2 124.237 3.6 124.297 4.65 ;
      RECT MASK 2 124.511 3.6 124.571 4.65 ;
      RECT MASK 2 124.785 3.6 124.845 4.65 ;
      RECT MASK 2 125.059 3.6 125.119 4.65 ;
      RECT MASK 2 125.333 3.6 125.393 4.65 ;
      RECT MASK 2 125.607 3.6 125.667 4.65 ;
      RECT MASK 2 125.881 3.6 125.941 4.65 ;
      RECT MASK 2 126.155 3.6 126.215 4.65 ;
      RECT MASK 2 126.429 3.6 126.489 4.65 ;
      RECT MASK 2 126.703 3.6 126.763 4.65 ;
      RECT MASK 2 126.977 3.6 127.037 4.65 ;
      RECT MASK 2 127.251 3.6 127.311 4.65 ;
      RECT MASK 2 127.525 3.6 127.585 4.65 ;
      RECT MASK 2 127.799 3.6 127.859 4.65 ;
      RECT MASK 2 128.073 3.6 128.133 4.65 ;
      RECT MASK 2 57.789 3.6175 57.969 3.6575 ;
      RECT MASK 2 60.995 3.6175 61.404 3.6575 ;
      RECT MASK 2 61.911 3.6175 62.091 3.6575 ;
      RECT MASK 2 58.765 3.662 58.825 3.842 ;
      RECT MASK 2 59.223 3.662 59.283 3.842 ;
      RECT MASK 2 59.681 3.662 59.741 3.842 ;
      RECT MASK 2 60.139 3.662 60.199 3.842 ;
      RECT MASK 2 62.658 3.662 62.718 3.842 ;
      RECT MASK 2 63.116 3.662 63.176 3.842 ;
      RECT MASK 2 63.574 3.662 63.634 3.842 ;
      RECT MASK 2 64.032 3.662 64.092 3.842 ;
      RECT MASK 2 64.49 3.662 64.55 3.842 ;
      RECT MASK 2 64.948 3.662 65.008 3.842 ;
      RECT MASK 2 65.406 3.662 65.466 3.842 ;
      RECT MASK 2 65.864 3.662 65.924 3.842 ;
      RECT MASK 2 46.6605 3.68 49.2605 3.7 ;
      RECT MASK 2 49.9415 3.69 52.6875 3.75 ;
      RECT MASK 2 72.7245 3.72 76.9845 3.76 ;
      RECT MASK 2 77.4385 3.72 82.3625 3.76 ;
      RECT MASK 2 104.3425 3.72 109.2665 3.76 ;
      RECT MASK 2 109.7205 3.72 113.9805 3.76 ;
      RECT MASK 2 1.6805 3.75 13.9525 3.79 ;
      RECT MASK 2 14.3195 3.75 21.7575 3.79 ;
      RECT MASK 2 25.1795 3.75 32.6175 3.79 ;
      RECT MASK 2 32.9845 3.75 45.2565 3.79 ;
      RECT MASK 2 46.6605 3.76 49.2605 3.78 ;
      RECT MASK 2 83.7885 3.8 93.0585 3.84 ;
      RECT MASK 2 93.6465 3.8 102.9165 3.84 ;
      RECT MASK 2 46.6605 3.84 49.2605 3.86 ;
      RECT MASK 2 22.2235 3.918 23.3135 3.942 ;
      RECT MASK 2 23.6235 3.918 24.7135 3.942 ;
      RECT MASK 2 46.6605 3.92 49.2605 3.94 ;
      RECT MASK 2 49.9415 3.93 52.6875 3.99 ;
      RECT MASK 2 83.7885 3.96 93.0585 4 ;
      RECT MASK 2 93.6465 3.96 102.9165 4 ;
      RECT MASK 2 46.6605 4 49.2605 4.02 ;
      RECT MASK 2 2.2045 4.032 2.4335 4.06 ;
      RECT MASK 2 2.961 4.032 3.28 4.06 ;
      RECT MASK 2 5.251 4.032 5.57 4.06 ;
      RECT MASK 2 8.457 4.032 8.776 4.06 ;
      RECT MASK 2 9.831 4.032 10.0455 4.06 ;
      RECT MASK 2 11.1705 4.032 11.3505 4.06 ;
      RECT MASK 2 11.903 4.032 12.222 4.06 ;
      RECT MASK 2 12.7735 4.032 12.9535 4.06 ;
      RECT MASK 2 14.3195 4.032 14.534 4.06 ;
      RECT MASK 2 21.543 4.032 21.7575 4.06 ;
      RECT MASK 2 25.1795 4.032 25.394 4.06 ;
      RECT MASK 2 32.403 4.032 32.6175 4.06 ;
      RECT MASK 2 33.9835 4.032 34.1635 4.06 ;
      RECT MASK 2 34.715 4.032 35.034 4.06 ;
      RECT MASK 2 35.5865 4.032 35.7665 4.06 ;
      RECT MASK 2 36.8915 4.032 37.106 4.06 ;
      RECT MASK 2 38.161 4.032 38.48 4.06 ;
      RECT MASK 2 41.367 4.032 41.686 4.06 ;
      RECT MASK 2 43.657 4.032 43.976 4.06 ;
      RECT MASK 2 44.5035 4.032 44.7325 4.06 ;
      RECT MASK 2 73.8505 4.159 74.2885 4.339 ;
      RECT MASK 2 74.6165 4.159 75.1445 4.339 ;
      RECT MASK 2 75.4725 4.159 75.9105 4.339 ;
      RECT MASK 2 78.5035 4.159 78.9415 4.339 ;
      RECT MASK 2 79.2695 4.159 79.7575 4.339 ;
      RECT MASK 2 80.0855 4.159 80.5535 4.339 ;
      RECT MASK 2 80.8815 4.159 81.3195 4.339 ;
      RECT MASK 2 105.3855 4.159 105.8235 4.339 ;
      RECT MASK 2 106.1515 4.159 106.6195 4.339 ;
      RECT MASK 2 106.9475 4.159 107.4355 4.339 ;
      RECT MASK 2 107.7635 4.159 108.2015 4.339 ;
      RECT MASK 2 110.7945 4.159 111.2325 4.339 ;
      RECT MASK 2 111.5605 4.159 112.0885 4.339 ;
      RECT MASK 2 112.4165 4.159 112.8545 4.339 ;
      RECT MASK 2 2.6325 4.168 2.6925 4.348 ;
      RECT MASK 2 11.5745 4.168 11.6345 4.348 ;
      RECT MASK 2 12.4905 4.168 12.5505 4.348 ;
      RECT MASK 2 14.8025 4.168 14.8625 4.348 ;
      RECT MASK 2 15.2605 4.168 15.3205 4.348 ;
      RECT MASK 2 15.7185 4.168 15.7785 4.348 ;
      RECT MASK 2 16.1765 4.168 16.2365 4.348 ;
      RECT MASK 2 16.6345 4.168 16.6945 4.348 ;
      RECT MASK 2 17.0925 4.168 17.1525 4.348 ;
      RECT MASK 2 17.5505 4.168 17.6105 4.348 ;
      RECT MASK 2 18.0085 4.168 18.0685 4.348 ;
      RECT MASK 2 18.4665 4.168 18.5265 4.348 ;
      RECT MASK 2 18.9245 4.168 18.9845 4.348 ;
      RECT MASK 2 19.3825 4.168 19.4425 4.348 ;
      RECT MASK 2 19.8405 4.168 19.9005 4.348 ;
      RECT MASK 2 20.2985 4.168 20.3585 4.348 ;
      RECT MASK 2 20.7565 4.168 20.8165 4.348 ;
      RECT MASK 2 21.2145 4.168 21.2745 4.348 ;
      RECT MASK 2 25.6625 4.168 25.7225 4.348 ;
      RECT MASK 2 26.1205 4.168 26.1805 4.348 ;
      RECT MASK 2 26.5785 4.168 26.6385 4.348 ;
      RECT MASK 2 27.0365 4.168 27.0965 4.348 ;
      RECT MASK 2 27.4945 4.168 27.5545 4.348 ;
      RECT MASK 2 27.9525 4.168 28.0125 4.348 ;
      RECT MASK 2 28.4105 4.168 28.4705 4.348 ;
      RECT MASK 2 28.8685 4.168 28.9285 4.348 ;
      RECT MASK 2 29.3265 4.168 29.3865 4.348 ;
      RECT MASK 2 29.7845 4.168 29.8445 4.348 ;
      RECT MASK 2 30.2425 4.168 30.3025 4.348 ;
      RECT MASK 2 30.7005 4.168 30.7605 4.348 ;
      RECT MASK 2 31.1585 4.168 31.2185 4.348 ;
      RECT MASK 2 31.6165 4.168 31.6765 4.348 ;
      RECT MASK 2 32.0745 4.168 32.1345 4.348 ;
      RECT MASK 2 34.3865 4.168 34.4465 4.348 ;
      RECT MASK 2 35.3025 4.168 35.3625 4.348 ;
      RECT MASK 2 44.2445 4.168 44.3045 4.348 ;
      RECT MASK 2 49.9735 4.2 50.3705 4.26 ;
      RECT MASK 2 50.6375 4.2 51.0345 4.26 ;
      RECT MASK 2 51.3015 4.2 51.6985 4.26 ;
      RECT MASK 2 51.9655 4.2 52.3625 4.26 ;
      RECT MASK 2 52.6025 4.2 52.7825 4.26 ;
      RECT MASK 2 22.4135 4.263 22.7135 4.287 ;
      RECT MASK 2 22.8235 4.263 23.1235 4.287 ;
      RECT MASK 2 23.8135 4.263 24.1135 4.287 ;
      RECT MASK 2 24.2235 4.263 24.5235 4.287 ;
      RECT MASK 2 58.765 4.318 58.825 4.498 ;
      RECT MASK 2 59.223 4.318 59.283 4.498 ;
      RECT MASK 2 59.681 4.318 59.741 4.498 ;
      RECT MASK 2 60.139 4.318 60.199 4.498 ;
      RECT MASK 2 62.658 4.318 62.718 4.498 ;
      RECT MASK 2 63.116 4.318 63.176 4.498 ;
      RECT MASK 2 63.574 4.318 63.634 4.498 ;
      RECT MASK 2 64.032 4.318 64.092 4.498 ;
      RECT MASK 2 64.49 4.318 64.55 4.498 ;
      RECT MASK 2 64.948 4.318 65.008 4.498 ;
      RECT MASK 2 65.406 4.318 65.466 4.498 ;
      RECT MASK 2 65.864 4.318 65.924 4.498 ;
      RECT MASK 2 10.107 4.3525 10.7505 4.3925 ;
      RECT MASK 2 13.5865 4.3525 13.7665 4.3925 ;
      RECT MASK 2 33.1705 4.3525 33.3505 4.3925 ;
      RECT MASK 2 36.3985 4.3525 36.5785 4.3925 ;
      RECT MASK 2 22.4135 4.353 22.7135 4.377 ;
      RECT MASK 2 22.8235 4.353 23.1235 4.377 ;
      RECT MASK 2 23.8135 4.353 24.1135 4.377 ;
      RECT MASK 2 24.2235 4.353 24.5235 4.377 ;
      RECT MASK 2 49.9735 4.38 50.3575 4.44 ;
      RECT MASK 2 50.6375 4.38 51.0215 4.44 ;
      RECT MASK 2 51.3015 4.38 51.6855 4.44 ;
      RECT MASK 2 51.9655 4.38 52.3495 4.44 ;
      RECT MASK 2 52.6025 4.38 52.7825 4.44 ;
      RECT MASK 2 1.6135 4.4125 1.8575 4.4525 ;
      RECT MASK 2 45.0795 4.4125 45.3235 4.4525 ;
      RECT MASK 2 22.4135 4.443 22.7135 4.467 ;
      RECT MASK 2 22.8235 4.443 23.1235 4.467 ;
      RECT MASK 2 23.8135 4.443 24.1135 4.467 ;
      RECT MASK 2 24.2235 4.443 24.5235 4.467 ;
      RECT MASK 2 2.3785 4.488 2.8505 4.528 ;
      RECT MASK 2 3.3985 4.488 3.738 4.528 ;
      RECT MASK 2 4.3185 4.488 5.4655 4.528 ;
      RECT MASK 2 5.938 4.488 6.3815 4.528 ;
      RECT MASK 2 6.854 4.488 7.2975 4.528 ;
      RECT MASK 2 7.77 4.488 8.6715 4.528 ;
      RECT MASK 2 12.361 4.488 13.0765 4.528 ;
      RECT MASK 2 33.8605 4.488 34.576 4.528 ;
      RECT MASK 2 38.2655 4.488 39.167 4.528 ;
      RECT MASK 2 39.6395 4.488 40.083 4.528 ;
      RECT MASK 2 40.5555 4.488 40.999 4.528 ;
      RECT MASK 2 41.4715 4.488 42.6185 4.528 ;
      RECT MASK 2 43.199 4.488 43.5385 4.528 ;
      RECT MASK 2 44.0865 4.488 44.5585 4.528 ;
      RECT MASK 2 84.4855 4.498 88.2395 4.558 ;
      RECT MASK 2 88.6075 4.498 92.3615 4.558 ;
      RECT MASK 2 94.3435 4.498 98.0975 4.558 ;
      RECT MASK 2 98.4655 4.498 102.2195 4.558 ;
      RECT MASK 2 57.789 4.5025 57.969 4.5425 ;
      RECT MASK 2 60.995 4.5025 61.404 4.5425 ;
      RECT MASK 2 61.911 4.5025 62.091 4.5425 ;
      RECT MASK 2 22.2135 4.533 23.3235 4.557 ;
      RECT MASK 2 23.6135 4.533 24.7235 4.557 ;
      RECT MASK 2 22.3735 4.623 22.7635 4.647 ;
      RECT MASK 2 24.1735 4.623 24.5635 4.647 ;
      RECT MASK 2 49.9415 4.65 52.6875 4.71 ;
      RECT MASK 2 58.4065 4.739 58.9545 4.779 ;
      RECT MASK 2 59.0935 4.739 59.4225 4.779 ;
      RECT MASK 2 59.5415 4.739 59.8705 4.779 ;
      RECT MASK 2 60.0095 4.739 60.5575 4.779 ;
      RECT MASK 2 62.862 4.739 63.557 4.779 ;
      RECT MASK 2 63.6735 4.739 64.473 4.779 ;
      RECT MASK 2 64.8185 4.739 65.491 4.779 ;
      RECT MASK 2 84.1235 4.74 84.461 4.8 ;
      RECT MASK 2 84.6 4.74 88.125 4.8 ;
      RECT MASK 2 88.264 4.74 88.583 4.8 ;
      RECT MASK 2 88.722 4.74 92.247 4.8 ;
      RECT MASK 2 92.386 4.74 92.705 4.8 ;
      RECT MASK 2 94 4.74 94.319 4.8 ;
      RECT MASK 2 94.458 4.74 97.983 4.8 ;
      RECT MASK 2 98.122 4.74 98.441 4.8 ;
      RECT MASK 2 98.58 4.74 102.105 4.8 ;
      RECT MASK 2 102.244 4.74 102.5815 4.8 ;
      RECT MASK 2 49.9415 4.89 52.6875 4.95 ;
      RECT MASK 2 2.3785 4.892 2.8505 4.932 ;
      RECT MASK 2 3.3985 4.892 3.738 4.932 ;
      RECT MASK 2 4.3185 4.892 5.4655 4.932 ;
      RECT MASK 2 5.938 4.892 6.3815 4.932 ;
      RECT MASK 2 6.854 4.892 7.2975 4.932 ;
      RECT MASK 2 7.77 4.892 8.6715 4.932 ;
      RECT MASK 2 8.915 4.892 10.1875 4.932 ;
      RECT MASK 2 36.7495 4.892 38.022 4.932 ;
      RECT MASK 2 38.2655 4.892 39.167 4.932 ;
      RECT MASK 2 39.6395 4.892 40.083 4.932 ;
      RECT MASK 2 40.5555 4.892 40.999 4.932 ;
      RECT MASK 2 41.4715 4.892 42.6185 4.932 ;
      RECT MASK 2 43.199 4.892 43.5385 4.932 ;
      RECT MASK 2 44.0865 4.892 44.5585 4.932 ;
      RECT MASK 2 58.6355 4.941 59.4225 4.981 ;
      RECT MASK 2 59.5415 4.941 60.3285 4.981 ;
      RECT MASK 2 62.862 4.941 64.4505 4.981 ;
      RECT MASK 2 64.5795 4.941 64.9085 4.981 ;
      RECT MASK 2 1.6135 4.9675 1.8575 5.0075 ;
      RECT MASK 2 45.0795 4.9675 45.3235 5.0075 ;
      RECT MASK 2 22.2135 4.983 23.3235 5.007 ;
      RECT MASK 2 23.6135 4.983 24.7235 5.007 ;
      RECT MASK 2 10.3585 5.0275 10.5385 5.0675 ;
      RECT MASK 2 13.5865 5.0275 13.7665 5.0675 ;
      RECT MASK 2 33.1705 5.0275 33.3505 5.0675 ;
      RECT MASK 2 36.3985 5.0275 36.5785 5.0675 ;
      RECT MASK 2 2.6325 5.072 2.6925 5.252 ;
      RECT MASK 2 11.5745 5.072 11.6345 5.252 ;
      RECT MASK 2 12.4905 5.072 12.5505 5.252 ;
      RECT MASK 2 14.8025 5.072 14.8625 5.252 ;
      RECT MASK 2 15.2605 5.072 15.3205 5.252 ;
      RECT MASK 2 15.7185 5.072 15.7785 5.252 ;
      RECT MASK 2 16.1765 5.072 16.2365 5.252 ;
      RECT MASK 2 16.6345 5.072 16.6945 5.252 ;
      RECT MASK 2 17.0925 5.072 17.1525 5.252 ;
      RECT MASK 2 17.5505 5.072 17.6105 5.252 ;
      RECT MASK 2 18.0085 5.072 18.0685 5.252 ;
      RECT MASK 2 18.4665 5.072 18.5265 5.252 ;
      RECT MASK 2 18.9245 5.072 18.9845 5.252 ;
      RECT MASK 2 19.3825 5.072 19.4425 5.252 ;
      RECT MASK 2 19.8405 5.072 19.9005 5.252 ;
      RECT MASK 2 20.2985 5.072 20.3585 5.252 ;
      RECT MASK 2 20.7565 5.072 20.8165 5.252 ;
      RECT MASK 2 21.2145 5.072 21.2745 5.252 ;
      RECT MASK 2 25.6625 5.072 25.7225 5.252 ;
      RECT MASK 2 26.1205 5.072 26.1805 5.252 ;
      RECT MASK 2 26.5785 5.072 26.6385 5.252 ;
      RECT MASK 2 27.0365 5.072 27.0965 5.252 ;
      RECT MASK 2 27.4945 5.072 27.5545 5.252 ;
      RECT MASK 2 27.9525 5.072 28.0125 5.252 ;
      RECT MASK 2 28.4105 5.072 28.4705 5.252 ;
      RECT MASK 2 28.8685 5.072 28.9285 5.252 ;
      RECT MASK 2 29.3265 5.072 29.3865 5.252 ;
      RECT MASK 2 29.7845 5.072 29.8445 5.252 ;
      RECT MASK 2 30.2425 5.072 30.3025 5.252 ;
      RECT MASK 2 30.7005 5.072 30.7605 5.252 ;
      RECT MASK 2 31.1585 5.072 31.2185 5.252 ;
      RECT MASK 2 31.6165 5.072 31.6765 5.252 ;
      RECT MASK 2 32.0745 5.072 32.1345 5.252 ;
      RECT MASK 2 34.3865 5.072 34.4465 5.252 ;
      RECT MASK 2 35.3025 5.072 35.3625 5.252 ;
      RECT MASK 2 44.2445 5.072 44.3045 5.252 ;
      RECT MASK 2 22.2135 5.073 23.3235 5.097 ;
      RECT MASK 2 23.6135 5.073 24.7235 5.097 ;
      RECT MASK 2 49.9415 5.13 52.6875 5.19 ;
      RECT MASK 2 46.7745 5.15 48.9595 5.19 ;
      RECT MASK 2 22.2135 5.163 23.3235 5.187 ;
      RECT MASK 2 23.6135 5.163 24.7235 5.187 ;
      RECT MASK 2 57.789 5.1775 57.969 5.2175 ;
      RECT MASK 2 84.7145 5.219 86.3865 5.279 ;
      RECT MASK 2 86.5465 5.219 90.3005 5.279 ;
      RECT MASK 2 90.6685 5.219 92.1325 5.279 ;
      RECT MASK 2 94.5725 5.219 96.0365 5.279 ;
      RECT MASK 2 96.4045 5.219 100.1585 5.279 ;
      RECT MASK 2 100.3185 5.219 101.9905 5.279 ;
      RECT MASK 2 58.765 5.222 58.825 5.402 ;
      RECT MASK 2 59.223 5.222 59.283 5.402 ;
      RECT MASK 2 59.681 5.222 59.741 5.402 ;
      RECT MASK 2 60.139 5.222 60.199 5.402 ;
      RECT MASK 2 62.658 5.222 62.718 5.402 ;
      RECT MASK 2 63.116 5.222 63.176 5.402 ;
      RECT MASK 2 63.574 5.222 63.634 5.402 ;
      RECT MASK 2 64.032 5.222 64.092 5.402 ;
      RECT MASK 2 64.49 5.222 64.55 5.402 ;
      RECT MASK 2 64.948 5.222 65.008 5.402 ;
      RECT MASK 2 65.406 5.222 65.466 5.402 ;
      RECT MASK 2 65.864 5.222 65.924 5.402 ;
      RECT MASK 2 53.9045 5.27 56.1725 5.31 ;
      RECT MASK 2 60.995 5.2975 61.404 5.3375 ;
      RECT MASK 2 61.911 5.2975 62.091 5.3375 ;
      RECT MASK 2 46.7745 5.31 48.9595 5.35 ;
      RECT MASK 2 116.291 5.31 116.351 6.36 ;
      RECT MASK 2 116.565 5.31 116.625 6.36 ;
      RECT MASK 2 116.839 5.31 116.899 6.36 ;
      RECT MASK 2 117.113 5.31 117.173 6.36 ;
      RECT MASK 2 117.387 5.31 117.447 6.36 ;
      RECT MASK 2 117.661 5.31 117.721 6.36 ;
      RECT MASK 2 117.935 5.31 117.995 6.36 ;
      RECT MASK 2 118.209 5.31 118.269 6.36 ;
      RECT MASK 2 118.483 5.31 118.543 6.36 ;
      RECT MASK 2 118.757 5.31 118.817 6.36 ;
      RECT MASK 2 119.031 5.31 119.091 6.36 ;
      RECT MASK 2 119.305 5.31 119.365 6.36 ;
      RECT MASK 2 119.579 5.31 119.639 6.36 ;
      RECT MASK 2 119.853 5.31 119.913 6.36 ;
      RECT MASK 2 120.127 5.31 120.187 6.36 ;
      RECT MASK 2 120.401 5.31 120.461 6.36 ;
      RECT MASK 2 120.675 5.31 120.735 6.36 ;
      RECT MASK 2 120.949 5.31 121.009 6.36 ;
      RECT MASK 2 121.223 5.31 121.283 6.36 ;
      RECT MASK 2 121.497 5.31 121.557 6.36 ;
      RECT MASK 2 121.771 5.31 121.831 6.36 ;
      RECT MASK 2 122.045 5.31 122.105 6.36 ;
      RECT MASK 2 122.319 5.31 122.379 6.36 ;
      RECT MASK 2 122.593 5.31 122.653 6.36 ;
      RECT MASK 2 122.867 5.31 122.927 6.36 ;
      RECT MASK 2 123.141 5.31 123.201 6.36 ;
      RECT MASK 2 123.415 5.31 123.475 6.36 ;
      RECT MASK 2 123.689 5.31 123.749 6.36 ;
      RECT MASK 2 123.963 5.31 124.023 6.36 ;
      RECT MASK 2 124.237 5.31 124.297 6.36 ;
      RECT MASK 2 124.511 5.31 124.571 6.36 ;
      RECT MASK 2 124.785 5.31 124.845 6.36 ;
      RECT MASK 2 125.059 5.31 125.119 6.36 ;
      RECT MASK 2 125.333 5.31 125.393 6.36 ;
      RECT MASK 2 125.607 5.31 125.667 6.36 ;
      RECT MASK 2 125.881 5.31 125.941 6.36 ;
      RECT MASK 2 126.155 5.31 126.215 6.36 ;
      RECT MASK 2 126.429 5.31 126.489 6.36 ;
      RECT MASK 2 126.703 5.31 126.763 6.36 ;
      RECT MASK 2 126.977 5.31 127.037 6.36 ;
      RECT MASK 2 127.251 5.31 127.311 6.36 ;
      RECT MASK 2 127.525 5.31 127.585 6.36 ;
      RECT MASK 2 127.799 5.31 127.859 6.36 ;
      RECT MASK 2 128.073 5.31 128.133 6.36 ;
      RECT MASK 2 2.2045 5.36 2.4335 5.388 ;
      RECT MASK 2 2.961 5.36 3.28 5.388 ;
      RECT MASK 2 5.251 5.36 5.57 5.388 ;
      RECT MASK 2 8.457 5.36 8.776 5.388 ;
      RECT MASK 2 9.831 5.36 10.0455 5.388 ;
      RECT MASK 2 11.1705 5.36 11.3505 5.388 ;
      RECT MASK 2 11.903 5.36 12.222 5.388 ;
      RECT MASK 2 12.7735 5.36 12.9535 5.388 ;
      RECT MASK 2 14.3195 5.36 14.534 5.388 ;
      RECT MASK 2 21.543 5.36 21.7575 5.388 ;
      RECT MASK 2 25.1795 5.36 25.394 5.388 ;
      RECT MASK 2 32.403 5.36 32.6175 5.388 ;
      RECT MASK 2 33.9835 5.36 34.1635 5.388 ;
      RECT MASK 2 34.715 5.36 35.034 5.388 ;
      RECT MASK 2 35.5865 5.36 35.7665 5.388 ;
      RECT MASK 2 36.8915 5.36 37.106 5.388 ;
      RECT MASK 2 38.161 5.36 38.48 5.388 ;
      RECT MASK 2 41.367 5.36 41.686 5.388 ;
      RECT MASK 2 43.657 5.36 43.976 5.388 ;
      RECT MASK 2 44.5035 5.36 44.7325 5.388 ;
      RECT MASK 2 49.9465 5.37 52.7045 5.43 ;
      RECT MASK 2 53.9045 5.43 56.1725 5.47 ;
      RECT MASK 2 58.4175 5.522 58.621 5.55 ;
      RECT MASK 2 60.343 5.522 60.546 5.55 ;
      RECT MASK 2 50.1675 5.61 50.4465 5.67 ;
      RECT MASK 2 50.8315 5.61 51.1105 5.67 ;
      RECT MASK 2 51.4955 5.61 51.7745 5.67 ;
      RECT MASK 2 52.1595 5.61 52.4385 5.67 ;
      RECT MASK 2 1.6805 5.63 10.7245 5.67 ;
      RECT MASK 2 11.1705 5.63 12.9295 5.67 ;
      RECT MASK 2 13.4005 5.63 21.7575 5.67 ;
      RECT MASK 2 25.1795 5.63 33.5365 5.67 ;
      RECT MASK 2 34.0075 5.63 35.7665 5.67 ;
      RECT MASK 2 36.2125 5.63 45.2565 5.67 ;
      RECT MASK 2 46.7465 5.651 49.0705 5.691 ;
      RECT MASK 2 86.5465 5.698 92.705 5.758 ;
      RECT MASK 2 94 5.698 100.1585 5.758 ;
      RECT MASK 2 58.6465 5.73 58.85 5.758 ;
      RECT MASK 2 59.656 5.73 60.775 5.758 ;
      RECT MASK 2 63.2265 5.73 63.888 5.758 ;
      RECT MASK 2 53.7935 5.771 56.2835 5.811 ;
      RECT MASK 2 1.6805 5.79 10.7245 5.83 ;
      RECT MASK 2 11.1705 5.79 12.9295 5.83 ;
      RECT MASK 2 13.4005 5.79 21.7575 5.83 ;
      RECT MASK 2 25.1795 5.79 33.5365 5.83 ;
      RECT MASK 2 34.0075 5.79 35.7665 5.83 ;
      RECT MASK 2 36.2125 5.79 45.2565 5.83 ;
      RECT MASK 2 46.9055 5.818 47.1235 5.858 ;
      RECT MASK 2 47.2375 5.818 47.4555 5.858 ;
      RECT MASK 2 50.1905 5.85 50.4695 5.91 ;
      RECT MASK 2 50.8545 5.85 51.1335 5.91 ;
      RECT MASK 2 51.5185 5.85 51.7975 5.91 ;
      RECT MASK 2 52.1825 5.85 52.4615 5.91 ;
      RECT MASK 2 58.994 5.878 59.054 6.058 ;
      RECT MASK 2 59.452 5.878 59.512 6.058 ;
      RECT MASK 2 61.055 5.878 61.115 6.058 ;
      RECT MASK 2 61.513 5.878 61.573 6.058 ;
      RECT MASK 2 61.971 5.878 62.031 6.058 ;
      RECT MASK 2 62.429 5.878 62.489 6.058 ;
      RECT MASK 2 62.887 5.878 62.947 6.058 ;
      RECT MASK 2 64.032 5.878 64.092 6.058 ;
      RECT MASK 2 64.49 5.878 64.55 6.058 ;
      RECT MASK 2 64.948 5.878 65.008 6.058 ;
      RECT MASK 2 48.8145 5.9125 48.9945 5.9525 ;
      RECT MASK 2 54.4505 5.938 54.6685 5.978 ;
      RECT MASK 2 55.2805 5.938 55.4985 5.978 ;
      RECT MASK 2 84.1235 5.94 84.461 6 ;
      RECT MASK 2 84.6 5.94 86.293 6 ;
      RECT MASK 2 86.432 5.94 88.125 6 ;
      RECT MASK 2 88.264 5.94 88.583 6 ;
      RECT MASK 2 88.722 5.94 89.041 6 ;
      RECT MASK 2 89.18 5.94 89.499 6 ;
      RECT MASK 2 89.638 5.94 89.957 6 ;
      RECT MASK 2 90.0845 5.94 90.415 6 ;
      RECT MASK 2 90.554 5.94 90.904 6 ;
      RECT MASK 2 91.012 5.94 92.705 6 ;
      RECT MASK 2 94 5.94 95.693 6 ;
      RECT MASK 2 95.801 5.94 96.151 6 ;
      RECT MASK 2 96.29 5.94 96.6205 6 ;
      RECT MASK 2 96.748 5.94 97.067 6 ;
      RECT MASK 2 97.206 5.94 97.525 6 ;
      RECT MASK 2 97.664 5.94 97.983 6 ;
      RECT MASK 2 98.122 5.94 98.441 6 ;
      RECT MASK 2 98.58 5.94 100.273 6 ;
      RECT MASK 2 100.412 5.94 102.105 6 ;
      RECT MASK 2 102.244 5.94 102.5815 6 ;
      RECT MASK 2 60.1675 5.9425 60.3475 5.9825 ;
      RECT MASK 2 65.575 5.9425 65.984 5.9825 ;
      RECT MASK 2 54.8175 5.952 55.0275 6.032 ;
      RECT MASK 2 53.8695 6.0325 54.0495 6.0725 ;
      RECT MASK 2 56.0275 6.0325 56.2075 6.0725 ;
      RECT MASK 2 57.789 6.0625 57.969 6.1025 ;
      RECT MASK 2 2.2045 6.072 2.4335 6.1 ;
      RECT MASK 2 2.961 6.072 3.28 6.1 ;
      RECT MASK 2 5.251 6.072 5.57 6.1 ;
      RECT MASK 2 8.457 6.072 8.776 6.1 ;
      RECT MASK 2 9.831 6.072 10.0455 6.1 ;
      RECT MASK 2 11.1705 6.072 11.3505 6.1 ;
      RECT MASK 2 11.903 6.072 12.222 6.1 ;
      RECT MASK 2 12.7735 6.072 12.9535 6.1 ;
      RECT MASK 2 14.3195 6.072 14.534 6.1 ;
      RECT MASK 2 21.543 6.072 21.7575 6.1 ;
      RECT MASK 2 25.1795 6.072 25.394 6.1 ;
      RECT MASK 2 32.403 6.072 32.6175 6.1 ;
      RECT MASK 2 33.9835 6.072 34.1635 6.1 ;
      RECT MASK 2 34.715 6.072 35.034 6.1 ;
      RECT MASK 2 35.5865 6.072 35.7665 6.1 ;
      RECT MASK 2 36.8915 6.072 37.106 6.1 ;
      RECT MASK 2 38.161 6.072 38.48 6.1 ;
      RECT MASK 2 41.367 6.072 41.686 6.1 ;
      RECT MASK 2 43.657 6.072 43.976 6.1 ;
      RECT MASK 2 44.5035 6.072 44.7325 6.1 ;
      RECT MASK 2 49.9465 6.09 52.7045 6.15 ;
      RECT MASK 2 55.1145 6.197 55.2945 6.237 ;
      RECT MASK 2 2.6325 6.208 2.6925 6.388 ;
      RECT MASK 2 11.5745 6.208 11.6345 6.388 ;
      RECT MASK 2 12.4905 6.208 12.5505 6.388 ;
      RECT MASK 2 14.8025 6.208 14.8625 6.388 ;
      RECT MASK 2 15.2605 6.208 15.3205 6.388 ;
      RECT MASK 2 15.7185 6.208 15.7785 6.388 ;
      RECT MASK 2 16.1765 6.208 16.2365 6.388 ;
      RECT MASK 2 16.6345 6.208 16.6945 6.388 ;
      RECT MASK 2 17.0925 6.208 17.1525 6.388 ;
      RECT MASK 2 17.5505 6.208 17.6105 6.388 ;
      RECT MASK 2 18.0085 6.208 18.0685 6.388 ;
      RECT MASK 2 18.4665 6.208 18.5265 6.388 ;
      RECT MASK 2 18.9245 6.208 18.9845 6.388 ;
      RECT MASK 2 19.3825 6.208 19.4425 6.388 ;
      RECT MASK 2 19.8405 6.208 19.9005 6.388 ;
      RECT MASK 2 20.2985 6.208 20.3585 6.388 ;
      RECT MASK 2 20.7565 6.208 20.8165 6.388 ;
      RECT MASK 2 21.2145 6.208 21.2745 6.388 ;
      RECT MASK 2 25.6625 6.208 25.7225 6.388 ;
      RECT MASK 2 26.1205 6.208 26.1805 6.388 ;
      RECT MASK 2 26.5785 6.208 26.6385 6.388 ;
      RECT MASK 2 27.0365 6.208 27.0965 6.388 ;
      RECT MASK 2 27.4945 6.208 27.5545 6.388 ;
      RECT MASK 2 27.9525 6.208 28.0125 6.388 ;
      RECT MASK 2 28.4105 6.208 28.4705 6.388 ;
      RECT MASK 2 28.8685 6.208 28.9285 6.388 ;
      RECT MASK 2 29.3265 6.208 29.3865 6.388 ;
      RECT MASK 2 29.7845 6.208 29.8445 6.388 ;
      RECT MASK 2 30.2425 6.208 30.3025 6.388 ;
      RECT MASK 2 30.7005 6.208 30.7605 6.388 ;
      RECT MASK 2 31.1585 6.208 31.2185 6.388 ;
      RECT MASK 2 31.6165 6.208 31.6765 6.388 ;
      RECT MASK 2 32.0745 6.208 32.1345 6.388 ;
      RECT MASK 2 34.3865 6.208 34.4465 6.388 ;
      RECT MASK 2 35.3025 6.208 35.3625 6.388 ;
      RECT MASK 2 44.2445 6.208 44.3045 6.388 ;
      RECT MASK 2 22.2135 6.273 23.3235 6.297 ;
      RECT MASK 2 23.6135 6.273 24.7235 6.297 ;
      RECT MASK 2 58.74 6.299 59.766 6.339 ;
      RECT MASK 2 60.9255 6.299 63.0765 6.339 ;
      RECT MASK 2 63.778 6.299 64.9085 6.339 ;
      RECT MASK 2 83.7885 6.32 93.0585 6.36 ;
      RECT MASK 2 93.6465 6.32 102.9165 6.36 ;
      RECT MASK 2 49.9395 6.35 52.6895 6.39 ;
      RECT MASK 2 22.2135 6.363 23.3235 6.387 ;
      RECT MASK 2 23.6135 6.363 24.7235 6.387 ;
      RECT MASK 2 10.3585 6.3925 10.5385 6.4325 ;
      RECT MASK 2 13.5865 6.3925 13.7665 6.4325 ;
      RECT MASK 2 33.1705 6.3925 33.3505 6.4325 ;
      RECT MASK 2 36.3985 6.3925 36.5785 6.4325 ;
      RECT MASK 2 55.1145 6.423 55.2945 6.463 ;
      RECT MASK 2 1.6135 6.4525 1.8575 6.4925 ;
      RECT MASK 2 45.0795 6.4525 45.3235 6.4925 ;
      RECT MASK 2 22.2135 6.453 23.3235 6.477 ;
      RECT MASK 2 23.6135 6.453 24.7235 6.477 ;
      RECT MASK 2 48.8145 6.4675 48.9945 6.5075 ;
      RECT MASK 2 83.7885 6.48 93.0585 6.52 ;
      RECT MASK 2 93.6465 6.48 102.9165 6.52 ;
      RECT MASK 2 58.74 6.501 59.766 6.541 ;
      RECT MASK 2 60.9255 6.501 63.0765 6.541 ;
      RECT MASK 2 63.778 6.501 64.9085 6.541 ;
      RECT MASK 2 49.9395 6.51 52.6895 6.55 ;
      RECT MASK 2 2.3785 6.528 2.8505 6.568 ;
      RECT MASK 2 3.3985 6.528 3.738 6.568 ;
      RECT MASK 2 4.3185 6.528 5.4655 6.568 ;
      RECT MASK 2 5.938 6.528 6.3815 6.568 ;
      RECT MASK 2 6.854 6.528 7.2975 6.568 ;
      RECT MASK 2 7.77 6.528 8.6715 6.568 ;
      RECT MASK 2 8.915 6.528 10.1875 6.568 ;
      RECT MASK 2 36.7495 6.528 38.022 6.568 ;
      RECT MASK 2 38.2655 6.528 39.167 6.568 ;
      RECT MASK 2 39.6395 6.528 40.083 6.568 ;
      RECT MASK 2 40.5555 6.528 40.999 6.568 ;
      RECT MASK 2 41.4715 6.528 42.6185 6.568 ;
      RECT MASK 2 43.199 6.528 43.5385 6.568 ;
      RECT MASK 2 44.0865 6.528 44.5585 6.568 ;
      RECT MASK 2 46.9055 6.562 47.1235 6.602 ;
      RECT MASK 2 47.2375 6.562 47.4555 6.602 ;
      RECT MASK 2 53.8695 6.5875 54.0495 6.6275 ;
      RECT MASK 2 56.0275 6.5875 56.2075 6.6275 ;
      RECT MASK 2 54.8175 6.628 55.1665 6.708 ;
      RECT MASK 2 54.4505 6.682 54.6685 6.722 ;
      RECT MASK 2 55.2805 6.682 55.4985 6.722 ;
      RECT MASK 2 46.7465 6.729 49.0705 6.769 ;
      RECT MASK 2 57.789 6.7375 57.969 6.7775 ;
      RECT MASK 2 60.1675 6.7375 60.3475 6.7775 ;
      RECT MASK 2 65.575 6.7375 65.984 6.7775 ;
      RECT MASK 2 49.9395 6.77 52.6895 6.81 ;
      RECT MASK 2 58.994 6.782 59.054 6.962 ;
      RECT MASK 2 59.452 6.782 59.512 6.962 ;
      RECT MASK 2 61.055 6.782 61.115 6.962 ;
      RECT MASK 2 61.513 6.782 61.573 6.962 ;
      RECT MASK 2 61.971 6.782 62.031 6.962 ;
      RECT MASK 2 62.429 6.782 62.489 6.962 ;
      RECT MASK 2 62.887 6.782 62.947 6.962 ;
      RECT MASK 2 64.032 6.782 64.092 6.962 ;
      RECT MASK 2 64.49 6.782 64.55 6.962 ;
      RECT MASK 2 64.948 6.782 65.008 6.962 ;
      RECT MASK 2 22.3735 6.813 22.7635 6.837 ;
      RECT MASK 2 24.1735 6.813 24.5635 6.837 ;
      RECT MASK 2 53.7935 6.849 56.2835 6.889 ;
      RECT MASK 2 22.2135 6.903 23.3235 6.927 ;
      RECT MASK 2 23.6135 6.903 24.7235 6.927 ;
      RECT MASK 2 49.9395 6.93 52.6895 6.97 ;
      RECT MASK 2 2.3785 6.932 2.8505 6.972 ;
      RECT MASK 2 3.3985 6.932 3.738 6.972 ;
      RECT MASK 2 4.3185 6.932 5.4655 6.972 ;
      RECT MASK 2 5.938 6.932 6.3815 6.972 ;
      RECT MASK 2 6.854 6.932 7.2975 6.972 ;
      RECT MASK 2 7.77 6.932 8.6715 6.972 ;
      RECT MASK 2 12.361 6.932 13.0765 6.972 ;
      RECT MASK 2 33.8605 6.932 34.576 6.972 ;
      RECT MASK 2 38.2655 6.932 39.167 6.972 ;
      RECT MASK 2 39.6395 6.932 40.083 6.972 ;
      RECT MASK 2 40.5555 6.932 40.999 6.972 ;
      RECT MASK 2 41.4715 6.932 42.6185 6.972 ;
      RECT MASK 2 43.199 6.932 43.5385 6.972 ;
      RECT MASK 2 44.0865 6.932 44.5585 6.972 ;
      RECT MASK 2 83.7875 6.98 91.6835 7.02 ;
      RECT MASK 2 95.0215 6.98 102.9175 7.02 ;
      RECT MASK 2 22.4135 6.993 22.7135 7.017 ;
      RECT MASK 2 22.8235 6.993 23.1235 7.017 ;
      RECT MASK 2 23.8135 6.993 24.1135 7.017 ;
      RECT MASK 2 24.2235 6.993 24.5235 7.017 ;
      RECT MASK 2 1.6135 7.0075 1.8575 7.0475 ;
      RECT MASK 2 45.0795 7.0075 45.3235 7.0475 ;
      RECT MASK 2 116.291 7.02 116.351 8.07 ;
      RECT MASK 2 116.565 7.02 116.625 8.07 ;
      RECT MASK 2 116.839 7.02 116.899 8.07 ;
      RECT MASK 2 117.113 7.02 117.173 8.07 ;
      RECT MASK 2 117.387 7.02 117.447 8.07 ;
      RECT MASK 2 117.661 7.02 117.721 8.07 ;
      RECT MASK 2 117.935 7.02 117.995 8.07 ;
      RECT MASK 2 118.209 7.02 118.269 8.07 ;
      RECT MASK 2 118.483 7.02 118.543 8.07 ;
      RECT MASK 2 118.757 7.02 118.817 8.07 ;
      RECT MASK 2 119.031 7.02 119.091 8.07 ;
      RECT MASK 2 119.305 7.02 119.365 8.07 ;
      RECT MASK 2 119.579 7.02 119.639 8.07 ;
      RECT MASK 2 119.853 7.02 119.913 8.07 ;
      RECT MASK 2 120.127 7.02 120.187 8.07 ;
      RECT MASK 2 120.401 7.02 120.461 8.07 ;
      RECT MASK 2 120.675 7.02 120.735 8.07 ;
      RECT MASK 2 120.949 7.02 121.009 8.07 ;
      RECT MASK 2 121.223 7.02 121.283 8.07 ;
      RECT MASK 2 121.497 7.02 121.557 8.07 ;
      RECT MASK 2 121.771 7.02 121.831 8.07 ;
      RECT MASK 2 122.045 7.02 122.105 8.07 ;
      RECT MASK 2 122.319 7.02 122.379 8.07 ;
      RECT MASK 2 122.593 7.02 122.653 8.07 ;
      RECT MASK 2 122.867 7.02 122.927 8.07 ;
      RECT MASK 2 123.141 7.02 123.201 8.07 ;
      RECT MASK 2 123.415 7.02 123.475 8.07 ;
      RECT MASK 2 123.689 7.02 123.749 8.07 ;
      RECT MASK 2 123.963 7.02 124.023 8.07 ;
      RECT MASK 2 124.237 7.02 124.297 8.07 ;
      RECT MASK 2 124.511 7.02 124.571 8.07 ;
      RECT MASK 2 124.785 7.02 124.845 8.07 ;
      RECT MASK 2 125.059 7.02 125.119 8.07 ;
      RECT MASK 2 125.333 7.02 125.393 8.07 ;
      RECT MASK 2 125.607 7.02 125.667 8.07 ;
      RECT MASK 2 125.881 7.02 125.941 8.07 ;
      RECT MASK 2 126.155 7.02 126.215 8.07 ;
      RECT MASK 2 126.429 7.02 126.489 8.07 ;
      RECT MASK 2 126.703 7.02 126.763 8.07 ;
      RECT MASK 2 126.977 7.02 127.037 8.07 ;
      RECT MASK 2 127.251 7.02 127.311 8.07 ;
      RECT MASK 2 127.525 7.02 127.585 8.07 ;
      RECT MASK 2 127.799 7.02 127.859 8.07 ;
      RECT MASK 2 128.073 7.02 128.133 8.07 ;
      RECT MASK 2 10.3585 7.0675 10.5385 7.1075 ;
      RECT MASK 2 13.5865 7.0675 13.7665 7.1075 ;
      RECT MASK 2 33.1705 7.0675 33.3505 7.1075 ;
      RECT MASK 2 36.3985 7.0675 36.5785 7.1075 ;
      RECT MASK 2 58.6465 7.082 58.85 7.11 ;
      RECT MASK 2 59.656 7.082 60.775 7.11 ;
      RECT MASK 2 63.2265 7.082 63.888 7.11 ;
      RECT MASK 2 22.4135 7.083 22.7135 7.107 ;
      RECT MASK 2 22.8235 7.083 23.1235 7.107 ;
      RECT MASK 2 23.8135 7.083 24.1135 7.107 ;
      RECT MASK 2 24.2235 7.083 24.5235 7.107 ;
      RECT MASK 2 46.7465 7.091 49.0705 7.131 ;
      RECT MASK 2 2.6325 7.112 2.6925 7.292 ;
      RECT MASK 2 11.5745 7.112 11.6345 7.292 ;
      RECT MASK 2 12.4905 7.112 12.5505 7.292 ;
      RECT MASK 2 14.8025 7.112 14.8625 7.292 ;
      RECT MASK 2 15.2605 7.112 15.3205 7.292 ;
      RECT MASK 2 15.7185 7.112 15.7785 7.292 ;
      RECT MASK 2 16.1765 7.112 16.2365 7.292 ;
      RECT MASK 2 16.6345 7.112 16.6945 7.292 ;
      RECT MASK 2 17.0925 7.112 17.1525 7.292 ;
      RECT MASK 2 17.5505 7.112 17.6105 7.292 ;
      RECT MASK 2 18.0085 7.112 18.0685 7.292 ;
      RECT MASK 2 18.4665 7.112 18.5265 7.292 ;
      RECT MASK 2 18.9245 7.112 18.9845 7.292 ;
      RECT MASK 2 19.3825 7.112 19.4425 7.292 ;
      RECT MASK 2 19.8405 7.112 19.9005 7.292 ;
      RECT MASK 2 20.2985 7.112 20.3585 7.292 ;
      RECT MASK 2 20.7565 7.112 20.8165 7.292 ;
      RECT MASK 2 21.2145 7.112 21.2745 7.292 ;
      RECT MASK 2 25.6625 7.112 25.7225 7.292 ;
      RECT MASK 2 26.1205 7.112 26.1805 7.292 ;
      RECT MASK 2 26.5785 7.112 26.6385 7.292 ;
      RECT MASK 2 27.0365 7.112 27.0965 7.292 ;
      RECT MASK 2 27.4945 7.112 27.5545 7.292 ;
      RECT MASK 2 27.9525 7.112 28.0125 7.292 ;
      RECT MASK 2 28.4105 7.112 28.4705 7.292 ;
      RECT MASK 2 28.8685 7.112 28.9285 7.292 ;
      RECT MASK 2 29.3265 7.112 29.3865 7.292 ;
      RECT MASK 2 29.7845 7.112 29.8445 7.292 ;
      RECT MASK 2 30.2425 7.112 30.3025 7.292 ;
      RECT MASK 2 30.7005 7.112 30.7605 7.292 ;
      RECT MASK 2 31.1585 7.112 31.2185 7.292 ;
      RECT MASK 2 31.6165 7.112 31.6765 7.292 ;
      RECT MASK 2 32.0745 7.112 32.1345 7.292 ;
      RECT MASK 2 34.3865 7.112 34.4465 7.292 ;
      RECT MASK 2 35.3025 7.112 35.3625 7.292 ;
      RECT MASK 2 44.2445 7.112 44.3045 7.292 ;
      RECT MASK 2 83.7875 7.14 91.6835 7.18 ;
      RECT MASK 2 95.0215 7.14 102.9175 7.18 ;
      RECT MASK 2 22.4135 7.173 22.7135 7.197 ;
      RECT MASK 2 22.8235 7.173 23.1235 7.197 ;
      RECT MASK 2 23.8135 7.173 24.1135 7.197 ;
      RECT MASK 2 24.2235 7.173 24.5235 7.197 ;
      RECT MASK 2 53.9045 7.19 56.1725 7.23 ;
      RECT MASK 2 46.9055 7.258 47.1235 7.298 ;
      RECT MASK 2 47.2375 7.258 47.4555 7.298 ;
      RECT MASK 2 47.5695 7.258 47.7875 7.298 ;
      RECT MASK 2 47.9365 7.258 48.2855 7.298 ;
      RECT MASK 2 49.9465 7.29 52.6825 7.35 ;
      RECT MASK 2 58.6465 7.29 58.85 7.318 ;
      RECT MASK 2 59.656 7.29 60.775 7.318 ;
      RECT MASK 2 63.2265 7.29 63.888 7.318 ;
      RECT MASK 2 53.9045 7.35 56.1725 7.39 ;
      RECT MASK 2 48.8145 7.3525 48.9945 7.3925 ;
      RECT MASK 2 2.2045 7.4 2.4335 7.428 ;
      RECT MASK 2 2.961 7.4 3.28 7.428 ;
      RECT MASK 2 5.251 7.4 5.57 7.428 ;
      RECT MASK 2 8.457 7.4 8.776 7.428 ;
      RECT MASK 2 9.831 7.4 10.0455 7.428 ;
      RECT MASK 2 11.1705 7.4 11.3505 7.428 ;
      RECT MASK 2 11.903 7.4 12.222 7.428 ;
      RECT MASK 2 12.7735 7.4 12.9535 7.428 ;
      RECT MASK 2 14.3195 7.4 14.534 7.428 ;
      RECT MASK 2 21.543 7.4 21.7575 7.428 ;
      RECT MASK 2 25.1795 7.4 25.394 7.428 ;
      RECT MASK 2 32.403 7.4 32.6175 7.428 ;
      RECT MASK 2 33.9835 7.4 34.1635 7.428 ;
      RECT MASK 2 34.715 7.4 35.034 7.428 ;
      RECT MASK 2 35.5865 7.4 35.7665 7.428 ;
      RECT MASK 2 36.8915 7.4 37.106 7.428 ;
      RECT MASK 2 38.161 7.4 38.48 7.428 ;
      RECT MASK 2 41.367 7.4 41.686 7.428 ;
      RECT MASK 2 43.657 7.4 43.976 7.428 ;
      RECT MASK 2 44.5035 7.4 44.7325 7.428 ;
      RECT MASK 2 48.0675 7.425 48.2475 7.465 ;
      RECT MASK 2 58.994 7.438 59.054 7.618 ;
      RECT MASK 2 59.452 7.438 59.512 7.618 ;
      RECT MASK 2 61.055 7.438 61.115 7.618 ;
      RECT MASK 2 61.513 7.438 61.573 7.618 ;
      RECT MASK 2 61.971 7.438 62.031 7.618 ;
      RECT MASK 2 62.429 7.438 62.489 7.618 ;
      RECT MASK 2 62.887 7.438 62.947 7.618 ;
      RECT MASK 2 64.032 7.438 64.092 7.618 ;
      RECT MASK 2 64.49 7.438 64.55 7.618 ;
      RECT MASK 2 64.948 7.438 65.008 7.618 ;
      RECT MASK 2 22.2235 7.518 23.3135 7.542 ;
      RECT MASK 2 23.6235 7.518 24.7135 7.542 ;
      RECT MASK 2 50.1075 7.53 50.2875 7.59 ;
      RECT MASK 2 50.7715 7.53 50.9515 7.59 ;
      RECT MASK 2 51.4355 7.53 51.6155 7.59 ;
      RECT MASK 2 52.0995 7.53 52.2795 7.59 ;
      RECT MASK 2 57.789 7.6225 57.969 7.6625 ;
      RECT MASK 2 60.1675 7.6225 60.3475 7.6625 ;
      RECT MASK 2 65.575 7.6225 65.984 7.6625 ;
      RECT MASK 2 84.406 7.651 88.312 7.711 ;
      RECT MASK 2 88.5295 7.651 88.9265 7.711 ;
      RECT MASK 2 89.158 7.651 89.6485 7.711 ;
      RECT MASK 2 90.1785 7.651 90.4035 7.711 ;
      RECT MASK 2 90.6685 7.651 91.065 7.711 ;
      RECT MASK 2 95.64 7.651 96.0365 7.711 ;
      RECT MASK 2 96.3015 7.651 96.5265 7.711 ;
      RECT MASK 2 97.0565 7.651 97.547 7.711 ;
      RECT MASK 2 97.7785 7.651 98.1755 7.711 ;
      RECT MASK 2 98.393 7.651 102.299 7.711 ;
      RECT MASK 2 1.6805 7.67 13.9525 7.71 ;
      RECT MASK 2 14.3195 7.67 21.7575 7.71 ;
      RECT MASK 2 25.1795 7.67 32.6175 7.71 ;
      RECT MASK 2 32.9845 7.67 45.2565 7.71 ;
      RECT MASK 2 49.9465 7.77 52.6825 7.83 ;
      RECT MASK 2 1.6805 7.83 13.9525 7.87 ;
      RECT MASK 2 14.3195 7.83 21.7575 7.87 ;
      RECT MASK 2 25.1795 7.83 32.6175 7.87 ;
      RECT MASK 2 32.9845 7.83 45.2565 7.87 ;
      RECT MASK 2 48.0675 7.835 48.2475 7.875 ;
      RECT MASK 2 58.74 7.859 59.766 7.899 ;
      RECT MASK 2 60.9255 7.859 63.0765 7.899 ;
      RECT MASK 2 63.778 7.859 64.9085 7.899 ;
      RECT MASK 2 48.8145 7.9075 48.9945 7.9475 ;
      RECT MASK 2 73.8505 7.999 74.2885 8.179 ;
      RECT MASK 2 74.6165 7.999 75.1445 8.179 ;
      RECT MASK 2 75.4725 7.999 75.9105 8.179 ;
      RECT MASK 2 110.7945 7.999 111.2325 8.179 ;
      RECT MASK 2 111.5605 7.999 112.0885 8.179 ;
      RECT MASK 2 112.4165 7.999 112.8545 8.179 ;
      RECT MASK 2 46.9055 8.002 47.1235 8.042 ;
      RECT MASK 2 47.2375 8.002 47.4555 8.042 ;
      RECT MASK 2 47.5695 8.002 47.7875 8.042 ;
      RECT MASK 2 47.9365 8.002 48.1465 8.042 ;
      RECT MASK 2 50.3495 8.01 50.5295 8.07 ;
      RECT MASK 2 51.0135 8.01 51.1935 8.07 ;
      RECT MASK 2 51.6775 8.01 51.8575 8.07 ;
      RECT MASK 2 52.3415 8.01 52.5215 8.07 ;
      RECT MASK 2 58.74 8.061 59.766 8.101 ;
      RECT MASK 2 60.9255 8.061 63.0765 8.101 ;
      RECT MASK 2 63.778 8.061 64.9085 8.101 ;
      RECT MASK 2 1.6805 8.09 13.9525 8.13 ;
      RECT MASK 2 14.3195 8.09 21.7575 8.13 ;
      RECT MASK 2 46.7465 8.169 49.0705 8.209 ;
      RECT MASK 2 83.7875 8.24 91.6755 8.28 ;
      RECT MASK 2 95.0295 8.24 102.9175 8.28 ;
      RECT MASK 2 1.6805 8.25 13.9525 8.29 ;
      RECT MASK 2 14.3195 8.25 21.7575 8.29 ;
      RECT MASK 2 50.1525 8.25 50.4695 8.31 ;
      RECT MASK 2 50.8165 8.25 51.1335 8.31 ;
      RECT MASK 2 51.4805 8.25 51.7975 8.31 ;
      RECT MASK 2 52.1445 8.25 52.4615 8.31 ;
      RECT MASK 2 57.789 8.2975 57.969 8.3375 ;
      RECT MASK 2 58.994 8.342 59.054 8.522 ;
      RECT MASK 2 59.452 8.342 59.512 8.522 ;
      RECT MASK 2 61.055 8.342 61.115 8.522 ;
      RECT MASK 2 61.513 8.342 61.573 8.522 ;
      RECT MASK 2 61.971 8.342 62.031 8.522 ;
      RECT MASK 2 62.429 8.342 62.489 8.522 ;
      RECT MASK 2 62.887 8.342 62.947 8.522 ;
      RECT MASK 2 64.032 8.342 64.092 8.522 ;
      RECT MASK 2 64.49 8.342 64.55 8.522 ;
      RECT MASK 2 64.948 8.342 65.008 8.522 ;
      RECT MASK 2 83.7875 8.4 91.6835 8.44 ;
      RECT MASK 2 95.0215 8.4 102.9175 8.44 ;
      RECT MASK 2 60.1675 8.4175 60.3475 8.4575 ;
      RECT MASK 2 65.575 8.4175 65.984 8.4575 ;
      RECT MASK 2 22.2235 8.418 23.3135 8.442 ;
      RECT MASK 2 50.1675 8.49 50.4465 8.55 ;
      RECT MASK 2 50.8315 8.49 51.1105 8.55 ;
      RECT MASK 2 51.4955 8.49 51.7745 8.55 ;
      RECT MASK 2 52.1595 8.49 52.4385 8.55 ;
      RECT MASK 2 67.634 8.51 70.721 8.55 ;
      RECT MASK 2 46.7465 8.531 49.0705 8.571 ;
      RECT MASK 2 2.2045 8.532 2.4335 8.56 ;
      RECT MASK 2 2.961 8.532 3.28 8.56 ;
      RECT MASK 2 5.251 8.532 5.57 8.56 ;
      RECT MASK 2 8.457 8.532 8.776 8.56 ;
      RECT MASK 2 9.831 8.532 10.0455 8.56 ;
      RECT MASK 2 11.1705 8.532 11.3505 8.56 ;
      RECT MASK 2 11.903 8.532 12.222 8.56 ;
      RECT MASK 2 12.7735 8.532 12.9535 8.56 ;
      RECT MASK 2 14.3195 8.532 14.534 8.56 ;
      RECT MASK 2 21.543 8.532 21.7575 8.56 ;
      RECT MASK 2 31.5485 8.54 39.1995 8.58 ;
      RECT MASK 2 53.7665 8.54 56.1665 8.58 ;
      RECT MASK 2 72.7245 8.6 76.9845 8.64 ;
      RECT MASK 2 109.7205 8.6 113.9805 8.64 ;
      RECT MASK 2 58.6465 8.642 58.85 8.67 ;
      RECT MASK 2 59.656 8.642 60.775 8.67 ;
      RECT MASK 2 63.2265 8.642 63.888 8.67 ;
      RECT MASK 2 2.6325 8.668 2.6925 8.848 ;
      RECT MASK 2 11.5745 8.668 11.6345 8.848 ;
      RECT MASK 2 12.4905 8.668 12.5505 8.848 ;
      RECT MASK 2 14.8025 8.668 14.8625 8.848 ;
      RECT MASK 2 15.2605 8.668 15.3205 8.848 ;
      RECT MASK 2 15.7185 8.668 15.7785 8.848 ;
      RECT MASK 2 16.1765 8.668 16.2365 8.848 ;
      RECT MASK 2 16.6345 8.668 16.6945 8.848 ;
      RECT MASK 2 17.0925 8.668 17.1525 8.848 ;
      RECT MASK 2 17.5505 8.668 17.6105 8.848 ;
      RECT MASK 2 18.0085 8.668 18.0685 8.848 ;
      RECT MASK 2 18.4665 8.668 18.5265 8.848 ;
      RECT MASK 2 18.9245 8.668 18.9845 8.848 ;
      RECT MASK 2 19.3825 8.668 19.4425 8.848 ;
      RECT MASK 2 19.8405 8.668 19.9005 8.848 ;
      RECT MASK 2 20.2985 8.668 20.3585 8.848 ;
      RECT MASK 2 20.7565 8.668 20.8165 8.848 ;
      RECT MASK 2 21.2145 8.668 21.2745 8.848 ;
      RECT MASK 2 67.634 8.67 70.721 8.71 ;
      RECT MASK 2 46.9055 8.698 47.1235 8.738 ;
      RECT MASK 2 47.2375 8.698 47.4555 8.738 ;
      RECT MASK 2 47.6045 8.698 47.8145 8.738 ;
      RECT MASK 2 48.0675 8.698 48.2855 8.738 ;
      RECT MASK 2 31.5485 8.7 39.1995 8.74 ;
      RECT MASK 2 53.7665 8.7 56.1665 8.74 ;
      RECT MASK 2 116.291 8.73 116.351 9.78 ;
      RECT MASK 2 116.565 8.73 116.625 9.78 ;
      RECT MASK 2 116.839 8.73 116.899 9.78 ;
      RECT MASK 2 117.113 8.73 117.173 9.78 ;
      RECT MASK 2 117.387 8.73 117.447 9.78 ;
      RECT MASK 2 117.661 8.73 117.721 9.78 ;
      RECT MASK 2 117.935 8.73 117.995 9.78 ;
      RECT MASK 2 118.209 8.73 118.269 9.78 ;
      RECT MASK 2 118.483 8.73 118.543 9.78 ;
      RECT MASK 2 118.757 8.73 118.817 9.78 ;
      RECT MASK 2 119.031 8.73 119.091 9.78 ;
      RECT MASK 2 119.305 8.73 119.365 9.78 ;
      RECT MASK 2 119.579 8.73 119.639 9.78 ;
      RECT MASK 2 119.853 8.73 119.913 9.78 ;
      RECT MASK 2 120.127 8.73 120.187 9.78 ;
      RECT MASK 2 120.401 8.73 120.461 9.78 ;
      RECT MASK 2 120.675 8.73 120.735 9.78 ;
      RECT MASK 2 120.949 8.73 121.009 9.78 ;
      RECT MASK 2 121.223 8.73 121.283 9.78 ;
      RECT MASK 2 121.497 8.73 121.557 9.78 ;
      RECT MASK 2 121.771 8.73 121.831 9.78 ;
      RECT MASK 2 122.045 8.73 122.105 9.78 ;
      RECT MASK 2 122.319 8.73 122.379 9.78 ;
      RECT MASK 2 122.593 8.73 122.653 9.78 ;
      RECT MASK 2 122.867 8.73 122.927 9.78 ;
      RECT MASK 2 123.141 8.73 123.201 9.78 ;
      RECT MASK 2 123.415 8.73 123.475 9.78 ;
      RECT MASK 2 123.689 8.73 123.749 9.78 ;
      RECT MASK 2 123.963 8.73 124.023 9.78 ;
      RECT MASK 2 124.237 8.73 124.297 9.78 ;
      RECT MASK 2 124.511 8.73 124.571 9.78 ;
      RECT MASK 2 124.785 8.73 124.845 9.78 ;
      RECT MASK 2 125.059 8.73 125.119 9.78 ;
      RECT MASK 2 125.333 8.73 125.393 9.78 ;
      RECT MASK 2 125.607 8.73 125.667 9.78 ;
      RECT MASK 2 125.881 8.73 125.941 9.78 ;
      RECT MASK 2 126.155 8.73 126.215 9.78 ;
      RECT MASK 2 126.429 8.73 126.489 9.78 ;
      RECT MASK 2 126.703 8.73 126.763 9.78 ;
      RECT MASK 2 126.977 8.73 127.037 9.78 ;
      RECT MASK 2 127.251 8.73 127.311 9.78 ;
      RECT MASK 2 127.525 8.73 127.585 9.78 ;
      RECT MASK 2 127.799 8.73 127.859 9.78 ;
      RECT MASK 2 128.073 8.73 128.133 9.78 ;
      RECT MASK 2 72.7245 8.76 76.9845 8.8 ;
      RECT MASK 2 109.7205 8.76 113.9805 8.8 ;
      RECT MASK 2 22.4135 8.763 22.7135 8.787 ;
      RECT MASK 2 22.8235 8.763 23.1235 8.787 ;
      RECT MASK 2 48.8145 8.7925 48.9945 8.8325 ;
      RECT MASK 2 58.4175 8.85 58.621 8.878 ;
      RECT MASK 2 60.343 8.85 60.546 8.878 ;
      RECT MASK 2 10.3585 8.8525 10.5385 8.8925 ;
      RECT MASK 2 13.5865 8.8525 13.7665 8.8925 ;
      RECT MASK 2 22.4135 8.853 22.7135 8.877 ;
      RECT MASK 2 22.8235 8.853 23.1235 8.877 ;
      RECT MASK 2 47.7355 8.865 47.9155 8.905 ;
      RECT MASK 2 49.9395 8.9 52.6895 8.94 ;
      RECT MASK 2 1.6135 8.9125 1.8575 8.9525 ;
      RECT MASK 2 22.4135 8.943 22.7135 8.967 ;
      RECT MASK 2 22.8235 8.943 23.1235 8.967 ;
      RECT MASK 2 2.3785 8.988 2.8505 9.028 ;
      RECT MASK 2 3.3985 8.988 3.738 9.028 ;
      RECT MASK 2 4.3185 8.988 5.4655 9.028 ;
      RECT MASK 2 5.938 8.988 6.3815 9.028 ;
      RECT MASK 2 6.854 8.988 7.2975 9.028 ;
      RECT MASK 2 7.77 8.988 8.6715 9.028 ;
      RECT MASK 2 12.361 8.988 13.0765 9.028 ;
      RECT MASK 2 58.765 8.998 58.825 9.178 ;
      RECT MASK 2 59.223 8.998 59.283 9.178 ;
      RECT MASK 2 59.681 8.998 59.741 9.178 ;
      RECT MASK 2 60.139 8.998 60.199 9.178 ;
      RECT MASK 2 62.658 8.998 62.718 9.178 ;
      RECT MASK 2 63.116 8.998 63.176 9.178 ;
      RECT MASK 2 63.574 8.998 63.634 9.178 ;
      RECT MASK 2 64.032 8.998 64.092 9.178 ;
      RECT MASK 2 64.49 8.998 64.55 9.178 ;
      RECT MASK 2 64.948 8.998 65.008 9.178 ;
      RECT MASK 2 65.406 8.998 65.466 9.178 ;
      RECT MASK 2 65.864 8.998 65.924 9.178 ;
      RECT MASK 2 22.2135 9.033 23.3235 9.057 ;
      RECT MASK 2 32.0535 9.041 38.6945 9.081 ;
      RECT MASK 2 49.9395 9.06 52.6895 9.1 ;
      RECT MASK 2 60.995 9.0625 61.404 9.1025 ;
      RECT MASK 2 61.911 9.0625 62.091 9.1025 ;
      RECT MASK 2 22.3735 9.123 22.7635 9.147 ;
      RECT MASK 2 57.789 9.1825 57.969 9.2225 ;
      RECT MASK 2 32.342 9.222 32.7855 9.302 ;
      RECT MASK 2 33.258 9.222 33.7015 9.302 ;
      RECT MASK 2 34.174 9.222 34.6175 9.302 ;
      RECT MASK 2 35.09 9.222 35.5335 9.302 ;
      RECT MASK 2 36.006 9.222 36.4495 9.302 ;
      RECT MASK 2 36.922 9.222 37.3655 9.302 ;
      RECT MASK 2 37.838 9.222 38.2815 9.302 ;
      RECT MASK 2 67.567 9.2725 67.811 9.3125 ;
      RECT MASK 2 70.544 9.2725 70.788 9.3125 ;
      RECT MASK 2 47.7355 9.275 47.9155 9.315 ;
      RECT MASK 2 31.4735 9.3025 31.7175 9.3425 ;
      RECT MASK 2 39.0305 9.3025 39.2745 9.3425 ;
      RECT MASK 2 53.6995 9.3025 53.9435 9.3425 ;
      RECT MASK 2 55.9895 9.3025 56.2335 9.3425 ;
      RECT MASK 2 49.9395 9.32 52.6895 9.36 ;
      RECT MASK 2 48.8145 9.3475 48.9945 9.3875 ;
      RECT MASK 2 2.3785 9.392 2.8505 9.432 ;
      RECT MASK 2 3.3985 9.392 3.738 9.432 ;
      RECT MASK 2 4.3185 9.392 5.4655 9.432 ;
      RECT MASK 2 5.938 9.392 6.3815 9.432 ;
      RECT MASK 2 6.854 9.392 7.2975 9.432 ;
      RECT MASK 2 7.77 9.392 8.6715 9.432 ;
      RECT MASK 2 8.915 9.392 10.1875 9.432 ;
      RECT MASK 2 68.454 9.417 68.514 9.723 ;
      RECT MASK 2 68.696 9.417 68.756 9.723 ;
      RECT MASK 2 68.912 9.417 68.972 9.723 ;
      RECT MASK 2 69.154 9.417 69.214 9.723 ;
      RECT MASK 2 69.599 9.417 69.659 9.723 ;
      RECT MASK 2 69.841 9.417 69.901 9.723 ;
      RECT MASK 2 58.6355 9.419 59.4225 9.459 ;
      RECT MASK 2 59.5415 9.419 60.3285 9.459 ;
      RECT MASK 2 62.862 9.419 64.4505 9.459 ;
      RECT MASK 2 64.5795 9.419 64.9085 9.459 ;
      RECT MASK 2 46.9055 9.442 47.1235 9.482 ;
      RECT MASK 2 47.2375 9.442 47.4555 9.482 ;
      RECT MASK 2 47.6045 9.442 47.9535 9.482 ;
      RECT MASK 2 48.0675 9.442 48.2855 9.482 ;
      RECT MASK 2 54.5865 9.447 54.6465 9.753 ;
      RECT MASK 2 54.8285 9.447 54.8885 9.753 ;
      RECT MASK 2 55.0445 9.447 55.1045 9.753 ;
      RECT MASK 2 55.2865 9.447 55.3465 9.753 ;
      RECT MASK 2 32.7405 9.467 32.945 9.507 ;
      RECT MASK 2 33.6565 9.467 33.861 9.507 ;
      RECT MASK 2 34.5725 9.467 34.777 9.507 ;
      RECT MASK 2 35.4885 9.467 35.693 9.507 ;
      RECT MASK 2 36.4045 9.467 36.609 9.507 ;
      RECT MASK 2 37.3205 9.467 37.525 9.507 ;
      RECT MASK 2 38.2365 9.467 38.441 9.507 ;
      RECT MASK 2 1.6135 9.4675 1.8575 9.5075 ;
      RECT MASK 2 49.9395 9.48 52.6895 9.52 ;
      RECT MASK 2 22.2135 9.483 23.3235 9.507 ;
      RECT MASK 2 10.3585 9.5275 10.5385 9.5675 ;
      RECT MASK 2 13.5865 9.5275 13.7665 9.5675 ;
      RECT MASK 2 2.6325 9.572 2.6925 9.752 ;
      RECT MASK 2 11.5745 9.572 11.6345 9.752 ;
      RECT MASK 2 12.4905 9.572 12.5505 9.752 ;
      RECT MASK 2 14.8025 9.572 14.8625 9.752 ;
      RECT MASK 2 15.2605 9.572 15.3205 9.752 ;
      RECT MASK 2 15.7185 9.572 15.7785 9.752 ;
      RECT MASK 2 16.1765 9.572 16.2365 9.752 ;
      RECT MASK 2 16.6345 9.572 16.6945 9.752 ;
      RECT MASK 2 17.0925 9.572 17.1525 9.752 ;
      RECT MASK 2 17.5505 9.572 17.6105 9.752 ;
      RECT MASK 2 18.0085 9.572 18.0685 9.752 ;
      RECT MASK 2 18.4665 9.572 18.5265 9.752 ;
      RECT MASK 2 18.9245 9.572 18.9845 9.752 ;
      RECT MASK 2 19.3825 9.572 19.4425 9.752 ;
      RECT MASK 2 19.8405 9.572 19.9005 9.752 ;
      RECT MASK 2 20.2985 9.572 20.3585 9.752 ;
      RECT MASK 2 20.7565 9.572 20.8165 9.752 ;
      RECT MASK 2 21.2145 9.572 21.2745 9.752 ;
      RECT MASK 2 22.2135 9.573 23.3235 9.597 ;
      RECT MASK 2 46.7465 9.609 49.0705 9.649 ;
      RECT MASK 2 58.4065 9.621 58.9545 9.661 ;
      RECT MASK 2 59.0935 9.621 59.4225 9.661 ;
      RECT MASK 2 59.5415 9.621 59.8705 9.661 ;
      RECT MASK 2 60.0095 9.621 60.5575 9.661 ;
      RECT MASK 2 62.862 9.621 63.557 9.661 ;
      RECT MASK 2 63.6735 9.621 64.473 9.661 ;
      RECT MASK 2 64.8185 9.621 65.491 9.661 ;
      RECT MASK 2 22.2135 9.663 23.3235 9.687 ;
      RECT MASK 2 32.7405 9.693 32.945 9.733 ;
      RECT MASK 2 33.6565 9.693 33.861 9.733 ;
      RECT MASK 2 34.5725 9.693 34.777 9.733 ;
      RECT MASK 2 35.4885 9.693 35.693 9.733 ;
      RECT MASK 2 36.4045 9.693 36.609 9.733 ;
      RECT MASK 2 37.3205 9.693 37.525 9.733 ;
      RECT MASK 2 38.2365 9.693 38.441 9.733 ;
      RECT MASK 2 78.5035 9.749 78.9415 9.929 ;
      RECT MASK 2 79.2695 9.749 79.7575 9.929 ;
      RECT MASK 2 80.0855 9.749 80.5535 9.929 ;
      RECT MASK 2 80.8815 9.749 81.3195 9.929 ;
      RECT MASK 2 105.3855 9.749 105.8235 9.929 ;
      RECT MASK 2 106.1515 9.749 106.6195 9.929 ;
      RECT MASK 2 106.9475 9.749 107.4355 9.929 ;
      RECT MASK 2 107.7635 9.749 108.2015 9.929 ;
      RECT MASK 2 67.567 9.8275 67.811 9.8675 ;
      RECT MASK 2 70.544 9.8275 70.788 9.8675 ;
      RECT MASK 2 31.4735 9.8575 31.7175 9.8975 ;
      RECT MASK 2 39.0305 9.8575 39.2745 9.8975 ;
      RECT MASK 2 53.6995 9.8575 53.9435 9.8975 ;
      RECT MASK 2 55.9895 9.8575 56.2335 9.8975 ;
      RECT MASK 2 57.789 9.8575 57.969 9.8975 ;
      RECT MASK 2 60.995 9.8575 61.404 9.8975 ;
      RECT MASK 2 61.911 9.8575 62.091 9.8975 ;
      RECT MASK 2 2.2045 9.86 2.4335 9.888 ;
      RECT MASK 2 2.961 9.86 3.28 9.888 ;
      RECT MASK 2 5.251 9.86 5.57 9.888 ;
      RECT MASK 2 8.457 9.86 8.776 9.888 ;
      RECT MASK 2 9.831 9.86 10.0455 9.888 ;
      RECT MASK 2 11.1705 9.86 11.3505 9.888 ;
      RECT MASK 2 11.903 9.86 12.222 9.888 ;
      RECT MASK 2 12.7735 9.86 12.9535 9.888 ;
      RECT MASK 2 14.3195 9.86 14.534 9.888 ;
      RECT MASK 2 21.543 9.86 21.7575 9.888 ;
      RECT MASK 2 32.342 9.9 32.5565 9.98 ;
      RECT MASK 2 33.258 9.9 33.4725 9.98 ;
      RECT MASK 2 34.174 9.9 34.3885 9.98 ;
      RECT MASK 2 35.09 9.9 35.3045 9.98 ;
      RECT MASK 2 36.006 9.9 36.2205 9.98 ;
      RECT MASK 2 36.922 9.9 37.1365 9.98 ;
      RECT MASK 2 37.838 9.9 38.0525 9.98 ;
      RECT MASK 2 58.765 9.902 58.825 10.082 ;
      RECT MASK 2 59.223 9.902 59.283 10.082 ;
      RECT MASK 2 59.681 9.902 59.741 10.082 ;
      RECT MASK 2 60.139 9.902 60.199 10.082 ;
      RECT MASK 2 62.658 9.902 62.718 10.082 ;
      RECT MASK 2 63.116 9.902 63.176 10.082 ;
      RECT MASK 2 63.574 9.902 63.634 10.082 ;
      RECT MASK 2 64.032 9.902 64.092 10.082 ;
      RECT MASK 2 64.49 9.902 64.55 10.082 ;
      RECT MASK 2 64.948 9.902 65.008 10.082 ;
      RECT MASK 2 65.406 9.902 65.466 10.082 ;
      RECT MASK 2 65.864 9.902 65.924 10.082 ;
      RECT MASK 2 46.7745 9.95 48.9595 9.99 ;
      RECT MASK 2 49.9415 10.05 52.6875 10.11 ;
      RECT MASK 2 46.7745 10.11 48.9595 10.15 ;
      RECT MASK 2 32.0535 10.119 38.6945 10.159 ;
      RECT MASK 2 1.6805 10.13 10.7245 10.17 ;
      RECT MASK 2 11.1705 10.13 12.9295 10.17 ;
      RECT MASK 2 13.4005 10.13 21.7575 10.17 ;
      RECT MASK 2 1.6805 10.29 10.7245 10.33 ;
      RECT MASK 2 11.1705 10.29 12.9295 10.33 ;
      RECT MASK 2 13.4005 10.29 21.7575 10.33 ;
      RECT MASK 2 50.1675 10.29 50.4465 10.35 ;
      RECT MASK 2 50.8315 10.29 51.1105 10.35 ;
      RECT MASK 2 51.4955 10.29 51.7745 10.35 ;
      RECT MASK 2 52.1595 10.29 52.4385 10.35 ;
      RECT MASK 2 52.5905 10.29 52.7705 10.35 ;
      RECT MASK 2 77.4385 10.31 82.3625 10.35 ;
      RECT MASK 2 104.3425 10.31 109.2665 10.35 ;
      RECT MASK 2 67.634 10.43 70.721 10.47 ;
      RECT MASK 2 116.291 10.44 116.351 11.49 ;
      RECT MASK 2 116.565 10.44 116.625 11.49 ;
      RECT MASK 2 116.839 10.44 116.899 11.49 ;
      RECT MASK 2 117.113 10.44 117.173 11.49 ;
      RECT MASK 2 117.387 10.44 117.447 11.49 ;
      RECT MASK 2 117.661 10.44 117.721 11.49 ;
      RECT MASK 2 117.935 10.44 117.995 11.49 ;
      RECT MASK 2 118.209 10.44 118.269 11.49 ;
      RECT MASK 2 118.483 10.44 118.543 11.49 ;
      RECT MASK 2 118.757 10.44 118.817 11.49 ;
      RECT MASK 2 119.031 10.44 119.091 11.49 ;
      RECT MASK 2 119.305 10.44 119.365 11.49 ;
      RECT MASK 2 119.579 10.44 119.639 11.49 ;
      RECT MASK 2 119.853 10.44 119.913 11.49 ;
      RECT MASK 2 120.127 10.44 120.187 11.49 ;
      RECT MASK 2 120.401 10.44 120.461 11.49 ;
      RECT MASK 2 120.675 10.44 120.735 11.49 ;
      RECT MASK 2 120.949 10.44 121.009 11.49 ;
      RECT MASK 2 121.223 10.44 121.283 11.49 ;
      RECT MASK 2 121.497 10.44 121.557 11.49 ;
      RECT MASK 2 121.771 10.44 121.831 11.49 ;
      RECT MASK 2 122.045 10.44 122.105 11.49 ;
      RECT MASK 2 122.319 10.44 122.379 11.49 ;
      RECT MASK 2 122.593 10.44 122.653 11.49 ;
      RECT MASK 2 122.867 10.44 122.927 11.49 ;
      RECT MASK 2 123.141 10.44 123.201 11.49 ;
      RECT MASK 2 123.415 10.44 123.475 11.49 ;
      RECT MASK 2 123.689 10.44 123.749 11.49 ;
      RECT MASK 2 123.963 10.44 124.023 11.49 ;
      RECT MASK 2 124.237 10.44 124.297 11.49 ;
      RECT MASK 2 124.511 10.44 124.571 11.49 ;
      RECT MASK 2 124.785 10.44 124.845 11.49 ;
      RECT MASK 2 125.059 10.44 125.119 11.49 ;
      RECT MASK 2 125.333 10.44 125.393 11.49 ;
      RECT MASK 2 125.607 10.44 125.667 11.49 ;
      RECT MASK 2 125.881 10.44 125.941 11.49 ;
      RECT MASK 2 126.155 10.44 126.215 11.49 ;
      RECT MASK 2 126.429 10.44 126.489 11.49 ;
      RECT MASK 2 126.703 10.44 126.763 11.49 ;
      RECT MASK 2 126.977 10.44 127.037 11.49 ;
      RECT MASK 2 127.251 10.44 127.311 11.49 ;
      RECT MASK 2 127.525 10.44 127.585 11.49 ;
      RECT MASK 2 127.799 10.44 127.859 11.49 ;
      RECT MASK 2 128.073 10.44 128.133 11.49 ;
      RECT MASK 2 31.5485 10.46 39.1995 10.5 ;
      RECT MASK 2 53.7665 10.46 56.1665 10.5 ;
      RECT MASK 2 57.824 10.46 60.453 10.5 ;
      RECT MASK 2 61.946 10.46 65.984 10.5 ;
      RECT MASK 2 77.4385 10.47 82.3625 10.51 ;
      RECT MASK 2 104.3425 10.47 109.2665 10.51 ;
      RECT MASK 2 49.9395 10.55 52.6895 10.59 ;
      RECT MASK 2 67.634 10.59 70.721 10.63 ;
      RECT MASK 2 31.5485 10.62 39.1995 10.66 ;
      RECT MASK 2 53.7665 10.62 56.1665 10.66 ;
      RECT MASK 2 57.824 10.62 60.453 10.66 ;
      RECT MASK 2 61.946 10.62 65.984 10.66 ;
      RECT MASK 2 49.9395 10.71 52.6895 10.75 ;
      RECT MASK 2 4.362 11.78 111.8065 11.82 ;
      RECT MASK 2 4.362 11.94 111.8085 11.98 ;
      RECT MASK 2 116.291 12.15 116.351 13.2 ;
      RECT MASK 2 116.565 12.15 116.625 13.2 ;
      RECT MASK 2 116.839 12.15 116.899 13.2 ;
      RECT MASK 2 117.113 12.15 117.173 13.2 ;
      RECT MASK 2 117.387 12.15 117.447 13.2 ;
      RECT MASK 2 117.661 12.15 117.721 13.2 ;
      RECT MASK 2 117.935 12.15 117.995 13.2 ;
      RECT MASK 2 118.209 12.15 118.269 13.2 ;
      RECT MASK 2 118.483 12.15 118.543 13.2 ;
      RECT MASK 2 118.757 12.15 118.817 13.2 ;
      RECT MASK 2 119.031 12.15 119.091 13.2 ;
      RECT MASK 2 119.305 12.15 119.365 13.2 ;
      RECT MASK 2 119.579 12.15 119.639 13.2 ;
      RECT MASK 2 119.853 12.15 119.913 13.2 ;
      RECT MASK 2 120.127 12.15 120.187 13.2 ;
      RECT MASK 2 120.401 12.15 120.461 13.2 ;
      RECT MASK 2 120.675 12.15 120.735 13.2 ;
      RECT MASK 2 120.949 12.15 121.009 13.2 ;
      RECT MASK 2 121.223 12.15 121.283 13.2 ;
      RECT MASK 2 121.497 12.15 121.557 13.2 ;
      RECT MASK 2 121.771 12.15 121.831 13.2 ;
      RECT MASK 2 122.045 12.15 122.105 13.2 ;
      RECT MASK 2 122.319 12.15 122.379 13.2 ;
      RECT MASK 2 122.593 12.15 122.653 13.2 ;
      RECT MASK 2 122.867 12.15 122.927 13.2 ;
      RECT MASK 2 123.141 12.15 123.201 13.2 ;
      RECT MASK 2 123.415 12.15 123.475 13.2 ;
      RECT MASK 2 123.689 12.15 123.749 13.2 ;
      RECT MASK 2 123.963 12.15 124.023 13.2 ;
      RECT MASK 2 124.237 12.15 124.297 13.2 ;
      RECT MASK 2 124.511 12.15 124.571 13.2 ;
      RECT MASK 2 124.785 12.15 124.845 13.2 ;
      RECT MASK 2 125.059 12.15 125.119 13.2 ;
      RECT MASK 2 125.333 12.15 125.393 13.2 ;
      RECT MASK 2 125.607 12.15 125.667 13.2 ;
      RECT MASK 2 125.881 12.15 125.941 13.2 ;
      RECT MASK 2 126.155 12.15 126.215 13.2 ;
      RECT MASK 2 126.429 12.15 126.489 13.2 ;
      RECT MASK 2 126.703 12.15 126.763 13.2 ;
      RECT MASK 2 126.977 12.15 127.037 13.2 ;
      RECT MASK 2 127.251 12.15 127.311 13.2 ;
      RECT MASK 2 127.525 12.15 127.585 13.2 ;
      RECT MASK 2 127.799 12.15 127.859 13.2 ;
      RECT MASK 2 128.073 12.15 128.133 13.2 ;
      RECT MASK 2 4.251 12.281 111.819 12.321 ;
      RECT MASK 2 8.356 12.448 8.871 12.488 ;
      RECT MASK 2 9.093 12.448 9.608 12.488 ;
      RECT MASK 2 10.016 12.448 10.531 12.488 ;
      RECT MASK 2 10.753 12.448 11.268 12.488 ;
      RECT MASK 2 22.373 12.448 22.888 12.488 ;
      RECT MASK 2 23.296 12.448 23.811 12.488 ;
      RECT MASK 2 24.033 12.448 24.548 12.488 ;
      RECT MASK 2 24.956 12.448 25.471 12.488 ;
      RECT MASK 2 25.659 12.448 26.081 12.488 ;
      RECT MASK 2 26.743 12.448 27.165 12.488 ;
      RECT MASK 2 27.446 12.448 27.629 12.488 ;
      RECT MASK 2 28.403 12.448 28.825 12.488 ;
      RECT MASK 2 28.979 12.448 29.401 12.488 ;
      RECT MASK 2 30.009 12.448 30.192 12.488 ;
      RECT MASK 2 30.639 12.448 31.061 12.488 ;
      RECT MASK 2 31.723 12.448 32.145 12.488 ;
      RECT MASK 2 32.299 12.448 32.721 12.488 ;
      RECT MASK 2 33.383 12.448 33.805 12.488 ;
      RECT MASK 2 34.086 12.448 34.601 12.488 ;
      RECT MASK 2 34.823 12.448 35.338 12.488 ;
      RECT MASK 2 35.653 12.448 36.168 12.488 ;
      RECT MASK 2 36.576 12.448 37.091 12.488 ;
      RECT MASK 2 37.279 12.448 37.701 12.488 ;
      RECT MASK 2 38.363 12.448 38.785 12.488 ;
      RECT MASK 2 38.939 12.448 39.361 12.488 ;
      RECT MASK 2 40.023 12.448 40.445 12.488 ;
      RECT MASK 2 40.726 12.448 40.909 12.488 ;
      RECT MASK 2 41.556 12.448 41.739 12.488 ;
      RECT MASK 2 42.259 12.448 42.681 12.488 ;
      RECT MASK 2 43.343 12.448 43.765 12.488 ;
      RECT MASK 2 43.953 12.448 44.468 12.488 ;
      RECT MASK 2 44.876 12.448 45.391 12.488 ;
      RECT MASK 2 45.706 12.448 46.221 12.488 ;
      RECT MASK 2 46.536 12.448 47.051 12.488 ;
      RECT MASK 2 47.239 12.448 47.661 12.488 ;
      RECT MASK 2 48.323 12.448 48.745 12.488 ;
      RECT MASK 2 48.933 12.448 49.448 12.488 ;
      RECT MASK 2 49.856 12.448 50.371 12.488 ;
      RECT MASK 2 50.593 12.448 51.108 12.488 ;
      RECT MASK 2 51.516 12.448 52.031 12.488 ;
      RECT MASK 2 52.253 12.448 52.768 12.488 ;
      RECT MASK 2 53.176 12.448 53.691 12.488 ;
      RECT MASK 2 53.879 12.448 54.301 12.488 ;
      RECT MASK 2 54.963 12.448 55.385 12.488 ;
      RECT MASK 2 55.573 12.448 55.756 12.488 ;
      RECT MASK 2 56.789 12.448 57.211 12.488 ;
      RECT MASK 2 57.365 12.448 57.787 12.488 ;
      RECT MASK 2 58.322 12.448 58.837 12.488 ;
      RECT MASK 2 59.059 12.448 59.574 12.488 ;
      RECT MASK 2 60.055 12.448 60.238 12.488 ;
      RECT MASK 2 60.719 12.448 61.234 12.488 ;
      RECT MASK 2 61.642 12.448 62.157 12.488 ;
      RECT MASK 2 62.472 12.448 62.655 12.488 ;
      RECT MASK 2 63.429 12.448 63.851 12.488 ;
      RECT MASK 2 64.005 12.448 64.427 12.488 ;
      RECT MASK 2 64.962 12.448 65.477 12.488 ;
      RECT MASK 2 65.699 12.448 66.214 12.488 ;
      RECT MASK 2 66.622 12.448 67.137 12.488 ;
      RECT MASK 2 67.359 12.448 67.874 12.488 ;
      RECT MASK 2 68.282 12.448 68.797 12.488 ;
      RECT MASK 2 69.019 12.448 69.534 12.488 ;
      RECT MASK 2 69.942 12.448 70.457 12.488 ;
      RECT MASK 2 70.679 12.448 71.194 12.488 ;
      RECT MASK 2 71.602 12.448 72.117 12.488 ;
      RECT MASK 2 72.339 12.448 72.854 12.488 ;
      RECT MASK 2 77.319 12.448 77.834 12.488 ;
      RECT MASK 2 78.242 12.448 78.757 12.488 ;
      RECT MASK 2 78.979 12.448 79.494 12.488 ;
      RECT MASK 2 79.902 12.448 80.417 12.488 ;
      RECT MASK 2 83.349 12.448 83.771 12.488 ;
      RECT MASK 2 83.925 12.448 84.347 12.488 ;
      RECT MASK 2 88.939 12.448 89.454 12.488 ;
      RECT MASK 2 89.862 12.448 90.377 12.488 ;
      RECT MASK 2 90.599 12.448 91.114 12.488 ;
      RECT MASK 2 91.522 12.448 92.037 12.488 ;
      RECT MASK 2 101.482 12.448 101.997 12.488 ;
      RECT MASK 2 102.219 12.448 102.734 12.488 ;
      RECT MASK 2 103.142 12.448 103.657 12.488 ;
      RECT MASK 2 103.879 12.448 104.394 12.488 ;
      RECT MASK 2 4.327 12.5425 4.507 12.5825 ;
      RECT MASK 2 111.563 12.5425 111.743 12.5825 ;
      RECT MASK 2 8.56 12.615 8.906 12.655 ;
      RECT MASK 2 9.058 12.615 9.404 12.655 ;
      RECT MASK 2 10.22 12.615 10.566 12.655 ;
      RECT MASK 2 10.718 12.615 11.064 12.655 ;
      RECT MASK 2 22.338 12.615 22.684 12.655 ;
      RECT MASK 2 23.5 12.615 23.846 12.655 ;
      RECT MASK 2 23.998 12.615 24.344 12.655 ;
      RECT MASK 2 25.16 12.615 25.506 12.655 ;
      RECT MASK 2 25.842 12.615 26.145 12.655 ;
      RECT MASK 2 26.679 12.615 26.982 12.655 ;
      RECT MASK 2 28.339 12.615 28.642 12.655 ;
      RECT MASK 2 29.162 12.615 29.465 12.655 ;
      RECT MASK 2 30.822 12.615 31.125 12.655 ;
      RECT MASK 2 31.659 12.615 31.962 12.655 ;
      RECT MASK 2 32.482 12.615 32.785 12.655 ;
      RECT MASK 2 33.319 12.615 33.622 12.655 ;
      RECT MASK 2 34.29 12.615 34.636 12.655 ;
      RECT MASK 2 34.788 12.615 35.134 12.655 ;
      RECT MASK 2 35.618 12.615 35.964 12.655 ;
      RECT MASK 2 36.78 12.615 37.126 12.655 ;
      RECT MASK 2 37.462 12.615 37.765 12.655 ;
      RECT MASK 2 38.299 12.615 38.602 12.655 ;
      RECT MASK 2 39.122 12.615 39.425 12.655 ;
      RECT MASK 2 39.959 12.615 40.262 12.655 ;
      RECT MASK 2 42.442 12.615 42.745 12.655 ;
      RECT MASK 2 43.279 12.615 43.582 12.655 ;
      RECT MASK 2 43.918 12.615 44.264 12.655 ;
      RECT MASK 2 45.08 12.615 45.426 12.655 ;
      RECT MASK 2 45.91 12.615 46.256 12.655 ;
      RECT MASK 2 46.74 12.615 47.086 12.655 ;
      RECT MASK 2 47.422 12.615 47.725 12.655 ;
      RECT MASK 2 48.259 12.615 48.562 12.655 ;
      RECT MASK 2 48.898 12.615 49.244 12.655 ;
      RECT MASK 2 50.06 12.615 50.406 12.655 ;
      RECT MASK 2 50.558 12.615 50.904 12.655 ;
      RECT MASK 2 51.72 12.615 52.066 12.655 ;
      RECT MASK 2 52.218 12.615 52.564 12.655 ;
      RECT MASK 2 53.38 12.615 53.726 12.655 ;
      RECT MASK 2 54.062 12.615 54.365 12.655 ;
      RECT MASK 2 54.899 12.615 55.202 12.655 ;
      RECT MASK 2 56.725 12.615 57.028 12.655 ;
      RECT MASK 2 57.548 12.615 57.851 12.655 ;
      RECT MASK 2 58.526 12.615 58.872 12.655 ;
      RECT MASK 2 59.024 12.615 59.37 12.655 ;
      RECT MASK 2 60.684 12.615 61.03 12.655 ;
      RECT MASK 2 61.846 12.615 62.192 12.655 ;
      RECT MASK 2 63.365 12.615 63.668 12.655 ;
      RECT MASK 2 64.188 12.615 64.491 12.655 ;
      RECT MASK 2 65.166 12.615 65.512 12.655 ;
      RECT MASK 2 65.664 12.615 66.01 12.655 ;
      RECT MASK 2 66.826 12.615 67.172 12.655 ;
      RECT MASK 2 67.324 12.615 67.67 12.655 ;
      RECT MASK 2 68.486 12.615 68.832 12.655 ;
      RECT MASK 2 68.984 12.615 69.33 12.655 ;
      RECT MASK 2 70.146 12.615 70.492 12.655 ;
      RECT MASK 2 70.644 12.615 70.99 12.655 ;
      RECT MASK 2 71.806 12.615 72.152 12.655 ;
      RECT MASK 2 72.304 12.615 72.65 12.655 ;
      RECT MASK 2 77.284 12.615 77.63 12.655 ;
      RECT MASK 2 78.446 12.615 78.792 12.655 ;
      RECT MASK 2 78.944 12.615 79.29 12.655 ;
      RECT MASK 2 80.106 12.615 80.452 12.655 ;
      RECT MASK 2 83.285 12.615 83.588 12.655 ;
      RECT MASK 2 84.108 12.615 84.411 12.655 ;
      RECT MASK 2 88.904 12.615 89.25 12.655 ;
      RECT MASK 2 90.066 12.615 90.412 12.655 ;
      RECT MASK 2 90.564 12.615 90.91 12.655 ;
      RECT MASK 2 91.726 12.615 92.072 12.655 ;
      RECT MASK 2 101.686 12.615 102.032 12.655 ;
      RECT MASK 2 102.184 12.615 102.53 12.655 ;
      RECT MASK 2 103.346 12.615 103.692 12.655 ;
      RECT MASK 2 103.844 12.615 104.19 12.655 ;
      RECT MASK 2 8.394 13.025 8.74 13.065 ;
      RECT MASK 2 9.224 13.025 9.57 13.065 ;
      RECT MASK 2 10.054 13.025 10.4 13.065 ;
      RECT MASK 2 10.884 13.025 11.23 13.065 ;
      RECT MASK 2 22.504 13.025 22.85 13.065 ;
      RECT MASK 2 23.334 13.025 23.68 13.065 ;
      RECT MASK 2 24.164 13.025 24.51 13.065 ;
      RECT MASK 2 24.994 13.025 25.34 13.065 ;
      RECT MASK 2 25.843 13.025 26.162 13.065 ;
      RECT MASK 2 26.662 13.025 26.981 13.065 ;
      RECT MASK 2 28.322 13.025 28.641 13.065 ;
      RECT MASK 2 29.163 13.025 29.482 13.065 ;
      RECT MASK 2 30.823 13.025 31.142 13.065 ;
      RECT MASK 2 31.642 13.025 31.961 13.065 ;
      RECT MASK 2 32.483 13.025 32.802 13.065 ;
      RECT MASK 2 33.302 13.025 33.621 13.065 ;
      RECT MASK 2 34.124 13.025 34.47 13.065 ;
      RECT MASK 2 34.954 13.025 35.3 13.065 ;
      RECT MASK 2 35.784 13.025 36.13 13.065 ;
      RECT MASK 2 36.614 13.025 36.96 13.065 ;
      RECT MASK 2 37.463 13.025 37.782 13.065 ;
      RECT MASK 2 38.282 13.025 38.601 13.065 ;
      RECT MASK 2 39.123 13.025 39.442 13.065 ;
      RECT MASK 2 39.942 13.025 40.261 13.065 ;
      RECT MASK 2 42.443 13.025 42.762 13.065 ;
      RECT MASK 2 43.262 13.025 43.581 13.065 ;
      RECT MASK 2 44.084 13.025 44.43 13.065 ;
      RECT MASK 2 44.914 13.025 45.26 13.065 ;
      RECT MASK 2 45.744 13.025 46.09 13.065 ;
      RECT MASK 2 46.574 13.025 46.92 13.065 ;
      RECT MASK 2 47.423 13.025 47.742 13.065 ;
      RECT MASK 2 48.242 13.025 48.561 13.065 ;
      RECT MASK 2 49.064 13.025 49.41 13.065 ;
      RECT MASK 2 49.894 13.025 50.24 13.065 ;
      RECT MASK 2 50.724 13.025 51.07 13.065 ;
      RECT MASK 2 51.554 13.025 51.9 13.065 ;
      RECT MASK 2 52.384 13.025 52.73 13.065 ;
      RECT MASK 2 53.214 13.025 53.56 13.065 ;
      RECT MASK 2 54.063 13.025 54.382 13.065 ;
      RECT MASK 2 54.882 13.025 55.201 13.065 ;
      RECT MASK 2 56.708 13.025 57.027 13.065 ;
      RECT MASK 2 57.549 13.025 57.868 13.065 ;
      RECT MASK 2 58.36 13.025 58.706 13.065 ;
      RECT MASK 2 59.19 13.025 59.536 13.065 ;
      RECT MASK 2 60.85 13.025 61.196 13.065 ;
      RECT MASK 2 61.68 13.025 62.026 13.065 ;
      RECT MASK 2 63.348 13.025 63.667 13.065 ;
      RECT MASK 2 64.189 13.025 64.508 13.065 ;
      RECT MASK 2 65 13.025 65.346 13.065 ;
      RECT MASK 2 65.83 13.025 66.176 13.065 ;
      RECT MASK 2 66.66 13.025 67.006 13.065 ;
      RECT MASK 2 67.49 13.025 67.836 13.065 ;
      RECT MASK 2 68.32 13.025 68.666 13.065 ;
      RECT MASK 2 69.15 13.025 69.496 13.065 ;
      RECT MASK 2 69.98 13.025 70.326 13.065 ;
      RECT MASK 2 70.81 13.025 71.156 13.065 ;
      RECT MASK 2 71.64 13.025 71.986 13.065 ;
      RECT MASK 2 72.47 13.025 72.816 13.065 ;
      RECT MASK 2 77.45 13.025 77.796 13.065 ;
      RECT MASK 2 78.28 13.025 78.626 13.065 ;
      RECT MASK 2 79.11 13.025 79.456 13.065 ;
      RECT MASK 2 79.94 13.025 80.286 13.065 ;
      RECT MASK 2 83.268 13.025 83.587 13.065 ;
      RECT MASK 2 84.109 13.025 84.428 13.065 ;
      RECT MASK 2 89.07 13.025 89.416 13.065 ;
      RECT MASK 2 89.9 13.025 90.246 13.065 ;
      RECT MASK 2 90.73 13.025 91.076 13.065 ;
      RECT MASK 2 91.56 13.025 91.906 13.065 ;
      RECT MASK 2 101.52 13.025 101.866 13.065 ;
      RECT MASK 2 102.35 13.025 102.696 13.065 ;
      RECT MASK 2 103.18 13.025 103.526 13.065 ;
      RECT MASK 2 104.01 13.025 104.356 13.065 ;
      RECT MASK 2 4.327 13.0975 4.507 13.1375 ;
      RECT MASK 2 111.563 13.0975 111.743 13.1375 ;
      RECT MASK 2 8.522 13.192 8.871 13.232 ;
      RECT MASK 2 9.093 13.192 9.442 13.232 ;
      RECT MASK 2 10.182 13.192 10.531 13.232 ;
      RECT MASK 2 10.753 13.192 11.102 13.232 ;
      RECT MASK 2 22.373 13.192 22.722 13.232 ;
      RECT MASK 2 23.462 13.192 23.811 13.232 ;
      RECT MASK 2 24.033 13.192 24.382 13.232 ;
      RECT MASK 2 25.122 13.192 25.471 13.232 ;
      RECT MASK 2 25.658 13.192 26.208 13.232 ;
      RECT MASK 2 26.616 13.192 27.166 13.232 ;
      RECT MASK 2 27.446 13.192 27.629 13.232 ;
      RECT MASK 2 28.276 13.192 28.826 13.232 ;
      RECT MASK 2 28.978 13.192 29.528 13.232 ;
      RECT MASK 2 30.009 13.192 30.192 13.232 ;
      RECT MASK 2 30.638 13.192 31.188 13.232 ;
      RECT MASK 2 31.596 13.192 32.146 13.232 ;
      RECT MASK 2 32.298 13.192 32.848 13.232 ;
      RECT MASK 2 33.256 13.192 33.806 13.232 ;
      RECT MASK 2 34.252 13.192 34.601 13.232 ;
      RECT MASK 2 34.823 13.192 35.172 13.232 ;
      RECT MASK 2 35.653 13.192 36.002 13.232 ;
      RECT MASK 2 36.742 13.192 37.091 13.232 ;
      RECT MASK 2 37.278 13.192 37.828 13.232 ;
      RECT MASK 2 38.236 13.192 38.786 13.232 ;
      RECT MASK 2 38.938 13.192 39.488 13.232 ;
      RECT MASK 2 39.896 13.192 40.446 13.232 ;
      RECT MASK 2 40.726 13.192 40.909 13.232 ;
      RECT MASK 2 41.556 13.192 41.739 13.232 ;
      RECT MASK 2 42.258 13.192 42.808 13.232 ;
      RECT MASK 2 43.216 13.192 43.766 13.232 ;
      RECT MASK 2 43.953 13.192 44.302 13.232 ;
      RECT MASK 2 45.042 13.192 45.391 13.232 ;
      RECT MASK 2 45.872 13.192 46.221 13.232 ;
      RECT MASK 2 46.702 13.192 47.051 13.232 ;
      RECT MASK 2 47.238 13.192 47.788 13.232 ;
      RECT MASK 2 48.196 13.192 48.746 13.232 ;
      RECT MASK 2 48.933 13.192 49.282 13.232 ;
      RECT MASK 2 50.022 13.192 50.371 13.232 ;
      RECT MASK 2 50.593 13.192 50.942 13.232 ;
      RECT MASK 2 51.682 13.192 52.031 13.232 ;
      RECT MASK 2 52.253 13.192 52.602 13.232 ;
      RECT MASK 2 53.342 13.192 53.691 13.232 ;
      RECT MASK 2 53.878 13.192 54.428 13.232 ;
      RECT MASK 2 54.836 13.192 55.386 13.232 ;
      RECT MASK 2 55.573 13.192 55.756 13.232 ;
      RECT MASK 2 56.662 13.192 57.212 13.232 ;
      RECT MASK 2 57.364 13.192 57.914 13.232 ;
      RECT MASK 2 58.488 13.192 58.837 13.232 ;
      RECT MASK 2 59.059 13.192 59.408 13.232 ;
      RECT MASK 2 60.055 13.192 60.238 13.232 ;
      RECT MASK 2 60.719 13.192 61.068 13.232 ;
      RECT MASK 2 61.808 13.192 62.157 13.232 ;
      RECT MASK 2 62.472 13.192 62.655 13.232 ;
      RECT MASK 2 63.302 13.192 63.852 13.232 ;
      RECT MASK 2 64.004 13.192 64.554 13.232 ;
      RECT MASK 2 65.128 13.192 65.477 13.232 ;
      RECT MASK 2 65.699 13.192 66.048 13.232 ;
      RECT MASK 2 66.788 13.192 67.137 13.232 ;
      RECT MASK 2 67.359 13.192 67.708 13.232 ;
      RECT MASK 2 68.448 13.192 68.797 13.232 ;
      RECT MASK 2 69.019 13.192 69.368 13.232 ;
      RECT MASK 2 70.108 13.192 70.457 13.232 ;
      RECT MASK 2 70.679 13.192 71.028 13.232 ;
      RECT MASK 2 71.768 13.192 72.117 13.232 ;
      RECT MASK 2 72.339 13.192 72.688 13.232 ;
      RECT MASK 2 77.319 13.192 77.668 13.232 ;
      RECT MASK 2 78.408 13.192 78.757 13.232 ;
      RECT MASK 2 78.979 13.192 79.328 13.232 ;
      RECT MASK 2 80.068 13.192 80.417 13.232 ;
      RECT MASK 2 83.222 13.192 83.772 13.232 ;
      RECT MASK 2 83.924 13.192 84.474 13.232 ;
      RECT MASK 2 88.939 13.192 89.288 13.232 ;
      RECT MASK 2 90.028 13.192 90.377 13.232 ;
      RECT MASK 2 90.599 13.192 90.948 13.232 ;
      RECT MASK 2 91.688 13.192 92.037 13.232 ;
      RECT MASK 2 101.648 13.192 101.997 13.232 ;
      RECT MASK 2 102.219 13.192 102.568 13.232 ;
      RECT MASK 2 103.308 13.192 103.657 13.232 ;
      RECT MASK 2 103.879 13.192 104.228 13.232 ;
      RECT MASK 2 4.251 13.359 111.819 13.399 ;
      RECT MASK 2 4.362 13.7 111.708 13.74 ;
      RECT MASK 2 4.362 13.86 111.708 13.9 ;
      RECT MASK 2 116.291 13.86 116.351 14.91 ;
      RECT MASK 2 116.565 13.86 116.625 14.91 ;
      RECT MASK 2 116.839 13.86 116.899 14.91 ;
      RECT MASK 2 117.113 13.86 117.173 14.91 ;
      RECT MASK 2 117.387 13.86 117.447 14.91 ;
      RECT MASK 2 117.661 13.86 117.721 14.91 ;
      RECT MASK 2 117.935 13.86 117.995 14.91 ;
      RECT MASK 2 118.209 13.86 118.269 14.91 ;
      RECT MASK 2 118.483 13.86 118.543 14.91 ;
      RECT MASK 2 118.757 13.86 118.817 14.91 ;
      RECT MASK 2 119.031 13.86 119.091 14.91 ;
      RECT MASK 2 119.305 13.86 119.365 14.91 ;
      RECT MASK 2 119.579 13.86 119.639 14.91 ;
      RECT MASK 2 119.853 13.86 119.913 14.91 ;
      RECT MASK 2 120.127 13.86 120.187 14.91 ;
      RECT MASK 2 120.401 13.86 120.461 14.91 ;
      RECT MASK 2 120.675 13.86 120.735 14.91 ;
      RECT MASK 2 120.949 13.86 121.009 14.91 ;
      RECT MASK 2 121.223 13.86 121.283 14.91 ;
      RECT MASK 2 121.497 13.86 121.557 14.91 ;
      RECT MASK 2 121.771 13.86 121.831 14.91 ;
      RECT MASK 2 122.045 13.86 122.105 14.91 ;
      RECT MASK 2 122.319 13.86 122.379 14.91 ;
      RECT MASK 2 122.593 13.86 122.653 14.91 ;
      RECT MASK 2 122.867 13.86 122.927 14.91 ;
      RECT MASK 2 123.141 13.86 123.201 14.91 ;
      RECT MASK 2 123.415 13.86 123.475 14.91 ;
      RECT MASK 2 123.689 13.86 123.749 14.91 ;
      RECT MASK 2 123.963 13.86 124.023 14.91 ;
      RECT MASK 2 124.237 13.86 124.297 14.91 ;
      RECT MASK 2 124.511 13.86 124.571 14.91 ;
      RECT MASK 2 124.785 13.86 124.845 14.91 ;
      RECT MASK 2 125.059 13.86 125.119 14.91 ;
      RECT MASK 2 125.333 13.86 125.393 14.91 ;
      RECT MASK 2 125.607 13.86 125.667 14.91 ;
      RECT MASK 2 125.881 13.86 125.941 14.91 ;
      RECT MASK 2 126.155 13.86 126.215 14.91 ;
      RECT MASK 2 126.429 13.86 126.489 14.91 ;
      RECT MASK 2 126.703 13.86 126.763 14.91 ;
      RECT MASK 2 126.977 13.86 127.037 14.91 ;
      RECT MASK 2 127.251 13.86 127.311 14.91 ;
      RECT MASK 2 127.525 13.86 127.585 14.91 ;
      RECT MASK 2 127.799 13.86 127.859 14.91 ;
      RECT MASK 2 128.073 13.86 128.133 14.91 ;
      RECT MASK 2 4.251 14.201 111.819 14.241 ;
      RECT MASK 2 5.036 14.368 5.586 14.408 ;
      RECT MASK 2 5.738 14.368 6.288 14.408 ;
      RECT MASK 2 6.696 14.368 7.246 14.408 ;
      RECT MASK 2 7.398 14.368 7.948 14.408 ;
      RECT MASK 2 8.356 14.368 8.906 14.408 ;
      RECT MASK 2 9.058 14.368 9.608 14.408 ;
      RECT MASK 2 10.016 14.368 10.566 14.408 ;
      RECT MASK 2 10.718 14.368 11.268 14.408 ;
      RECT MASK 2 11.676 14.368 12.226 14.408 ;
      RECT MASK 2 12.378 14.368 12.928 14.408 ;
      RECT MASK 2 13.336 14.368 13.886 14.408 ;
      RECT MASK 2 14.038 14.368 14.588 14.408 ;
      RECT MASK 2 14.996 14.368 15.546 14.408 ;
      RECT MASK 2 15.698 14.368 16.248 14.408 ;
      RECT MASK 2 16.656 14.368 17.206 14.408 ;
      RECT MASK 2 17.358 14.368 17.908 14.408 ;
      RECT MASK 2 18.316 14.368 18.866 14.408 ;
      RECT MASK 2 19.018 14.368 19.568 14.408 ;
      RECT MASK 2 19.976 14.368 20.526 14.408 ;
      RECT MASK 2 20.678 14.368 21.228 14.408 ;
      RECT MASK 2 21.636 14.368 22.186 14.408 ;
      RECT MASK 2 22.338 14.368 22.888 14.408 ;
      RECT MASK 2 23.296 14.368 23.846 14.408 ;
      RECT MASK 2 23.998 14.368 24.548 14.408 ;
      RECT MASK 2 24.956 14.368 25.506 14.408 ;
      RECT MASK 2 25.658 14.368 26.208 14.408 ;
      RECT MASK 2 26.616 14.368 27.166 14.408 ;
      RECT MASK 2 27.318 14.368 27.868 14.408 ;
      RECT MASK 2 28.276 14.368 28.826 14.408 ;
      RECT MASK 2 28.978 14.368 29.528 14.408 ;
      RECT MASK 2 29.936 14.368 30.486 14.408 ;
      RECT MASK 2 30.638 14.368 31.188 14.408 ;
      RECT MASK 2 31.596 14.368 32.146 14.408 ;
      RECT MASK 2 32.298 14.368 32.848 14.408 ;
      RECT MASK 2 33.256 14.368 33.806 14.408 ;
      RECT MASK 2 33.958 14.368 34.508 14.408 ;
      RECT MASK 2 34.916 14.368 35.466 14.408 ;
      RECT MASK 2 35.618 14.368 36.168 14.408 ;
      RECT MASK 2 36.576 14.368 37.126 14.408 ;
      RECT MASK 2 37.278 14.368 37.828 14.408 ;
      RECT MASK 2 38.236 14.368 38.786 14.408 ;
      RECT MASK 2 38.938 14.368 39.488 14.408 ;
      RECT MASK 2 39.896 14.368 40.446 14.408 ;
      RECT MASK 2 40.598 14.368 41.148 14.408 ;
      RECT MASK 2 41.556 14.368 42.106 14.408 ;
      RECT MASK 2 42.258 14.368 42.808 14.408 ;
      RECT MASK 2 43.216 14.368 43.766 14.408 ;
      RECT MASK 2 43.918 14.368 44.468 14.408 ;
      RECT MASK 2 44.876 14.368 45.426 14.408 ;
      RECT MASK 2 45.578 14.368 46.128 14.408 ;
      RECT MASK 2 46.536 14.368 47.086 14.408 ;
      RECT MASK 2 47.238 14.368 47.788 14.408 ;
      RECT MASK 2 48.196 14.368 48.746 14.408 ;
      RECT MASK 2 48.898 14.368 49.448 14.408 ;
      RECT MASK 2 49.856 14.368 50.406 14.408 ;
      RECT MASK 2 50.558 14.368 51.108 14.408 ;
      RECT MASK 2 51.516 14.368 52.066 14.408 ;
      RECT MASK 2 52.218 14.368 52.768 14.408 ;
      RECT MASK 2 53.176 14.368 53.726 14.408 ;
      RECT MASK 2 53.878 14.368 54.428 14.408 ;
      RECT MASK 2 54.836 14.368 55.386 14.408 ;
      RECT MASK 2 55.538 14.368 56.088 14.408 ;
      RECT MASK 2 56.662 14.368 57.212 14.408 ;
      RECT MASK 2 57.364 14.368 57.914 14.408 ;
      RECT MASK 2 58.322 14.368 58.872 14.408 ;
      RECT MASK 2 59.024 14.368 59.574 14.408 ;
      RECT MASK 2 59.982 14.368 60.532 14.408 ;
      RECT MASK 2 60.684 14.368 61.234 14.408 ;
      RECT MASK 2 61.642 14.368 62.192 14.408 ;
      RECT MASK 2 62.344 14.368 62.894 14.408 ;
      RECT MASK 2 63.302 14.368 63.852 14.408 ;
      RECT MASK 2 64.004 14.368 64.554 14.408 ;
      RECT MASK 2 64.962 14.368 65.512 14.408 ;
      RECT MASK 2 65.664 14.368 66.214 14.408 ;
      RECT MASK 2 66.622 14.368 67.172 14.408 ;
      RECT MASK 2 67.324 14.368 67.874 14.408 ;
      RECT MASK 2 68.282 14.368 68.832 14.408 ;
      RECT MASK 2 68.984 14.368 69.534 14.408 ;
      RECT MASK 2 69.942 14.368 70.492 14.408 ;
      RECT MASK 2 70.644 14.368 71.194 14.408 ;
      RECT MASK 2 71.602 14.368 72.152 14.408 ;
      RECT MASK 2 72.304 14.368 72.854 14.408 ;
      RECT MASK 2 73.262 14.368 73.812 14.408 ;
      RECT MASK 2 73.964 14.368 74.514 14.408 ;
      RECT MASK 2 74.922 14.368 75.472 14.408 ;
      RECT MASK 2 75.624 14.368 76.174 14.408 ;
      RECT MASK 2 76.582 14.368 77.132 14.408 ;
      RECT MASK 2 77.284 14.368 77.834 14.408 ;
      RECT MASK 2 78.242 14.368 78.792 14.408 ;
      RECT MASK 2 78.944 14.368 79.494 14.408 ;
      RECT MASK 2 79.902 14.368 80.452 14.408 ;
      RECT MASK 2 80.604 14.368 81.154 14.408 ;
      RECT MASK 2 81.562 14.368 82.112 14.408 ;
      RECT MASK 2 82.264 14.368 82.814 14.408 ;
      RECT MASK 2 83.222 14.368 83.772 14.408 ;
      RECT MASK 2 83.924 14.368 84.474 14.408 ;
      RECT MASK 2 84.882 14.368 85.432 14.408 ;
      RECT MASK 2 85.584 14.368 86.134 14.408 ;
      RECT MASK 2 86.542 14.368 87.092 14.408 ;
      RECT MASK 2 87.244 14.368 87.794 14.408 ;
      RECT MASK 2 88.202 14.368 88.752 14.408 ;
      RECT MASK 2 88.904 14.368 89.454 14.408 ;
      RECT MASK 2 89.862 14.368 90.412 14.408 ;
      RECT MASK 2 90.564 14.368 91.114 14.408 ;
      RECT MASK 2 91.522 14.368 92.072 14.408 ;
      RECT MASK 2 92.224 14.368 92.774 14.408 ;
      RECT MASK 2 93.182 14.368 93.732 14.408 ;
      RECT MASK 2 93.884 14.368 94.434 14.408 ;
      RECT MASK 2 94.842 14.368 95.392 14.408 ;
      RECT MASK 2 95.544 14.368 96.094 14.408 ;
      RECT MASK 2 96.502 14.368 97.052 14.408 ;
      RECT MASK 2 97.204 14.368 97.754 14.408 ;
      RECT MASK 2 98.162 14.368 98.712 14.408 ;
      RECT MASK 2 98.864 14.368 99.414 14.408 ;
      RECT MASK 2 99.822 14.368 100.372 14.408 ;
      RECT MASK 2 100.524 14.368 101.074 14.408 ;
      RECT MASK 2 101.482 14.368 102.032 14.408 ;
      RECT MASK 2 102.184 14.368 102.734 14.408 ;
      RECT MASK 2 103.142 14.368 103.692 14.408 ;
      RECT MASK 2 103.844 14.368 104.394 14.408 ;
      RECT MASK 2 104.802 14.368 105.352 14.408 ;
      RECT MASK 2 105.504 14.368 106.054 14.408 ;
      RECT MASK 2 106.462 14.368 107.012 14.408 ;
      RECT MASK 2 107.164 14.368 107.714 14.408 ;
      RECT MASK 2 108.122 14.368 108.672 14.408 ;
      RECT MASK 2 108.824 14.368 109.374 14.408 ;
      RECT MASK 2 109.782 14.368 110.332 14.408 ;
      RECT MASK 2 110.484 14.368 111.034 14.408 ;
      RECT MASK 2 4.327 14.4625 4.507 14.5025 ;
      RECT MASK 2 111.563 14.4625 111.743 14.5025 ;
      RECT MASK 2 5.082 14.535 5.401 14.575 ;
      RECT MASK 2 5.923 14.535 6.242 14.575 ;
      RECT MASK 2 6.742 14.535 7.061 14.575 ;
      RECT MASK 2 7.583 14.535 7.902 14.575 ;
      RECT MASK 2 8.402 14.535 8.721 14.575 ;
      RECT MASK 2 9.243 14.535 9.562 14.575 ;
      RECT MASK 2 10.062 14.535 10.381 14.575 ;
      RECT MASK 2 10.903 14.535 11.222 14.575 ;
      RECT MASK 2 11.722 14.535 12.041 14.575 ;
      RECT MASK 2 12.563 14.535 12.882 14.575 ;
      RECT MASK 2 13.382 14.535 13.701 14.575 ;
      RECT MASK 2 14.223 14.535 14.542 14.575 ;
      RECT MASK 2 15.042 14.535 15.361 14.575 ;
      RECT MASK 2 15.883 14.535 16.202 14.575 ;
      RECT MASK 2 16.702 14.535 17.021 14.575 ;
      RECT MASK 2 17.543 14.535 17.862 14.575 ;
      RECT MASK 2 18.362 14.535 18.681 14.575 ;
      RECT MASK 2 19.203 14.535 19.522 14.575 ;
      RECT MASK 2 20.022 14.535 20.341 14.575 ;
      RECT MASK 2 20.863 14.535 21.182 14.575 ;
      RECT MASK 2 21.682 14.535 22.001 14.575 ;
      RECT MASK 2 22.523 14.535 22.842 14.575 ;
      RECT MASK 2 23.342 14.535 23.661 14.575 ;
      RECT MASK 2 24.183 14.535 24.502 14.575 ;
      RECT MASK 2 25.002 14.535 25.321 14.575 ;
      RECT MASK 2 25.843 14.535 26.162 14.575 ;
      RECT MASK 2 26.662 14.535 26.981 14.575 ;
      RECT MASK 2 27.503 14.535 27.822 14.575 ;
      RECT MASK 2 28.322 14.535 28.641 14.575 ;
      RECT MASK 2 29.163 14.535 29.482 14.575 ;
      RECT MASK 2 29.982 14.535 30.301 14.575 ;
      RECT MASK 2 30.823 14.535 31.142 14.575 ;
      RECT MASK 2 31.642 14.535 31.961 14.575 ;
      RECT MASK 2 32.483 14.535 32.802 14.575 ;
      RECT MASK 2 33.302 14.535 33.621 14.575 ;
      RECT MASK 2 34.143 14.535 34.462 14.575 ;
      RECT MASK 2 34.962 14.535 35.281 14.575 ;
      RECT MASK 2 35.803 14.535 36.122 14.575 ;
      RECT MASK 2 36.622 14.535 36.941 14.575 ;
      RECT MASK 2 37.463 14.535 37.782 14.575 ;
      RECT MASK 2 38.282 14.535 38.601 14.575 ;
      RECT MASK 2 39.123 14.535 39.442 14.575 ;
      RECT MASK 2 39.942 14.535 40.261 14.575 ;
      RECT MASK 2 40.783 14.535 41.102 14.575 ;
      RECT MASK 2 41.602 14.535 41.921 14.575 ;
      RECT MASK 2 42.443 14.535 42.762 14.575 ;
      RECT MASK 2 43.262 14.535 43.581 14.575 ;
      RECT MASK 2 44.103 14.535 44.422 14.575 ;
      RECT MASK 2 44.922 14.535 45.241 14.575 ;
      RECT MASK 2 45.763 14.535 46.082 14.575 ;
      RECT MASK 2 46.582 14.535 46.901 14.575 ;
      RECT MASK 2 47.423 14.535 47.742 14.575 ;
      RECT MASK 2 48.242 14.535 48.561 14.575 ;
      RECT MASK 2 49.083 14.535 49.402 14.575 ;
      RECT MASK 2 49.902 14.535 50.221 14.575 ;
      RECT MASK 2 50.743 14.535 51.062 14.575 ;
      RECT MASK 2 51.562 14.535 51.881 14.575 ;
      RECT MASK 2 52.403 14.535 52.722 14.575 ;
      RECT MASK 2 53.222 14.535 53.541 14.575 ;
      RECT MASK 2 54.063 14.535 54.382 14.575 ;
      RECT MASK 2 54.882 14.535 55.201 14.575 ;
      RECT MASK 2 55.723 14.535 56.042 14.575 ;
      RECT MASK 2 56.708 14.535 57.027 14.575 ;
      RECT MASK 2 57.549 14.535 57.868 14.575 ;
      RECT MASK 2 58.368 14.535 58.687 14.575 ;
      RECT MASK 2 59.209 14.535 59.528 14.575 ;
      RECT MASK 2 60.028 14.535 60.347 14.575 ;
      RECT MASK 2 60.869 14.535 61.188 14.575 ;
      RECT MASK 2 61.688 14.535 62.007 14.575 ;
      RECT MASK 2 62.529 14.535 62.848 14.575 ;
      RECT MASK 2 63.348 14.535 63.667 14.575 ;
      RECT MASK 2 64.189 14.535 64.508 14.575 ;
      RECT MASK 2 65.008 14.535 65.327 14.575 ;
      RECT MASK 2 65.849 14.535 66.168 14.575 ;
      RECT MASK 2 66.668 14.535 66.987 14.575 ;
      RECT MASK 2 67.509 14.535 67.828 14.575 ;
      RECT MASK 2 68.328 14.535 68.647 14.575 ;
      RECT MASK 2 69.169 14.535 69.488 14.575 ;
      RECT MASK 2 69.988 14.535 70.307 14.575 ;
      RECT MASK 2 70.829 14.535 71.148 14.575 ;
      RECT MASK 2 71.648 14.535 71.967 14.575 ;
      RECT MASK 2 72.489 14.535 72.808 14.575 ;
      RECT MASK 2 73.308 14.535 73.627 14.575 ;
      RECT MASK 2 74.149 14.535 74.468 14.575 ;
      RECT MASK 2 74.968 14.535 75.287 14.575 ;
      RECT MASK 2 75.809 14.535 76.128 14.575 ;
      RECT MASK 2 76.628 14.535 76.947 14.575 ;
      RECT MASK 2 77.469 14.535 77.788 14.575 ;
      RECT MASK 2 78.288 14.535 78.607 14.575 ;
      RECT MASK 2 79.129 14.535 79.448 14.575 ;
      RECT MASK 2 79.948 14.535 80.267 14.575 ;
      RECT MASK 2 80.789 14.535 81.108 14.575 ;
      RECT MASK 2 81.608 14.535 81.927 14.575 ;
      RECT MASK 2 82.449 14.535 82.768 14.575 ;
      RECT MASK 2 83.268 14.535 83.587 14.575 ;
      RECT MASK 2 84.109 14.535 84.428 14.575 ;
      RECT MASK 2 84.928 14.535 85.247 14.575 ;
      RECT MASK 2 85.769 14.535 86.088 14.575 ;
      RECT MASK 2 86.588 14.535 86.907 14.575 ;
      RECT MASK 2 87.429 14.535 87.748 14.575 ;
      RECT MASK 2 88.248 14.535 88.567 14.575 ;
      RECT MASK 2 89.089 14.535 89.408 14.575 ;
      RECT MASK 2 89.908 14.535 90.227 14.575 ;
      RECT MASK 2 90.749 14.535 91.068 14.575 ;
      RECT MASK 2 91.568 14.535 91.887 14.575 ;
      RECT MASK 2 92.409 14.535 92.728 14.575 ;
      RECT MASK 2 93.228 14.535 93.547 14.575 ;
      RECT MASK 2 94.069 14.535 94.388 14.575 ;
      RECT MASK 2 94.888 14.535 95.207 14.575 ;
      RECT MASK 2 95.729 14.535 96.048 14.575 ;
      RECT MASK 2 96.548 14.535 96.867 14.575 ;
      RECT MASK 2 97.389 14.535 97.708 14.575 ;
      RECT MASK 2 98.208 14.535 98.527 14.575 ;
      RECT MASK 2 99.049 14.535 99.368 14.575 ;
      RECT MASK 2 99.868 14.535 100.187 14.575 ;
      RECT MASK 2 100.709 14.535 101.028 14.575 ;
      RECT MASK 2 101.528 14.535 101.847 14.575 ;
      RECT MASK 2 102.369 14.535 102.688 14.575 ;
      RECT MASK 2 103.188 14.535 103.507 14.575 ;
      RECT MASK 2 104.029 14.535 104.348 14.575 ;
      RECT MASK 2 104.848 14.535 105.167 14.575 ;
      RECT MASK 2 105.689 14.535 106.008 14.575 ;
      RECT MASK 2 106.508 14.535 106.827 14.575 ;
      RECT MASK 2 107.349 14.535 107.668 14.575 ;
      RECT MASK 2 108.168 14.535 108.487 14.575 ;
      RECT MASK 2 109.009 14.535 109.328 14.575 ;
      RECT MASK 2 109.828 14.535 110.147 14.575 ;
      RECT MASK 2 110.669 14.535 110.988 14.575 ;
      RECT MASK 2 5.099 14.945 5.402 14.985 ;
      RECT MASK 2 5.922 14.945 6.225 14.985 ;
      RECT MASK 2 6.759 14.945 7.062 14.985 ;
      RECT MASK 2 7.582 14.945 7.885 14.985 ;
      RECT MASK 2 8.419 14.945 8.722 14.985 ;
      RECT MASK 2 9.242 14.945 9.545 14.985 ;
      RECT MASK 2 10.079 14.945 10.382 14.985 ;
      RECT MASK 2 10.902 14.945 11.205 14.985 ;
      RECT MASK 2 11.739 14.945 12.042 14.985 ;
      RECT MASK 2 12.562 14.945 12.865 14.985 ;
      RECT MASK 2 13.399 14.945 13.702 14.985 ;
      RECT MASK 2 14.222 14.945 14.525 14.985 ;
      RECT MASK 2 15.059 14.945 15.362 14.985 ;
      RECT MASK 2 15.882 14.945 16.185 14.985 ;
      RECT MASK 2 16.719 14.945 17.022 14.985 ;
      RECT MASK 2 17.542 14.945 17.845 14.985 ;
      RECT MASK 2 18.379 14.945 18.682 14.985 ;
      RECT MASK 2 19.202 14.945 19.505 14.985 ;
      RECT MASK 2 20.039 14.945 20.342 14.985 ;
      RECT MASK 2 20.862 14.945 21.165 14.985 ;
      RECT MASK 2 21.699 14.945 22.002 14.985 ;
      RECT MASK 2 22.522 14.945 22.825 14.985 ;
      RECT MASK 2 23.359 14.945 23.662 14.985 ;
      RECT MASK 2 24.182 14.945 24.485 14.985 ;
      RECT MASK 2 25.019 14.945 25.322 14.985 ;
      RECT MASK 2 25.842 14.945 26.145 14.985 ;
      RECT MASK 2 26.679 14.945 26.982 14.985 ;
      RECT MASK 2 27.502 14.945 27.805 14.985 ;
      RECT MASK 2 28.339 14.945 28.642 14.985 ;
      RECT MASK 2 29.162 14.945 29.465 14.985 ;
      RECT MASK 2 29.999 14.945 30.302 14.985 ;
      RECT MASK 2 30.822 14.945 31.125 14.985 ;
      RECT MASK 2 31.659 14.945 31.962 14.985 ;
      RECT MASK 2 32.482 14.945 32.785 14.985 ;
      RECT MASK 2 33.319 14.945 33.622 14.985 ;
      RECT MASK 2 34.142 14.945 34.445 14.985 ;
      RECT MASK 2 34.979 14.945 35.282 14.985 ;
      RECT MASK 2 35.802 14.945 36.105 14.985 ;
      RECT MASK 2 36.639 14.945 36.942 14.985 ;
      RECT MASK 2 37.462 14.945 37.765 14.985 ;
      RECT MASK 2 38.299 14.945 38.602 14.985 ;
      RECT MASK 2 39.122 14.945 39.425 14.985 ;
      RECT MASK 2 39.959 14.945 40.262 14.985 ;
      RECT MASK 2 40.782 14.945 41.085 14.985 ;
      RECT MASK 2 41.619 14.945 41.922 14.985 ;
      RECT MASK 2 42.442 14.945 42.745 14.985 ;
      RECT MASK 2 43.279 14.945 43.582 14.985 ;
      RECT MASK 2 44.102 14.945 44.405 14.985 ;
      RECT MASK 2 44.939 14.945 45.242 14.985 ;
      RECT MASK 2 45.762 14.945 46.065 14.985 ;
      RECT MASK 2 46.599 14.945 46.902 14.985 ;
      RECT MASK 2 47.422 14.945 47.725 14.985 ;
      RECT MASK 2 48.259 14.945 48.562 14.985 ;
      RECT MASK 2 49.082 14.945 49.385 14.985 ;
      RECT MASK 2 49.919 14.945 50.222 14.985 ;
      RECT MASK 2 50.742 14.945 51.045 14.985 ;
      RECT MASK 2 51.579 14.945 51.882 14.985 ;
      RECT MASK 2 52.402 14.945 52.705 14.985 ;
      RECT MASK 2 53.239 14.945 53.542 14.985 ;
      RECT MASK 2 54.062 14.945 54.365 14.985 ;
      RECT MASK 2 54.899 14.945 55.202 14.985 ;
      RECT MASK 2 55.722 14.945 56.025 14.985 ;
      RECT MASK 2 56.725 14.945 57.028 14.985 ;
      RECT MASK 2 57.548 14.945 57.851 14.985 ;
      RECT MASK 2 58.385 14.945 58.688 14.985 ;
      RECT MASK 2 59.208 14.945 59.511 14.985 ;
      RECT MASK 2 60.045 14.945 60.348 14.985 ;
      RECT MASK 2 60.868 14.945 61.171 14.985 ;
      RECT MASK 2 61.705 14.945 62.008 14.985 ;
      RECT MASK 2 62.528 14.945 62.831 14.985 ;
      RECT MASK 2 63.365 14.945 63.668 14.985 ;
      RECT MASK 2 64.188 14.945 64.491 14.985 ;
      RECT MASK 2 65.025 14.945 65.328 14.985 ;
      RECT MASK 2 65.848 14.945 66.151 14.985 ;
      RECT MASK 2 66.685 14.945 66.988 14.985 ;
      RECT MASK 2 67.508 14.945 67.811 14.985 ;
      RECT MASK 2 68.345 14.945 68.648 14.985 ;
      RECT MASK 2 69.168 14.945 69.471 14.985 ;
      RECT MASK 2 70.005 14.945 70.308 14.985 ;
      RECT MASK 2 70.828 14.945 71.131 14.985 ;
      RECT MASK 2 71.665 14.945 71.968 14.985 ;
      RECT MASK 2 72.488 14.945 72.791 14.985 ;
      RECT MASK 2 73.325 14.945 73.628 14.985 ;
      RECT MASK 2 74.148 14.945 74.451 14.985 ;
      RECT MASK 2 74.985 14.945 75.288 14.985 ;
      RECT MASK 2 75.808 14.945 76.111 14.985 ;
      RECT MASK 2 76.645 14.945 76.948 14.985 ;
      RECT MASK 2 77.468 14.945 77.771 14.985 ;
      RECT MASK 2 78.305 14.945 78.608 14.985 ;
      RECT MASK 2 79.128 14.945 79.431 14.985 ;
      RECT MASK 2 79.965 14.945 80.268 14.985 ;
      RECT MASK 2 80.788 14.945 81.091 14.985 ;
      RECT MASK 2 81.625 14.945 81.928 14.985 ;
      RECT MASK 2 82.448 14.945 82.751 14.985 ;
      RECT MASK 2 83.285 14.945 83.588 14.985 ;
      RECT MASK 2 84.108 14.945 84.411 14.985 ;
      RECT MASK 2 84.945 14.945 85.248 14.985 ;
      RECT MASK 2 85.768 14.945 86.071 14.985 ;
      RECT MASK 2 86.605 14.945 86.908 14.985 ;
      RECT MASK 2 87.428 14.945 87.731 14.985 ;
      RECT MASK 2 88.265 14.945 88.568 14.985 ;
      RECT MASK 2 89.088 14.945 89.391 14.985 ;
      RECT MASK 2 89.925 14.945 90.228 14.985 ;
      RECT MASK 2 90.748 14.945 91.051 14.985 ;
      RECT MASK 2 91.585 14.945 91.888 14.985 ;
      RECT MASK 2 92.408 14.945 92.711 14.985 ;
      RECT MASK 2 93.245 14.945 93.548 14.985 ;
      RECT MASK 2 94.068 14.945 94.371 14.985 ;
      RECT MASK 2 94.905 14.945 95.208 14.985 ;
      RECT MASK 2 95.728 14.945 96.031 14.985 ;
      RECT MASK 2 96.565 14.945 96.868 14.985 ;
      RECT MASK 2 97.388 14.945 97.691 14.985 ;
      RECT MASK 2 98.225 14.945 98.528 14.985 ;
      RECT MASK 2 99.048 14.945 99.351 14.985 ;
      RECT MASK 2 99.885 14.945 100.188 14.985 ;
      RECT MASK 2 100.708 14.945 101.011 14.985 ;
      RECT MASK 2 101.545 14.945 101.848 14.985 ;
      RECT MASK 2 102.368 14.945 102.671 14.985 ;
      RECT MASK 2 103.205 14.945 103.508 14.985 ;
      RECT MASK 2 104.028 14.945 104.331 14.985 ;
      RECT MASK 2 104.865 14.945 105.168 14.985 ;
      RECT MASK 2 105.688 14.945 105.991 14.985 ;
      RECT MASK 2 106.525 14.945 106.828 14.985 ;
      RECT MASK 2 107.348 14.945 107.651 14.985 ;
      RECT MASK 2 108.185 14.945 108.488 14.985 ;
      RECT MASK 2 109.008 14.945 109.311 14.985 ;
      RECT MASK 2 109.845 14.945 110.148 14.985 ;
      RECT MASK 2 110.668 14.945 110.971 14.985 ;
      RECT MASK 2 4.327 15.0175 4.507 15.0575 ;
      RECT MASK 2 111.563 15.0175 111.743 15.0575 ;
      RECT MASK 2 5.163 15.112 5.585 15.152 ;
      RECT MASK 2 5.739 15.112 6.161 15.152 ;
      RECT MASK 2 6.823 15.112 7.245 15.152 ;
      RECT MASK 2 7.399 15.112 7.821 15.152 ;
      RECT MASK 2 8.483 15.112 8.905 15.152 ;
      RECT MASK 2 9.059 15.112 9.481 15.152 ;
      RECT MASK 2 10.143 15.112 10.565 15.152 ;
      RECT MASK 2 10.719 15.112 11.141 15.152 ;
      RECT MASK 2 11.803 15.112 12.225 15.152 ;
      RECT MASK 2 12.379 15.112 12.801 15.152 ;
      RECT MASK 2 13.463 15.112 13.885 15.152 ;
      RECT MASK 2 14.039 15.112 14.461 15.152 ;
      RECT MASK 2 15.123 15.112 15.545 15.152 ;
      RECT MASK 2 15.699 15.112 16.121 15.152 ;
      RECT MASK 2 16.783 15.112 17.205 15.152 ;
      RECT MASK 2 17.359 15.112 17.781 15.152 ;
      RECT MASK 2 18.443 15.112 18.865 15.152 ;
      RECT MASK 2 19.019 15.112 19.441 15.152 ;
      RECT MASK 2 20.103 15.112 20.525 15.152 ;
      RECT MASK 2 20.679 15.112 21.101 15.152 ;
      RECT MASK 2 21.763 15.112 22.185 15.152 ;
      RECT MASK 2 22.339 15.112 22.761 15.152 ;
      RECT MASK 2 23.423 15.112 23.845 15.152 ;
      RECT MASK 2 23.999 15.112 24.421 15.152 ;
      RECT MASK 2 25.083 15.112 25.505 15.152 ;
      RECT MASK 2 25.659 15.112 26.081 15.152 ;
      RECT MASK 2 26.743 15.112 27.165 15.152 ;
      RECT MASK 2 27.319 15.112 27.741 15.152 ;
      RECT MASK 2 28.403 15.112 28.825 15.152 ;
      RECT MASK 2 28.979 15.112 29.401 15.152 ;
      RECT MASK 2 30.063 15.112 30.485 15.152 ;
      RECT MASK 2 30.639 15.112 31.061 15.152 ;
      RECT MASK 2 31.723 15.112 32.145 15.152 ;
      RECT MASK 2 32.299 15.112 32.721 15.152 ;
      RECT MASK 2 33.383 15.112 33.805 15.152 ;
      RECT MASK 2 33.959 15.112 34.381 15.152 ;
      RECT MASK 2 35.043 15.112 35.465 15.152 ;
      RECT MASK 2 35.619 15.112 36.041 15.152 ;
      RECT MASK 2 36.703 15.112 37.125 15.152 ;
      RECT MASK 2 37.279 15.112 37.701 15.152 ;
      RECT MASK 2 38.363 15.112 38.785 15.152 ;
      RECT MASK 2 38.939 15.112 39.361 15.152 ;
      RECT MASK 2 40.023 15.112 40.445 15.152 ;
      RECT MASK 2 40.599 15.112 41.021 15.152 ;
      RECT MASK 2 41.683 15.112 42.105 15.152 ;
      RECT MASK 2 42.259 15.112 42.681 15.152 ;
      RECT MASK 2 43.343 15.112 43.765 15.152 ;
      RECT MASK 2 43.919 15.112 44.341 15.152 ;
      RECT MASK 2 45.003 15.112 45.425 15.152 ;
      RECT MASK 2 45.579 15.112 46.001 15.152 ;
      RECT MASK 2 46.663 15.112 47.085 15.152 ;
      RECT MASK 2 47.239 15.112 47.661 15.152 ;
      RECT MASK 2 48.323 15.112 48.745 15.152 ;
      RECT MASK 2 48.899 15.112 49.321 15.152 ;
      RECT MASK 2 49.983 15.112 50.405 15.152 ;
      RECT MASK 2 50.559 15.112 50.981 15.152 ;
      RECT MASK 2 51.643 15.112 52.065 15.152 ;
      RECT MASK 2 52.219 15.112 52.641 15.152 ;
      RECT MASK 2 53.303 15.112 53.725 15.152 ;
      RECT MASK 2 53.879 15.112 54.301 15.152 ;
      RECT MASK 2 54.963 15.112 55.385 15.152 ;
      RECT MASK 2 55.539 15.112 55.961 15.152 ;
      RECT MASK 2 56.789 15.112 57.211 15.152 ;
      RECT MASK 2 57.365 15.112 57.787 15.152 ;
      RECT MASK 2 58.449 15.112 58.871 15.152 ;
      RECT MASK 2 59.025 15.112 59.447 15.152 ;
      RECT MASK 2 60.109 15.112 60.531 15.152 ;
      RECT MASK 2 60.685 15.112 61.107 15.152 ;
      RECT MASK 2 61.769 15.112 62.191 15.152 ;
      RECT MASK 2 62.345 15.112 62.767 15.152 ;
      RECT MASK 2 63.429 15.112 63.851 15.152 ;
      RECT MASK 2 64.005 15.112 64.427 15.152 ;
      RECT MASK 2 65.089 15.112 65.511 15.152 ;
      RECT MASK 2 65.665 15.112 66.087 15.152 ;
      RECT MASK 2 66.749 15.112 67.171 15.152 ;
      RECT MASK 2 67.325 15.112 67.747 15.152 ;
      RECT MASK 2 68.409 15.112 68.831 15.152 ;
      RECT MASK 2 68.985 15.112 69.407 15.152 ;
      RECT MASK 2 70.069 15.112 70.491 15.152 ;
      RECT MASK 2 70.645 15.112 71.067 15.152 ;
      RECT MASK 2 71.729 15.112 72.151 15.152 ;
      RECT MASK 2 72.305 15.112 72.727 15.152 ;
      RECT MASK 2 73.389 15.112 73.811 15.152 ;
      RECT MASK 2 73.965 15.112 74.387 15.152 ;
      RECT MASK 2 75.049 15.112 75.471 15.152 ;
      RECT MASK 2 75.625 15.112 76.047 15.152 ;
      RECT MASK 2 76.709 15.112 77.131 15.152 ;
      RECT MASK 2 77.285 15.112 77.707 15.152 ;
      RECT MASK 2 78.369 15.112 78.791 15.152 ;
      RECT MASK 2 78.945 15.112 79.367 15.152 ;
      RECT MASK 2 80.029 15.112 80.451 15.152 ;
      RECT MASK 2 80.605 15.112 81.027 15.152 ;
      RECT MASK 2 81.689 15.112 82.111 15.152 ;
      RECT MASK 2 82.265 15.112 82.687 15.152 ;
      RECT MASK 2 83.349 15.112 83.771 15.152 ;
      RECT MASK 2 83.925 15.112 84.347 15.152 ;
      RECT MASK 2 85.009 15.112 85.431 15.152 ;
      RECT MASK 2 85.585 15.112 86.007 15.152 ;
      RECT MASK 2 86.669 15.112 87.091 15.152 ;
      RECT MASK 2 87.245 15.112 87.667 15.152 ;
      RECT MASK 2 88.329 15.112 88.751 15.152 ;
      RECT MASK 2 88.905 15.112 89.327 15.152 ;
      RECT MASK 2 89.989 15.112 90.411 15.152 ;
      RECT MASK 2 90.565 15.112 90.987 15.152 ;
      RECT MASK 2 91.649 15.112 92.071 15.152 ;
      RECT MASK 2 92.225 15.112 92.647 15.152 ;
      RECT MASK 2 93.309 15.112 93.731 15.152 ;
      RECT MASK 2 93.885 15.112 94.307 15.152 ;
      RECT MASK 2 94.969 15.112 95.391 15.152 ;
      RECT MASK 2 95.545 15.112 95.967 15.152 ;
      RECT MASK 2 96.629 15.112 97.051 15.152 ;
      RECT MASK 2 97.205 15.112 97.627 15.152 ;
      RECT MASK 2 98.289 15.112 98.711 15.152 ;
      RECT MASK 2 98.865 15.112 99.287 15.152 ;
      RECT MASK 2 99.949 15.112 100.371 15.152 ;
      RECT MASK 2 100.525 15.112 100.947 15.152 ;
      RECT MASK 2 101.609 15.112 102.031 15.152 ;
      RECT MASK 2 102.185 15.112 102.607 15.152 ;
      RECT MASK 2 103.269 15.112 103.691 15.152 ;
      RECT MASK 2 103.845 15.112 104.267 15.152 ;
      RECT MASK 2 104.929 15.112 105.351 15.152 ;
      RECT MASK 2 105.505 15.112 105.927 15.152 ;
      RECT MASK 2 106.589 15.112 107.011 15.152 ;
      RECT MASK 2 107.165 15.112 107.587 15.152 ;
      RECT MASK 2 108.249 15.112 108.671 15.152 ;
      RECT MASK 2 108.825 15.112 109.247 15.152 ;
      RECT MASK 2 109.909 15.112 110.331 15.152 ;
      RECT MASK 2 110.485 15.112 110.907 15.152 ;
      RECT MASK 2 4.251 15.279 111.819 15.319 ;
      RECT MASK 2 116.291 15.57 116.351 16.62 ;
      RECT MASK 2 116.565 15.57 116.625 16.62 ;
      RECT MASK 2 116.839 15.57 116.899 16.62 ;
      RECT MASK 2 117.113 15.57 117.173 16.62 ;
      RECT MASK 2 117.387 15.57 117.447 16.62 ;
      RECT MASK 2 117.661 15.57 117.721 16.62 ;
      RECT MASK 2 117.935 15.57 117.995 16.62 ;
      RECT MASK 2 118.209 15.57 118.269 16.62 ;
      RECT MASK 2 118.483 15.57 118.543 16.62 ;
      RECT MASK 2 118.757 15.57 118.817 16.62 ;
      RECT MASK 2 119.031 15.57 119.091 16.62 ;
      RECT MASK 2 119.305 15.57 119.365 16.62 ;
      RECT MASK 2 119.579 15.57 119.639 16.62 ;
      RECT MASK 2 119.853 15.57 119.913 16.62 ;
      RECT MASK 2 120.127 15.57 120.187 16.62 ;
      RECT MASK 2 120.401 15.57 120.461 16.62 ;
      RECT MASK 2 120.675 15.57 120.735 16.62 ;
      RECT MASK 2 120.949 15.57 121.009 16.62 ;
      RECT MASK 2 121.223 15.57 121.283 16.62 ;
      RECT MASK 2 121.497 15.57 121.557 16.62 ;
      RECT MASK 2 121.771 15.57 121.831 16.62 ;
      RECT MASK 2 122.045 15.57 122.105 16.62 ;
      RECT MASK 2 122.319 15.57 122.379 16.62 ;
      RECT MASK 2 122.593 15.57 122.653 16.62 ;
      RECT MASK 2 122.867 15.57 122.927 16.62 ;
      RECT MASK 2 123.141 15.57 123.201 16.62 ;
      RECT MASK 2 123.415 15.57 123.475 16.62 ;
      RECT MASK 2 123.689 15.57 123.749 16.62 ;
      RECT MASK 2 123.963 15.57 124.023 16.62 ;
      RECT MASK 2 124.237 15.57 124.297 16.62 ;
      RECT MASK 2 124.511 15.57 124.571 16.62 ;
      RECT MASK 2 124.785 15.57 124.845 16.62 ;
      RECT MASK 2 125.059 15.57 125.119 16.62 ;
      RECT MASK 2 125.333 15.57 125.393 16.62 ;
      RECT MASK 2 125.607 15.57 125.667 16.62 ;
      RECT MASK 2 125.881 15.57 125.941 16.62 ;
      RECT MASK 2 126.155 15.57 126.215 16.62 ;
      RECT MASK 2 126.429 15.57 126.489 16.62 ;
      RECT MASK 2 126.703 15.57 126.763 16.62 ;
      RECT MASK 2 126.977 15.57 127.037 16.62 ;
      RECT MASK 2 127.251 15.57 127.311 16.62 ;
      RECT MASK 2 127.525 15.57 127.585 16.62 ;
      RECT MASK 2 127.799 15.57 127.859 16.62 ;
      RECT MASK 2 128.073 15.57 128.133 16.62 ;
      RECT MASK 2 4.362 15.62 111.708 15.66 ;
      RECT MASK 2 4.362 15.78 111.708 15.82 ;
      RECT MASK 2 4.251 16.121 111.819 16.161 ;
      RECT MASK 2 5.163 16.288 5.585 16.328 ;
      RECT MASK 2 5.739 16.288 6.161 16.328 ;
      RECT MASK 2 6.823 16.288 7.245 16.328 ;
      RECT MASK 2 7.399 16.288 7.821 16.328 ;
      RECT MASK 2 8.483 16.288 8.905 16.328 ;
      RECT MASK 2 9.059 16.288 9.481 16.328 ;
      RECT MASK 2 10.143 16.288 10.565 16.328 ;
      RECT MASK 2 10.719 16.288 11.141 16.328 ;
      RECT MASK 2 11.803 16.288 12.225 16.328 ;
      RECT MASK 2 12.379 16.288 12.801 16.328 ;
      RECT MASK 2 13.463 16.288 13.885 16.328 ;
      RECT MASK 2 14.039 16.288 14.461 16.328 ;
      RECT MASK 2 15.123 16.288 15.545 16.328 ;
      RECT MASK 2 15.699 16.288 16.121 16.328 ;
      RECT MASK 2 16.783 16.288 17.205 16.328 ;
      RECT MASK 2 17.359 16.288 17.781 16.328 ;
      RECT MASK 2 18.443 16.288 18.865 16.328 ;
      RECT MASK 2 19.019 16.288 19.441 16.328 ;
      RECT MASK 2 20.103 16.288 20.525 16.328 ;
      RECT MASK 2 20.679 16.288 21.101 16.328 ;
      RECT MASK 2 21.763 16.288 22.185 16.328 ;
      RECT MASK 2 22.339 16.288 22.761 16.328 ;
      RECT MASK 2 23.423 16.288 23.845 16.328 ;
      RECT MASK 2 23.999 16.288 24.421 16.328 ;
      RECT MASK 2 25.083 16.288 25.505 16.328 ;
      RECT MASK 2 25.659 16.288 26.081 16.328 ;
      RECT MASK 2 26.743 16.288 27.165 16.328 ;
      RECT MASK 2 27.319 16.288 27.741 16.328 ;
      RECT MASK 2 28.403 16.288 28.825 16.328 ;
      RECT MASK 2 28.979 16.288 29.401 16.328 ;
      RECT MASK 2 30.063 16.288 30.485 16.328 ;
      RECT MASK 2 30.639 16.288 31.061 16.328 ;
      RECT MASK 2 31.723 16.288 32.145 16.328 ;
      RECT MASK 2 32.299 16.288 32.721 16.328 ;
      RECT MASK 2 33.383 16.288 33.805 16.328 ;
      RECT MASK 2 33.959 16.288 34.381 16.328 ;
      RECT MASK 2 35.043 16.288 35.465 16.328 ;
      RECT MASK 2 35.619 16.288 36.041 16.328 ;
      RECT MASK 2 36.703 16.288 37.125 16.328 ;
      RECT MASK 2 37.279 16.288 37.701 16.328 ;
      RECT MASK 2 38.363 16.288 38.785 16.328 ;
      RECT MASK 2 38.939 16.288 39.361 16.328 ;
      RECT MASK 2 40.023 16.288 40.445 16.328 ;
      RECT MASK 2 40.599 16.288 41.021 16.328 ;
      RECT MASK 2 41.683 16.288 42.105 16.328 ;
      RECT MASK 2 42.259 16.288 42.681 16.328 ;
      RECT MASK 2 43.343 16.288 43.765 16.328 ;
      RECT MASK 2 43.919 16.288 44.341 16.328 ;
      RECT MASK 2 45.003 16.288 45.425 16.328 ;
      RECT MASK 2 45.579 16.288 46.001 16.328 ;
      RECT MASK 2 46.663 16.288 47.085 16.328 ;
      RECT MASK 2 47.239 16.288 47.661 16.328 ;
      RECT MASK 2 48.323 16.288 48.745 16.328 ;
      RECT MASK 2 48.899 16.288 49.321 16.328 ;
      RECT MASK 2 49.983 16.288 50.405 16.328 ;
      RECT MASK 2 50.559 16.288 50.981 16.328 ;
      RECT MASK 2 51.643 16.288 52.065 16.328 ;
      RECT MASK 2 52.219 16.288 52.641 16.328 ;
      RECT MASK 2 53.303 16.288 53.725 16.328 ;
      RECT MASK 2 53.879 16.288 54.301 16.328 ;
      RECT MASK 2 54.963 16.288 55.385 16.328 ;
      RECT MASK 2 55.539 16.288 55.961 16.328 ;
      RECT MASK 2 56.789 16.288 57.211 16.328 ;
      RECT MASK 2 57.365 16.288 57.787 16.328 ;
      RECT MASK 2 58.449 16.288 58.871 16.328 ;
      RECT MASK 2 59.025 16.288 59.447 16.328 ;
      RECT MASK 2 60.109 16.288 60.531 16.328 ;
      RECT MASK 2 60.685 16.288 61.107 16.328 ;
      RECT MASK 2 61.769 16.288 62.191 16.328 ;
      RECT MASK 2 62.345 16.288 62.767 16.328 ;
      RECT MASK 2 63.429 16.288 63.851 16.328 ;
      RECT MASK 2 64.005 16.288 64.427 16.328 ;
      RECT MASK 2 65.089 16.288 65.511 16.328 ;
      RECT MASK 2 65.665 16.288 66.087 16.328 ;
      RECT MASK 2 66.749 16.288 67.171 16.328 ;
      RECT MASK 2 67.325 16.288 67.747 16.328 ;
      RECT MASK 2 68.409 16.288 68.831 16.328 ;
      RECT MASK 2 68.985 16.288 69.407 16.328 ;
      RECT MASK 2 70.069 16.288 70.491 16.328 ;
      RECT MASK 2 70.645 16.288 71.067 16.328 ;
      RECT MASK 2 71.729 16.288 72.151 16.328 ;
      RECT MASK 2 72.305 16.288 72.727 16.328 ;
      RECT MASK 2 73.389 16.288 73.811 16.328 ;
      RECT MASK 2 73.965 16.288 74.387 16.328 ;
      RECT MASK 2 75.049 16.288 75.471 16.328 ;
      RECT MASK 2 75.625 16.288 76.047 16.328 ;
      RECT MASK 2 76.709 16.288 77.131 16.328 ;
      RECT MASK 2 77.285 16.288 77.707 16.328 ;
      RECT MASK 2 78.369 16.288 78.791 16.328 ;
      RECT MASK 2 78.945 16.288 79.367 16.328 ;
      RECT MASK 2 80.029 16.288 80.451 16.328 ;
      RECT MASK 2 80.605 16.288 81.027 16.328 ;
      RECT MASK 2 81.689 16.288 82.111 16.328 ;
      RECT MASK 2 82.265 16.288 82.687 16.328 ;
      RECT MASK 2 83.349 16.288 83.771 16.328 ;
      RECT MASK 2 83.925 16.288 84.347 16.328 ;
      RECT MASK 2 85.009 16.288 85.431 16.328 ;
      RECT MASK 2 85.585 16.288 86.007 16.328 ;
      RECT MASK 2 86.669 16.288 87.091 16.328 ;
      RECT MASK 2 87.245 16.288 87.667 16.328 ;
      RECT MASK 2 88.329 16.288 88.751 16.328 ;
      RECT MASK 2 88.905 16.288 89.327 16.328 ;
      RECT MASK 2 89.989 16.288 90.411 16.328 ;
      RECT MASK 2 90.565 16.288 90.987 16.328 ;
      RECT MASK 2 91.649 16.288 92.071 16.328 ;
      RECT MASK 2 92.225 16.288 92.647 16.328 ;
      RECT MASK 2 93.309 16.288 93.731 16.328 ;
      RECT MASK 2 93.885 16.288 94.307 16.328 ;
      RECT MASK 2 94.969 16.288 95.391 16.328 ;
      RECT MASK 2 95.545 16.288 95.967 16.328 ;
      RECT MASK 2 96.629 16.288 97.051 16.328 ;
      RECT MASK 2 97.205 16.288 97.627 16.328 ;
      RECT MASK 2 98.289 16.288 98.711 16.328 ;
      RECT MASK 2 98.865 16.288 99.287 16.328 ;
      RECT MASK 2 99.949 16.288 100.371 16.328 ;
      RECT MASK 2 100.525 16.288 100.947 16.328 ;
      RECT MASK 2 101.609 16.288 102.031 16.328 ;
      RECT MASK 2 102.185 16.288 102.607 16.328 ;
      RECT MASK 2 103.269 16.288 103.691 16.328 ;
      RECT MASK 2 103.845 16.288 104.267 16.328 ;
      RECT MASK 2 104.929 16.288 105.351 16.328 ;
      RECT MASK 2 105.505 16.288 105.927 16.328 ;
      RECT MASK 2 106.589 16.288 107.011 16.328 ;
      RECT MASK 2 107.165 16.288 107.587 16.328 ;
      RECT MASK 2 108.249 16.288 108.671 16.328 ;
      RECT MASK 2 108.825 16.288 109.247 16.328 ;
      RECT MASK 2 109.909 16.288 110.331 16.328 ;
      RECT MASK 2 110.485 16.288 110.907 16.328 ;
      RECT MASK 2 4.327 16.3825 4.507 16.4225 ;
      RECT MASK 2 111.563 16.3825 111.743 16.4225 ;
      RECT MASK 2 5.099 16.455 5.402 16.495 ;
      RECT MASK 2 5.922 16.455 6.225 16.495 ;
      RECT MASK 2 6.759 16.455 7.062 16.495 ;
      RECT MASK 2 7.582 16.455 7.885 16.495 ;
      RECT MASK 2 8.419 16.455 8.722 16.495 ;
      RECT MASK 2 9.242 16.455 9.545 16.495 ;
      RECT MASK 2 10.079 16.455 10.382 16.495 ;
      RECT MASK 2 10.902 16.455 11.205 16.495 ;
      RECT MASK 2 11.739 16.455 12.042 16.495 ;
      RECT MASK 2 12.562 16.455 12.865 16.495 ;
      RECT MASK 2 13.399 16.455 13.702 16.495 ;
      RECT MASK 2 14.222 16.455 14.525 16.495 ;
      RECT MASK 2 15.059 16.455 15.362 16.495 ;
      RECT MASK 2 15.882 16.455 16.185 16.495 ;
      RECT MASK 2 16.719 16.455 17.022 16.495 ;
      RECT MASK 2 17.542 16.455 17.845 16.495 ;
      RECT MASK 2 18.379 16.455 18.682 16.495 ;
      RECT MASK 2 19.202 16.455 19.505 16.495 ;
      RECT MASK 2 20.039 16.455 20.342 16.495 ;
      RECT MASK 2 20.862 16.455 21.165 16.495 ;
      RECT MASK 2 21.699 16.455 22.002 16.495 ;
      RECT MASK 2 22.522 16.455 22.825 16.495 ;
      RECT MASK 2 23.359 16.455 23.662 16.495 ;
      RECT MASK 2 24.182 16.455 24.485 16.495 ;
      RECT MASK 2 25.019 16.455 25.322 16.495 ;
      RECT MASK 2 25.842 16.455 26.145 16.495 ;
      RECT MASK 2 26.679 16.455 26.982 16.495 ;
      RECT MASK 2 27.502 16.455 27.805 16.495 ;
      RECT MASK 2 28.339 16.455 28.642 16.495 ;
      RECT MASK 2 29.162 16.455 29.465 16.495 ;
      RECT MASK 2 29.999 16.455 30.302 16.495 ;
      RECT MASK 2 30.822 16.455 31.125 16.495 ;
      RECT MASK 2 31.659 16.455 31.962 16.495 ;
      RECT MASK 2 32.482 16.455 32.785 16.495 ;
      RECT MASK 2 33.319 16.455 33.622 16.495 ;
      RECT MASK 2 34.142 16.455 34.445 16.495 ;
      RECT MASK 2 34.979 16.455 35.282 16.495 ;
      RECT MASK 2 35.802 16.455 36.105 16.495 ;
      RECT MASK 2 36.639 16.455 36.942 16.495 ;
      RECT MASK 2 37.462 16.455 37.765 16.495 ;
      RECT MASK 2 38.299 16.455 38.602 16.495 ;
      RECT MASK 2 39.122 16.455 39.425 16.495 ;
      RECT MASK 2 39.959 16.455 40.262 16.495 ;
      RECT MASK 2 40.782 16.455 41.085 16.495 ;
      RECT MASK 2 41.619 16.455 41.922 16.495 ;
      RECT MASK 2 42.442 16.455 42.745 16.495 ;
      RECT MASK 2 43.279 16.455 43.582 16.495 ;
      RECT MASK 2 44.102 16.455 44.405 16.495 ;
      RECT MASK 2 44.939 16.455 45.242 16.495 ;
      RECT MASK 2 45.762 16.455 46.065 16.495 ;
      RECT MASK 2 46.599 16.455 46.902 16.495 ;
      RECT MASK 2 47.422 16.455 47.725 16.495 ;
      RECT MASK 2 48.259 16.455 48.562 16.495 ;
      RECT MASK 2 49.082 16.455 49.385 16.495 ;
      RECT MASK 2 49.919 16.455 50.222 16.495 ;
      RECT MASK 2 50.742 16.455 51.045 16.495 ;
      RECT MASK 2 51.579 16.455 51.882 16.495 ;
      RECT MASK 2 52.402 16.455 52.705 16.495 ;
      RECT MASK 2 53.239 16.455 53.542 16.495 ;
      RECT MASK 2 54.062 16.455 54.365 16.495 ;
      RECT MASK 2 54.899 16.455 55.202 16.495 ;
      RECT MASK 2 55.722 16.455 56.025 16.495 ;
      RECT MASK 2 56.725 16.455 57.028 16.495 ;
      RECT MASK 2 57.548 16.455 57.851 16.495 ;
      RECT MASK 2 58.385 16.455 58.688 16.495 ;
      RECT MASK 2 59.208 16.455 59.511 16.495 ;
      RECT MASK 2 60.045 16.455 60.348 16.495 ;
      RECT MASK 2 60.868 16.455 61.171 16.495 ;
      RECT MASK 2 61.705 16.455 62.008 16.495 ;
      RECT MASK 2 62.528 16.455 62.831 16.495 ;
      RECT MASK 2 63.365 16.455 63.668 16.495 ;
      RECT MASK 2 64.188 16.455 64.491 16.495 ;
      RECT MASK 2 65.025 16.455 65.328 16.495 ;
      RECT MASK 2 65.848 16.455 66.151 16.495 ;
      RECT MASK 2 66.685 16.455 66.988 16.495 ;
      RECT MASK 2 67.508 16.455 67.811 16.495 ;
      RECT MASK 2 68.345 16.455 68.648 16.495 ;
      RECT MASK 2 69.168 16.455 69.471 16.495 ;
      RECT MASK 2 70.005 16.455 70.308 16.495 ;
      RECT MASK 2 70.828 16.455 71.131 16.495 ;
      RECT MASK 2 71.665 16.455 71.968 16.495 ;
      RECT MASK 2 72.488 16.455 72.791 16.495 ;
      RECT MASK 2 73.325 16.455 73.628 16.495 ;
      RECT MASK 2 74.148 16.455 74.451 16.495 ;
      RECT MASK 2 74.985 16.455 75.288 16.495 ;
      RECT MASK 2 75.808 16.455 76.111 16.495 ;
      RECT MASK 2 76.645 16.455 76.948 16.495 ;
      RECT MASK 2 77.468 16.455 77.771 16.495 ;
      RECT MASK 2 78.305 16.455 78.608 16.495 ;
      RECT MASK 2 79.128 16.455 79.431 16.495 ;
      RECT MASK 2 79.965 16.455 80.268 16.495 ;
      RECT MASK 2 80.788 16.455 81.091 16.495 ;
      RECT MASK 2 81.625 16.455 81.928 16.495 ;
      RECT MASK 2 82.448 16.455 82.751 16.495 ;
      RECT MASK 2 83.285 16.455 83.588 16.495 ;
      RECT MASK 2 84.108 16.455 84.411 16.495 ;
      RECT MASK 2 84.945 16.455 85.248 16.495 ;
      RECT MASK 2 85.768 16.455 86.071 16.495 ;
      RECT MASK 2 86.605 16.455 86.908 16.495 ;
      RECT MASK 2 87.428 16.455 87.731 16.495 ;
      RECT MASK 2 88.265 16.455 88.568 16.495 ;
      RECT MASK 2 89.088 16.455 89.391 16.495 ;
      RECT MASK 2 89.925 16.455 90.228 16.495 ;
      RECT MASK 2 90.748 16.455 91.051 16.495 ;
      RECT MASK 2 91.585 16.455 91.888 16.495 ;
      RECT MASK 2 92.408 16.455 92.711 16.495 ;
      RECT MASK 2 93.245 16.455 93.548 16.495 ;
      RECT MASK 2 94.068 16.455 94.371 16.495 ;
      RECT MASK 2 94.905 16.455 95.208 16.495 ;
      RECT MASK 2 95.728 16.455 96.031 16.495 ;
      RECT MASK 2 96.565 16.455 96.868 16.495 ;
      RECT MASK 2 97.388 16.455 97.691 16.495 ;
      RECT MASK 2 98.225 16.455 98.528 16.495 ;
      RECT MASK 2 99.048 16.455 99.351 16.495 ;
      RECT MASK 2 99.885 16.455 100.188 16.495 ;
      RECT MASK 2 100.708 16.455 101.011 16.495 ;
      RECT MASK 2 101.545 16.455 101.848 16.495 ;
      RECT MASK 2 102.368 16.455 102.671 16.495 ;
      RECT MASK 2 103.205 16.455 103.508 16.495 ;
      RECT MASK 2 104.028 16.455 104.331 16.495 ;
      RECT MASK 2 104.865 16.455 105.168 16.495 ;
      RECT MASK 2 105.688 16.455 105.991 16.495 ;
      RECT MASK 2 106.525 16.455 106.828 16.495 ;
      RECT MASK 2 107.348 16.455 107.651 16.495 ;
      RECT MASK 2 108.185 16.455 108.488 16.495 ;
      RECT MASK 2 109.008 16.455 109.311 16.495 ;
      RECT MASK 2 109.845 16.455 110.148 16.495 ;
      RECT MASK 2 110.668 16.455 110.971 16.495 ;
      RECT MASK 2 5.082 16.865 5.401 16.905 ;
      RECT MASK 2 5.923 16.865 6.242 16.905 ;
      RECT MASK 2 6.742 16.865 7.061 16.905 ;
      RECT MASK 2 7.583 16.865 7.902 16.905 ;
      RECT MASK 2 8.402 16.865 8.721 16.905 ;
      RECT MASK 2 9.243 16.865 9.562 16.905 ;
      RECT MASK 2 10.062 16.865 10.381 16.905 ;
      RECT MASK 2 10.903 16.865 11.222 16.905 ;
      RECT MASK 2 11.722 16.865 12.041 16.905 ;
      RECT MASK 2 12.563 16.865 12.882 16.905 ;
      RECT MASK 2 13.382 16.865 13.701 16.905 ;
      RECT MASK 2 14.223 16.865 14.542 16.905 ;
      RECT MASK 2 15.042 16.865 15.361 16.905 ;
      RECT MASK 2 15.883 16.865 16.202 16.905 ;
      RECT MASK 2 16.702 16.865 17.021 16.905 ;
      RECT MASK 2 17.543 16.865 17.862 16.905 ;
      RECT MASK 2 18.362 16.865 18.681 16.905 ;
      RECT MASK 2 19.203 16.865 19.522 16.905 ;
      RECT MASK 2 20.022 16.865 20.341 16.905 ;
      RECT MASK 2 20.863 16.865 21.182 16.905 ;
      RECT MASK 2 21.682 16.865 22.001 16.905 ;
      RECT MASK 2 22.523 16.865 22.842 16.905 ;
      RECT MASK 2 23.342 16.865 23.661 16.905 ;
      RECT MASK 2 24.183 16.865 24.502 16.905 ;
      RECT MASK 2 25.002 16.865 25.321 16.905 ;
      RECT MASK 2 25.843 16.865 26.162 16.905 ;
      RECT MASK 2 26.662 16.865 26.981 16.905 ;
      RECT MASK 2 27.503 16.865 27.822 16.905 ;
      RECT MASK 2 28.322 16.865 28.641 16.905 ;
      RECT MASK 2 29.163 16.865 29.482 16.905 ;
      RECT MASK 2 29.982 16.865 30.301 16.905 ;
      RECT MASK 2 30.823 16.865 31.142 16.905 ;
      RECT MASK 2 31.642 16.865 31.961 16.905 ;
      RECT MASK 2 32.483 16.865 32.802 16.905 ;
      RECT MASK 2 33.302 16.865 33.621 16.905 ;
      RECT MASK 2 34.143 16.865 34.462 16.905 ;
      RECT MASK 2 34.962 16.865 35.281 16.905 ;
      RECT MASK 2 35.803 16.865 36.122 16.905 ;
      RECT MASK 2 36.622 16.865 36.941 16.905 ;
      RECT MASK 2 37.463 16.865 37.782 16.905 ;
      RECT MASK 2 38.282 16.865 38.601 16.905 ;
      RECT MASK 2 39.123 16.865 39.442 16.905 ;
      RECT MASK 2 39.942 16.865 40.261 16.905 ;
      RECT MASK 2 40.783 16.865 41.102 16.905 ;
      RECT MASK 2 41.602 16.865 41.921 16.905 ;
      RECT MASK 2 42.443 16.865 42.762 16.905 ;
      RECT MASK 2 43.262 16.865 43.581 16.905 ;
      RECT MASK 2 44.103 16.865 44.422 16.905 ;
      RECT MASK 2 44.922 16.865 45.241 16.905 ;
      RECT MASK 2 45.763 16.865 46.082 16.905 ;
      RECT MASK 2 46.582 16.865 46.901 16.905 ;
      RECT MASK 2 47.423 16.865 47.742 16.905 ;
      RECT MASK 2 48.242 16.865 48.561 16.905 ;
      RECT MASK 2 49.083 16.865 49.402 16.905 ;
      RECT MASK 2 49.902 16.865 50.221 16.905 ;
      RECT MASK 2 50.743 16.865 51.062 16.905 ;
      RECT MASK 2 51.562 16.865 51.881 16.905 ;
      RECT MASK 2 52.403 16.865 52.722 16.905 ;
      RECT MASK 2 53.222 16.865 53.541 16.905 ;
      RECT MASK 2 54.063 16.865 54.382 16.905 ;
      RECT MASK 2 54.882 16.865 55.201 16.905 ;
      RECT MASK 2 55.723 16.865 56.042 16.905 ;
      RECT MASK 2 56.708 16.865 57.027 16.905 ;
      RECT MASK 2 57.549 16.865 57.868 16.905 ;
      RECT MASK 2 58.368 16.865 58.687 16.905 ;
      RECT MASK 2 59.209 16.865 59.528 16.905 ;
      RECT MASK 2 60.028 16.865 60.347 16.905 ;
      RECT MASK 2 60.869 16.865 61.188 16.905 ;
      RECT MASK 2 61.688 16.865 62.007 16.905 ;
      RECT MASK 2 62.529 16.865 62.848 16.905 ;
      RECT MASK 2 63.348 16.865 63.667 16.905 ;
      RECT MASK 2 64.189 16.865 64.508 16.905 ;
      RECT MASK 2 65.008 16.865 65.327 16.905 ;
      RECT MASK 2 65.849 16.865 66.168 16.905 ;
      RECT MASK 2 66.668 16.865 66.987 16.905 ;
      RECT MASK 2 67.509 16.865 67.828 16.905 ;
      RECT MASK 2 68.328 16.865 68.647 16.905 ;
      RECT MASK 2 69.169 16.865 69.488 16.905 ;
      RECT MASK 2 69.988 16.865 70.307 16.905 ;
      RECT MASK 2 70.829 16.865 71.148 16.905 ;
      RECT MASK 2 71.648 16.865 71.967 16.905 ;
      RECT MASK 2 72.489 16.865 72.808 16.905 ;
      RECT MASK 2 73.308 16.865 73.627 16.905 ;
      RECT MASK 2 74.149 16.865 74.468 16.905 ;
      RECT MASK 2 74.968 16.865 75.287 16.905 ;
      RECT MASK 2 75.809 16.865 76.128 16.905 ;
      RECT MASK 2 76.628 16.865 76.947 16.905 ;
      RECT MASK 2 77.469 16.865 77.788 16.905 ;
      RECT MASK 2 78.288 16.865 78.607 16.905 ;
      RECT MASK 2 79.129 16.865 79.448 16.905 ;
      RECT MASK 2 79.948 16.865 80.267 16.905 ;
      RECT MASK 2 80.789 16.865 81.108 16.905 ;
      RECT MASK 2 81.608 16.865 81.927 16.905 ;
      RECT MASK 2 82.449 16.865 82.768 16.905 ;
      RECT MASK 2 83.268 16.865 83.587 16.905 ;
      RECT MASK 2 84.109 16.865 84.428 16.905 ;
      RECT MASK 2 84.928 16.865 85.247 16.905 ;
      RECT MASK 2 85.769 16.865 86.088 16.905 ;
      RECT MASK 2 86.588 16.865 86.907 16.905 ;
      RECT MASK 2 87.429 16.865 87.748 16.905 ;
      RECT MASK 2 88.248 16.865 88.567 16.905 ;
      RECT MASK 2 89.089 16.865 89.408 16.905 ;
      RECT MASK 2 89.908 16.865 90.227 16.905 ;
      RECT MASK 2 90.749 16.865 91.068 16.905 ;
      RECT MASK 2 91.568 16.865 91.887 16.905 ;
      RECT MASK 2 92.409 16.865 92.728 16.905 ;
      RECT MASK 2 93.228 16.865 93.547 16.905 ;
      RECT MASK 2 94.069 16.865 94.388 16.905 ;
      RECT MASK 2 94.888 16.865 95.207 16.905 ;
      RECT MASK 2 95.729 16.865 96.048 16.905 ;
      RECT MASK 2 96.548 16.865 96.867 16.905 ;
      RECT MASK 2 97.389 16.865 97.708 16.905 ;
      RECT MASK 2 98.208 16.865 98.527 16.905 ;
      RECT MASK 2 99.049 16.865 99.368 16.905 ;
      RECT MASK 2 99.868 16.865 100.187 16.905 ;
      RECT MASK 2 100.709 16.865 101.028 16.905 ;
      RECT MASK 2 101.528 16.865 101.847 16.905 ;
      RECT MASK 2 102.369 16.865 102.688 16.905 ;
      RECT MASK 2 103.188 16.865 103.507 16.905 ;
      RECT MASK 2 104.029 16.865 104.348 16.905 ;
      RECT MASK 2 104.848 16.865 105.167 16.905 ;
      RECT MASK 2 105.689 16.865 106.008 16.905 ;
      RECT MASK 2 106.508 16.865 106.827 16.905 ;
      RECT MASK 2 107.349 16.865 107.668 16.905 ;
      RECT MASK 2 108.168 16.865 108.487 16.905 ;
      RECT MASK 2 109.009 16.865 109.328 16.905 ;
      RECT MASK 2 109.828 16.865 110.147 16.905 ;
      RECT MASK 2 110.669 16.865 110.988 16.905 ;
      RECT MASK 2 4.327 16.9375 4.507 16.9775 ;
      RECT MASK 2 111.563 16.9375 111.743 16.9775 ;
      RECT MASK 2 5.036 17.032 5.586 17.072 ;
      RECT MASK 2 5.738 17.032 6.288 17.072 ;
      RECT MASK 2 6.696 17.032 7.246 17.072 ;
      RECT MASK 2 7.398 17.032 7.948 17.072 ;
      RECT MASK 2 8.356 17.032 8.906 17.072 ;
      RECT MASK 2 9.058 17.032 9.608 17.072 ;
      RECT MASK 2 10.016 17.032 10.566 17.072 ;
      RECT MASK 2 10.718 17.032 11.268 17.072 ;
      RECT MASK 2 11.676 17.032 12.226 17.072 ;
      RECT MASK 2 12.378 17.032 12.928 17.072 ;
      RECT MASK 2 13.336 17.032 13.886 17.072 ;
      RECT MASK 2 14.038 17.032 14.588 17.072 ;
      RECT MASK 2 14.996 17.032 15.546 17.072 ;
      RECT MASK 2 15.698 17.032 16.248 17.072 ;
      RECT MASK 2 16.656 17.032 17.206 17.072 ;
      RECT MASK 2 17.358 17.032 17.908 17.072 ;
      RECT MASK 2 18.316 17.032 18.866 17.072 ;
      RECT MASK 2 19.018 17.032 19.568 17.072 ;
      RECT MASK 2 19.976 17.032 20.526 17.072 ;
      RECT MASK 2 20.678 17.032 21.228 17.072 ;
      RECT MASK 2 21.636 17.032 22.186 17.072 ;
      RECT MASK 2 22.338 17.032 22.888 17.072 ;
      RECT MASK 2 23.296 17.032 23.846 17.072 ;
      RECT MASK 2 23.998 17.032 24.548 17.072 ;
      RECT MASK 2 24.956 17.032 25.506 17.072 ;
      RECT MASK 2 25.658 17.032 26.208 17.072 ;
      RECT MASK 2 26.616 17.032 27.166 17.072 ;
      RECT MASK 2 27.318 17.032 27.868 17.072 ;
      RECT MASK 2 28.276 17.032 28.826 17.072 ;
      RECT MASK 2 28.978 17.032 29.528 17.072 ;
      RECT MASK 2 29.936 17.032 30.486 17.072 ;
      RECT MASK 2 30.638 17.032 31.188 17.072 ;
      RECT MASK 2 31.596 17.032 32.146 17.072 ;
      RECT MASK 2 32.298 17.032 32.848 17.072 ;
      RECT MASK 2 33.256 17.032 33.806 17.072 ;
      RECT MASK 2 33.958 17.032 34.508 17.072 ;
      RECT MASK 2 34.916 17.032 35.466 17.072 ;
      RECT MASK 2 35.618 17.032 36.168 17.072 ;
      RECT MASK 2 36.576 17.032 37.126 17.072 ;
      RECT MASK 2 37.278 17.032 37.828 17.072 ;
      RECT MASK 2 38.236 17.032 38.786 17.072 ;
      RECT MASK 2 38.938 17.032 39.488 17.072 ;
      RECT MASK 2 39.896 17.032 40.446 17.072 ;
      RECT MASK 2 40.598 17.032 41.148 17.072 ;
      RECT MASK 2 41.556 17.032 42.106 17.072 ;
      RECT MASK 2 42.258 17.032 42.808 17.072 ;
      RECT MASK 2 43.216 17.032 43.766 17.072 ;
      RECT MASK 2 43.918 17.032 44.468 17.072 ;
      RECT MASK 2 44.876 17.032 45.426 17.072 ;
      RECT MASK 2 45.578 17.032 46.128 17.072 ;
      RECT MASK 2 46.536 17.032 47.086 17.072 ;
      RECT MASK 2 47.238 17.032 47.788 17.072 ;
      RECT MASK 2 48.196 17.032 48.746 17.072 ;
      RECT MASK 2 48.898 17.032 49.448 17.072 ;
      RECT MASK 2 49.856 17.032 50.406 17.072 ;
      RECT MASK 2 50.558 17.032 51.108 17.072 ;
      RECT MASK 2 51.516 17.032 52.066 17.072 ;
      RECT MASK 2 52.218 17.032 52.768 17.072 ;
      RECT MASK 2 53.176 17.032 53.726 17.072 ;
      RECT MASK 2 53.878 17.032 54.428 17.072 ;
      RECT MASK 2 54.836 17.032 55.386 17.072 ;
      RECT MASK 2 55.538 17.032 56.088 17.072 ;
      RECT MASK 2 56.662 17.032 57.212 17.072 ;
      RECT MASK 2 57.364 17.032 57.914 17.072 ;
      RECT MASK 2 58.322 17.032 58.872 17.072 ;
      RECT MASK 2 59.024 17.032 59.574 17.072 ;
      RECT MASK 2 59.982 17.032 60.532 17.072 ;
      RECT MASK 2 60.684 17.032 61.234 17.072 ;
      RECT MASK 2 61.642 17.032 62.192 17.072 ;
      RECT MASK 2 62.344 17.032 62.894 17.072 ;
      RECT MASK 2 63.302 17.032 63.852 17.072 ;
      RECT MASK 2 64.004 17.032 64.554 17.072 ;
      RECT MASK 2 64.962 17.032 65.512 17.072 ;
      RECT MASK 2 65.664 17.032 66.214 17.072 ;
      RECT MASK 2 66.622 17.032 67.172 17.072 ;
      RECT MASK 2 67.324 17.032 67.874 17.072 ;
      RECT MASK 2 68.282 17.032 68.832 17.072 ;
      RECT MASK 2 68.984 17.032 69.534 17.072 ;
      RECT MASK 2 69.942 17.032 70.492 17.072 ;
      RECT MASK 2 70.644 17.032 71.194 17.072 ;
      RECT MASK 2 71.602 17.032 72.152 17.072 ;
      RECT MASK 2 72.304 17.032 72.854 17.072 ;
      RECT MASK 2 73.262 17.032 73.812 17.072 ;
      RECT MASK 2 73.964 17.032 74.514 17.072 ;
      RECT MASK 2 74.922 17.032 75.472 17.072 ;
      RECT MASK 2 75.624 17.032 76.174 17.072 ;
      RECT MASK 2 76.582 17.032 77.132 17.072 ;
      RECT MASK 2 77.284 17.032 77.834 17.072 ;
      RECT MASK 2 78.242 17.032 78.792 17.072 ;
      RECT MASK 2 78.944 17.032 79.494 17.072 ;
      RECT MASK 2 79.902 17.032 80.452 17.072 ;
      RECT MASK 2 80.604 17.032 81.154 17.072 ;
      RECT MASK 2 81.562 17.032 82.112 17.072 ;
      RECT MASK 2 82.264 17.032 82.814 17.072 ;
      RECT MASK 2 83.222 17.032 83.772 17.072 ;
      RECT MASK 2 83.924 17.032 84.474 17.072 ;
      RECT MASK 2 84.882 17.032 85.432 17.072 ;
      RECT MASK 2 85.584 17.032 86.134 17.072 ;
      RECT MASK 2 86.542 17.032 87.092 17.072 ;
      RECT MASK 2 87.244 17.032 87.794 17.072 ;
      RECT MASK 2 88.202 17.032 88.752 17.072 ;
      RECT MASK 2 88.904 17.032 89.454 17.072 ;
      RECT MASK 2 89.862 17.032 90.412 17.072 ;
      RECT MASK 2 90.564 17.032 91.114 17.072 ;
      RECT MASK 2 91.522 17.032 92.072 17.072 ;
      RECT MASK 2 92.224 17.032 92.774 17.072 ;
      RECT MASK 2 93.182 17.032 93.732 17.072 ;
      RECT MASK 2 93.884 17.032 94.434 17.072 ;
      RECT MASK 2 94.842 17.032 95.392 17.072 ;
      RECT MASK 2 95.544 17.032 96.094 17.072 ;
      RECT MASK 2 96.502 17.032 97.052 17.072 ;
      RECT MASK 2 97.204 17.032 97.754 17.072 ;
      RECT MASK 2 98.162 17.032 98.712 17.072 ;
      RECT MASK 2 98.864 17.032 99.414 17.072 ;
      RECT MASK 2 99.822 17.032 100.372 17.072 ;
      RECT MASK 2 100.524 17.032 101.074 17.072 ;
      RECT MASK 2 101.482 17.032 102.032 17.072 ;
      RECT MASK 2 102.184 17.032 102.734 17.072 ;
      RECT MASK 2 103.142 17.032 103.692 17.072 ;
      RECT MASK 2 103.844 17.032 104.394 17.072 ;
      RECT MASK 2 104.802 17.032 105.352 17.072 ;
      RECT MASK 2 105.504 17.032 106.054 17.072 ;
      RECT MASK 2 106.462 17.032 107.012 17.072 ;
      RECT MASK 2 107.164 17.032 107.714 17.072 ;
      RECT MASK 2 108.122 17.032 108.672 17.072 ;
      RECT MASK 2 108.824 17.032 109.374 17.072 ;
      RECT MASK 2 109.782 17.032 110.332 17.072 ;
      RECT MASK 2 110.484 17.032 111.034 17.072 ;
      RECT MASK 2 4.251 17.199 111.819 17.239 ;
      RECT MASK 2 116.291 17.28 116.351 18.33 ;
      RECT MASK 2 116.565 17.28 116.625 18.33 ;
      RECT MASK 2 116.839 17.28 116.899 18.33 ;
      RECT MASK 2 117.113 17.28 117.173 18.33 ;
      RECT MASK 2 117.387 17.28 117.447 18.33 ;
      RECT MASK 2 117.661 17.28 117.721 18.33 ;
      RECT MASK 2 117.935 17.28 117.995 18.33 ;
      RECT MASK 2 118.209 17.28 118.269 18.33 ;
      RECT MASK 2 118.483 17.28 118.543 18.33 ;
      RECT MASK 2 118.757 17.28 118.817 18.33 ;
      RECT MASK 2 119.031 17.28 119.091 18.33 ;
      RECT MASK 2 119.305 17.28 119.365 18.33 ;
      RECT MASK 2 119.579 17.28 119.639 18.33 ;
      RECT MASK 2 119.853 17.28 119.913 18.33 ;
      RECT MASK 2 120.127 17.28 120.187 18.33 ;
      RECT MASK 2 120.401 17.28 120.461 18.33 ;
      RECT MASK 2 120.675 17.28 120.735 18.33 ;
      RECT MASK 2 120.949 17.28 121.009 18.33 ;
      RECT MASK 2 121.223 17.28 121.283 18.33 ;
      RECT MASK 2 121.497 17.28 121.557 18.33 ;
      RECT MASK 2 121.771 17.28 121.831 18.33 ;
      RECT MASK 2 122.045 17.28 122.105 18.33 ;
      RECT MASK 2 122.319 17.28 122.379 18.33 ;
      RECT MASK 2 122.593 17.28 122.653 18.33 ;
      RECT MASK 2 122.867 17.28 122.927 18.33 ;
      RECT MASK 2 123.141 17.28 123.201 18.33 ;
      RECT MASK 2 123.415 17.28 123.475 18.33 ;
      RECT MASK 2 123.689 17.28 123.749 18.33 ;
      RECT MASK 2 123.963 17.28 124.023 18.33 ;
      RECT MASK 2 124.237 17.28 124.297 18.33 ;
      RECT MASK 2 124.511 17.28 124.571 18.33 ;
      RECT MASK 2 124.785 17.28 124.845 18.33 ;
      RECT MASK 2 125.059 17.28 125.119 18.33 ;
      RECT MASK 2 125.333 17.28 125.393 18.33 ;
      RECT MASK 2 125.607 17.28 125.667 18.33 ;
      RECT MASK 2 125.881 17.28 125.941 18.33 ;
      RECT MASK 2 126.155 17.28 126.215 18.33 ;
      RECT MASK 2 126.429 17.28 126.489 18.33 ;
      RECT MASK 2 126.703 17.28 126.763 18.33 ;
      RECT MASK 2 126.977 17.28 127.037 18.33 ;
      RECT MASK 2 127.251 17.28 127.311 18.33 ;
      RECT MASK 2 127.525 17.28 127.585 18.33 ;
      RECT MASK 2 127.799 17.28 127.859 18.33 ;
      RECT MASK 2 128.073 17.28 128.133 18.33 ;
      RECT MASK 2 4.362 17.54 111.708 17.58 ;
      RECT MASK 2 4.362 17.7 111.708 17.74 ;
      RECT MASK 2 5.062 17.96 109.834 18 ;
      RECT MASK 2 5.062 18.15 109.834 18.19 ;
      RECT MASK 2 5.062 18.491 109.898 18.531 ;
      RECT MASK 2 5.062 18.659 109.898 18.699 ;
      RECT MASK 2 5.816 18.843 5.999 18.883 ;
      RECT MASK 2 6.221 18.843 6.404 18.883 ;
      RECT MASK 2 6.978 18.843 7.161 18.883 ;
      RECT MASK 2 7.383 18.843 7.566 18.883 ;
      RECT MASK 2 8.14 18.843 8.323 18.883 ;
      RECT MASK 2 8.545 18.843 8.728 18.883 ;
      RECT MASK 2 9.302 18.843 9.485 18.883 ;
      RECT MASK 2 9.707 18.843 9.89 18.883 ;
      RECT MASK 2 12.434 18.843 12.617 18.883 ;
      RECT MASK 2 12.839 18.843 13.022 18.883 ;
      RECT MASK 2 13.596 18.843 13.779 18.883 ;
      RECT MASK 2 14.001 18.843 14.184 18.883 ;
      RECT MASK 2 14.758 18.843 14.941 18.883 ;
      RECT MASK 2 15.163 18.843 15.346 18.883 ;
      RECT MASK 2 15.92 18.843 16.103 18.883 ;
      RECT MASK 2 16.325 18.843 16.508 18.883 ;
      RECT MASK 2 19.052 18.843 19.235 18.883 ;
      RECT MASK 2 19.457 18.843 19.64 18.883 ;
      RECT MASK 2 20.214 18.843 20.397 18.883 ;
      RECT MASK 2 20.619 18.843 20.802 18.883 ;
      RECT MASK 2 21.376 18.843 21.559 18.883 ;
      RECT MASK 2 21.781 18.843 21.964 18.883 ;
      RECT MASK 2 22.538 18.843 22.721 18.883 ;
      RECT MASK 2 22.943 18.843 23.126 18.883 ;
      RECT MASK 2 25.67 18.843 25.853 18.883 ;
      RECT MASK 2 26.075 18.843 26.258 18.883 ;
      RECT MASK 2 26.832 18.843 27.015 18.883 ;
      RECT MASK 2 27.237 18.843 27.42 18.883 ;
      RECT MASK 2 27.994 18.843 28.177 18.883 ;
      RECT MASK 2 28.399 18.843 28.582 18.883 ;
      RECT MASK 2 29.156 18.843 29.339 18.883 ;
      RECT MASK 2 29.561 18.843 29.744 18.883 ;
      RECT MASK 2 32.288 18.843 32.471 18.883 ;
      RECT MASK 2 32.693 18.843 32.876 18.883 ;
      RECT MASK 2 33.45 18.843 33.633 18.883 ;
      RECT MASK 2 33.855 18.843 34.038 18.883 ;
      RECT MASK 2 34.612 18.843 34.795 18.883 ;
      RECT MASK 2 35.017 18.843 35.2 18.883 ;
      RECT MASK 2 35.774 18.843 35.957 18.883 ;
      RECT MASK 2 36.179 18.843 36.362 18.883 ;
      RECT MASK 2 38.906 18.843 39.089 18.883 ;
      RECT MASK 2 39.311 18.843 39.494 18.883 ;
      RECT MASK 2 40.068 18.843 40.251 18.883 ;
      RECT MASK 2 40.473 18.843 40.656 18.883 ;
      RECT MASK 2 41.23 18.843 41.413 18.883 ;
      RECT MASK 2 41.635 18.843 41.818 18.883 ;
      RECT MASK 2 42.392 18.843 42.575 18.883 ;
      RECT MASK 2 42.797 18.843 42.98 18.883 ;
      RECT MASK 2 45.524 18.843 45.707 18.883 ;
      RECT MASK 2 45.929 18.843 46.112 18.883 ;
      RECT MASK 2 46.686 18.843 46.869 18.883 ;
      RECT MASK 2 47.091 18.843 47.274 18.883 ;
      RECT MASK 2 47.848 18.843 48.031 18.883 ;
      RECT MASK 2 48.253 18.843 48.436 18.883 ;
      RECT MASK 2 49.01 18.843 49.193 18.883 ;
      RECT MASK 2 49.415 18.843 49.598 18.883 ;
      RECT MASK 2 52.142 18.843 52.325 18.883 ;
      RECT MASK 2 52.547 18.843 52.73 18.883 ;
      RECT MASK 2 53.304 18.843 53.487 18.883 ;
      RECT MASK 2 53.709 18.843 53.892 18.883 ;
      RECT MASK 2 54.466 18.843 54.649 18.883 ;
      RECT MASK 2 54.871 18.843 55.054 18.883 ;
      RECT MASK 2 55.628 18.843 55.811 18.883 ;
      RECT MASK 2 56.033 18.843 56.216 18.883 ;
      RECT MASK 2 58.76 18.843 58.943 18.883 ;
      RECT MASK 2 59.165 18.843 59.348 18.883 ;
      RECT MASK 2 59.922 18.843 60.105 18.883 ;
      RECT MASK 2 60.327 18.843 60.51 18.883 ;
      RECT MASK 2 61.084 18.843 61.267 18.883 ;
      RECT MASK 2 61.489 18.843 61.672 18.883 ;
      RECT MASK 2 62.246 18.843 62.429 18.883 ;
      RECT MASK 2 62.651 18.843 62.834 18.883 ;
      RECT MASK 2 65.378 18.843 65.561 18.883 ;
      RECT MASK 2 65.783 18.843 65.966 18.883 ;
      RECT MASK 2 66.54 18.843 66.723 18.883 ;
      RECT MASK 2 66.945 18.843 67.128 18.883 ;
      RECT MASK 2 67.702 18.843 67.885 18.883 ;
      RECT MASK 2 68.107 18.843 68.29 18.883 ;
      RECT MASK 2 68.864 18.843 69.047 18.883 ;
      RECT MASK 2 69.269 18.843 69.452 18.883 ;
      RECT MASK 2 71.996 18.843 72.179 18.883 ;
      RECT MASK 2 72.401 18.843 72.584 18.883 ;
      RECT MASK 2 73.158 18.843 73.341 18.883 ;
      RECT MASK 2 73.563 18.843 73.746 18.883 ;
      RECT MASK 2 74.32 18.843 74.503 18.883 ;
      RECT MASK 2 74.725 18.843 74.908 18.883 ;
      RECT MASK 2 75.482 18.843 75.665 18.883 ;
      RECT MASK 2 75.887 18.843 76.07 18.883 ;
      RECT MASK 2 78.614 18.843 78.797 18.883 ;
      RECT MASK 2 79.019 18.843 79.202 18.883 ;
      RECT MASK 2 79.776 18.843 79.959 18.883 ;
      RECT MASK 2 80.181 18.843 80.364 18.883 ;
      RECT MASK 2 80.938 18.843 81.121 18.883 ;
      RECT MASK 2 81.343 18.843 81.526 18.883 ;
      RECT MASK 2 82.1 18.843 82.283 18.883 ;
      RECT MASK 2 82.505 18.843 82.688 18.883 ;
      RECT MASK 2 85.232 18.843 85.415 18.883 ;
      RECT MASK 2 85.637 18.843 85.82 18.883 ;
      RECT MASK 2 86.394 18.843 86.577 18.883 ;
      RECT MASK 2 86.799 18.843 86.982 18.883 ;
      RECT MASK 2 87.556 18.843 87.739 18.883 ;
      RECT MASK 2 87.961 18.843 88.144 18.883 ;
      RECT MASK 2 88.718 18.843 88.901 18.883 ;
      RECT MASK 2 89.123 18.843 89.306 18.883 ;
      RECT MASK 2 91.85 18.843 92.033 18.883 ;
      RECT MASK 2 92.255 18.843 92.438 18.883 ;
      RECT MASK 2 93.012 18.843 93.195 18.883 ;
      RECT MASK 2 93.417 18.843 93.6 18.883 ;
      RECT MASK 2 94.174 18.843 94.357 18.883 ;
      RECT MASK 2 94.579 18.843 94.762 18.883 ;
      RECT MASK 2 95.336 18.843 95.519 18.883 ;
      RECT MASK 2 95.741 18.843 95.924 18.883 ;
      RECT MASK 2 98.468 18.843 98.651 18.883 ;
      RECT MASK 2 98.873 18.843 99.056 18.883 ;
      RECT MASK 2 99.63 18.843 99.813 18.883 ;
      RECT MASK 2 100.035 18.843 100.218 18.883 ;
      RECT MASK 2 100.792 18.843 100.975 18.883 ;
      RECT MASK 2 101.197 18.843 101.38 18.883 ;
      RECT MASK 2 101.954 18.843 102.137 18.883 ;
      RECT MASK 2 102.359 18.843 102.542 18.883 ;
      RECT MASK 2 105.086 18.843 105.269 18.883 ;
      RECT MASK 2 105.491 18.843 105.674 18.883 ;
      RECT MASK 2 106.248 18.843 106.431 18.883 ;
      RECT MASK 2 106.653 18.843 106.836 18.883 ;
      RECT MASK 2 107.41 18.843 107.593 18.883 ;
      RECT MASK 2 107.815 18.843 107.998 18.883 ;
      RECT MASK 2 108.572 18.843 108.755 18.883 ;
      RECT MASK 2 108.977 18.843 109.16 18.883 ;
      RECT MASK 2 116.291 18.99 116.351 20.04 ;
      RECT MASK 2 116.565 18.99 116.625 20.04 ;
      RECT MASK 2 116.839 18.99 116.899 20.04 ;
      RECT MASK 2 117.113 18.99 117.173 20.04 ;
      RECT MASK 2 117.387 18.99 117.447 20.04 ;
      RECT MASK 2 117.661 18.99 117.721 20.04 ;
      RECT MASK 2 117.935 18.99 117.995 20.04 ;
      RECT MASK 2 118.209 18.99 118.269 20.04 ;
      RECT MASK 2 118.483 18.99 118.543 20.04 ;
      RECT MASK 2 118.757 18.99 118.817 20.04 ;
      RECT MASK 2 119.031 18.99 119.091 20.04 ;
      RECT MASK 2 119.305 18.99 119.365 20.04 ;
      RECT MASK 2 119.579 18.99 119.639 20.04 ;
      RECT MASK 2 119.853 18.99 119.913 20.04 ;
      RECT MASK 2 120.127 18.99 120.187 20.04 ;
      RECT MASK 2 120.401 18.99 120.461 20.04 ;
      RECT MASK 2 120.675 18.99 120.735 20.04 ;
      RECT MASK 2 120.949 18.99 121.009 20.04 ;
      RECT MASK 2 121.223 18.99 121.283 20.04 ;
      RECT MASK 2 121.497 18.99 121.557 20.04 ;
      RECT MASK 2 121.771 18.99 121.831 20.04 ;
      RECT MASK 2 122.045 18.99 122.105 20.04 ;
      RECT MASK 2 122.319 18.99 122.379 20.04 ;
      RECT MASK 2 122.593 18.99 122.653 20.04 ;
      RECT MASK 2 122.867 18.99 122.927 20.04 ;
      RECT MASK 2 123.141 18.99 123.201 20.04 ;
      RECT MASK 2 123.415 18.99 123.475 20.04 ;
      RECT MASK 2 123.689 18.99 123.749 20.04 ;
      RECT MASK 2 123.963 18.99 124.023 20.04 ;
      RECT MASK 2 124.237 18.99 124.297 20.04 ;
      RECT MASK 2 124.511 18.99 124.571 20.04 ;
      RECT MASK 2 124.785 18.99 124.845 20.04 ;
      RECT MASK 2 125.059 18.99 125.119 20.04 ;
      RECT MASK 2 125.333 18.99 125.393 20.04 ;
      RECT MASK 2 125.607 18.99 125.667 20.04 ;
      RECT MASK 2 125.881 18.99 125.941 20.04 ;
      RECT MASK 2 126.155 18.99 126.215 20.04 ;
      RECT MASK 2 126.429 18.99 126.489 20.04 ;
      RECT MASK 2 126.703 18.99 126.763 20.04 ;
      RECT MASK 2 126.977 18.99 127.037 20.04 ;
      RECT MASK 2 127.251 18.99 127.311 20.04 ;
      RECT MASK 2 127.525 18.99 127.585 20.04 ;
      RECT MASK 2 127.799 18.99 127.859 20.04 ;
      RECT MASK 2 128.073 18.99 128.133 20.04 ;
      RECT MASK 2 5.107 19.065 5.287 19.105 ;
      RECT MASK 2 10.419 19.065 10.599 19.105 ;
      RECT MASK 2 11.725 19.065 11.905 19.105 ;
      RECT MASK 2 17.037 19.065 17.217 19.105 ;
      RECT MASK 2 18.343 19.065 18.523 19.105 ;
      RECT MASK 2 23.655 19.065 23.835 19.105 ;
      RECT MASK 2 24.961 19.065 25.141 19.105 ;
      RECT MASK 2 30.273 19.065 30.453 19.105 ;
      RECT MASK 2 31.579 19.065 31.759 19.105 ;
      RECT MASK 2 36.891 19.065 37.071 19.105 ;
      RECT MASK 2 38.197 19.065 38.377 19.105 ;
      RECT MASK 2 43.509 19.065 43.689 19.105 ;
      RECT MASK 2 44.815 19.065 44.995 19.105 ;
      RECT MASK 2 50.127 19.065 50.307 19.105 ;
      RECT MASK 2 51.433 19.065 51.613 19.105 ;
      RECT MASK 2 56.745 19.065 56.925 19.105 ;
      RECT MASK 2 58.051 19.065 58.231 19.105 ;
      RECT MASK 2 63.363 19.065 63.543 19.105 ;
      RECT MASK 2 64.669 19.065 64.849 19.105 ;
      RECT MASK 2 69.981 19.065 70.161 19.105 ;
      RECT MASK 2 71.287 19.065 71.467 19.105 ;
      RECT MASK 2 76.599 19.065 76.779 19.105 ;
      RECT MASK 2 77.905 19.065 78.085 19.105 ;
      RECT MASK 2 83.217 19.065 83.397 19.105 ;
      RECT MASK 2 84.523 19.065 84.703 19.105 ;
      RECT MASK 2 89.835 19.065 90.015 19.105 ;
      RECT MASK 2 91.141 19.065 91.321 19.105 ;
      RECT MASK 2 96.453 19.065 96.633 19.105 ;
      RECT MASK 2 97.759 19.065 97.939 19.105 ;
      RECT MASK 2 103.071 19.065 103.251 19.105 ;
      RECT MASK 2 104.377 19.065 104.557 19.105 ;
      RECT MASK 2 109.689 19.065 109.869 19.105 ;
      RECT MASK 2 1.406 19.07 4.69 19.11 ;
      RECT MASK 2 1.406 19.26 4.69 19.3 ;
      RECT MASK 2 5.1135 19.475 109.836 19.515 ;
      RECT MASK 2 2.362 19.77 2.422 20.82 ;
      RECT MASK 2 2.636 19.77 2.696 20.82 ;
      RECT MASK 2 2.91 19.77 2.97 20.82 ;
      RECT MASK 2 3.184 19.77 3.244 20.82 ;
      RECT MASK 2 3.458 19.77 3.518 20.82 ;
      RECT MASK 2 3.732 19.77 3.792 20.82 ;
      RECT MASK 2 5.1135 19.995 109.836 20.035 ;
      RECT MASK 2 5.107 20.441 5.287 20.481 ;
      RECT MASK 2 10.419 20.441 10.599 20.481 ;
      RECT MASK 2 11.725 20.441 11.905 20.481 ;
      RECT MASK 2 17.037 20.441 17.217 20.481 ;
      RECT MASK 2 18.343 20.441 18.523 20.481 ;
      RECT MASK 2 23.655 20.441 23.835 20.481 ;
      RECT MASK 2 24.961 20.441 25.141 20.481 ;
      RECT MASK 2 30.273 20.441 30.453 20.481 ;
      RECT MASK 2 31.579 20.441 31.759 20.481 ;
      RECT MASK 2 36.891 20.441 37.071 20.481 ;
      RECT MASK 2 38.197 20.441 38.377 20.481 ;
      RECT MASK 2 43.509 20.441 43.689 20.481 ;
      RECT MASK 2 44.815 20.441 44.995 20.481 ;
      RECT MASK 2 50.127 20.441 50.307 20.481 ;
      RECT MASK 2 51.433 20.441 51.613 20.481 ;
      RECT MASK 2 56.745 20.441 56.925 20.481 ;
      RECT MASK 2 58.051 20.441 58.231 20.481 ;
      RECT MASK 2 63.363 20.441 63.543 20.481 ;
      RECT MASK 2 64.669 20.441 64.849 20.481 ;
      RECT MASK 2 69.981 20.441 70.161 20.481 ;
      RECT MASK 2 71.287 20.441 71.467 20.481 ;
      RECT MASK 2 76.599 20.441 76.779 20.481 ;
      RECT MASK 2 77.905 20.441 78.085 20.481 ;
      RECT MASK 2 83.217 20.441 83.397 20.481 ;
      RECT MASK 2 84.523 20.441 84.703 20.481 ;
      RECT MASK 2 89.835 20.441 90.015 20.481 ;
      RECT MASK 2 91.141 20.441 91.321 20.481 ;
      RECT MASK 2 96.453 20.441 96.633 20.481 ;
      RECT MASK 2 97.759 20.441 97.939 20.481 ;
      RECT MASK 2 103.071 20.441 103.251 20.481 ;
      RECT MASK 2 104.377 20.441 104.557 20.481 ;
      RECT MASK 2 109.689 20.441 109.869 20.481 ;
      RECT MASK 2 5.816 20.627 5.999 20.667 ;
      RECT MASK 2 6.221 20.627 6.404 20.667 ;
      RECT MASK 2 6.978 20.627 7.161 20.667 ;
      RECT MASK 2 7.383 20.627 7.566 20.667 ;
      RECT MASK 2 8.14 20.627 8.323 20.667 ;
      RECT MASK 2 8.545 20.627 8.728 20.667 ;
      RECT MASK 2 9.302 20.627 9.485 20.667 ;
      RECT MASK 2 9.707 20.627 9.89 20.667 ;
      RECT MASK 2 12.434 20.627 12.617 20.667 ;
      RECT MASK 2 12.839 20.627 13.022 20.667 ;
      RECT MASK 2 13.596 20.627 13.779 20.667 ;
      RECT MASK 2 14.001 20.627 14.184 20.667 ;
      RECT MASK 2 14.758 20.627 14.941 20.667 ;
      RECT MASK 2 15.163 20.627 15.346 20.667 ;
      RECT MASK 2 15.92 20.627 16.103 20.667 ;
      RECT MASK 2 16.325 20.627 16.508 20.667 ;
      RECT MASK 2 19.052 20.627 19.235 20.667 ;
      RECT MASK 2 19.457 20.627 19.64 20.667 ;
      RECT MASK 2 20.214 20.627 20.397 20.667 ;
      RECT MASK 2 20.619 20.627 20.802 20.667 ;
      RECT MASK 2 21.376 20.627 21.559 20.667 ;
      RECT MASK 2 21.781 20.627 21.964 20.667 ;
      RECT MASK 2 22.538 20.627 22.721 20.667 ;
      RECT MASK 2 22.943 20.627 23.126 20.667 ;
      RECT MASK 2 25.67 20.627 25.853 20.667 ;
      RECT MASK 2 26.075 20.627 26.258 20.667 ;
      RECT MASK 2 26.832 20.627 27.015 20.667 ;
      RECT MASK 2 27.237 20.627 27.42 20.667 ;
      RECT MASK 2 27.994 20.627 28.177 20.667 ;
      RECT MASK 2 28.399 20.627 28.582 20.667 ;
      RECT MASK 2 29.156 20.627 29.339 20.667 ;
      RECT MASK 2 29.561 20.627 29.744 20.667 ;
      RECT MASK 2 32.288 20.627 32.471 20.667 ;
      RECT MASK 2 32.693 20.627 32.876 20.667 ;
      RECT MASK 2 33.45 20.627 33.633 20.667 ;
      RECT MASK 2 33.855 20.627 34.038 20.667 ;
      RECT MASK 2 34.612 20.627 34.795 20.667 ;
      RECT MASK 2 35.017 20.627 35.2 20.667 ;
      RECT MASK 2 35.774 20.627 35.957 20.667 ;
      RECT MASK 2 36.179 20.627 36.362 20.667 ;
      RECT MASK 2 38.906 20.627 39.089 20.667 ;
      RECT MASK 2 39.311 20.627 39.494 20.667 ;
      RECT MASK 2 40.068 20.627 40.251 20.667 ;
      RECT MASK 2 40.473 20.627 40.656 20.667 ;
      RECT MASK 2 41.23 20.627 41.413 20.667 ;
      RECT MASK 2 41.635 20.627 41.818 20.667 ;
      RECT MASK 2 42.392 20.627 42.575 20.667 ;
      RECT MASK 2 42.797 20.627 42.98 20.667 ;
      RECT MASK 2 45.524 20.627 45.707 20.667 ;
      RECT MASK 2 45.929 20.627 46.112 20.667 ;
      RECT MASK 2 46.686 20.627 46.869 20.667 ;
      RECT MASK 2 47.091 20.627 47.274 20.667 ;
      RECT MASK 2 47.848 20.627 48.031 20.667 ;
      RECT MASK 2 48.253 20.627 48.436 20.667 ;
      RECT MASK 2 49.01 20.627 49.193 20.667 ;
      RECT MASK 2 49.415 20.627 49.598 20.667 ;
      RECT MASK 2 52.142 20.627 52.325 20.667 ;
      RECT MASK 2 52.547 20.627 52.73 20.667 ;
      RECT MASK 2 53.304 20.627 53.487 20.667 ;
      RECT MASK 2 53.709 20.627 53.892 20.667 ;
      RECT MASK 2 54.466 20.627 54.649 20.667 ;
      RECT MASK 2 54.871 20.627 55.054 20.667 ;
      RECT MASK 2 55.628 20.627 55.811 20.667 ;
      RECT MASK 2 56.033 20.627 56.216 20.667 ;
      RECT MASK 2 58.76 20.627 58.943 20.667 ;
      RECT MASK 2 59.165 20.627 59.348 20.667 ;
      RECT MASK 2 59.922 20.627 60.105 20.667 ;
      RECT MASK 2 60.327 20.627 60.51 20.667 ;
      RECT MASK 2 61.084 20.627 61.267 20.667 ;
      RECT MASK 2 61.489 20.627 61.672 20.667 ;
      RECT MASK 2 62.246 20.627 62.429 20.667 ;
      RECT MASK 2 62.651 20.627 62.834 20.667 ;
      RECT MASK 2 65.378 20.627 65.561 20.667 ;
      RECT MASK 2 65.783 20.627 65.966 20.667 ;
      RECT MASK 2 66.54 20.627 66.723 20.667 ;
      RECT MASK 2 66.945 20.627 67.128 20.667 ;
      RECT MASK 2 67.702 20.627 67.885 20.667 ;
      RECT MASK 2 68.107 20.627 68.29 20.667 ;
      RECT MASK 2 68.864 20.627 69.047 20.667 ;
      RECT MASK 2 69.269 20.627 69.452 20.667 ;
      RECT MASK 2 71.996 20.627 72.179 20.667 ;
      RECT MASK 2 72.401 20.627 72.584 20.667 ;
      RECT MASK 2 73.158 20.627 73.341 20.667 ;
      RECT MASK 2 73.563 20.627 73.746 20.667 ;
      RECT MASK 2 74.32 20.627 74.503 20.667 ;
      RECT MASK 2 74.725 20.627 74.908 20.667 ;
      RECT MASK 2 75.482 20.627 75.665 20.667 ;
      RECT MASK 2 75.887 20.627 76.07 20.667 ;
      RECT MASK 2 78.614 20.627 78.797 20.667 ;
      RECT MASK 2 79.019 20.627 79.202 20.667 ;
      RECT MASK 2 79.776 20.627 79.959 20.667 ;
      RECT MASK 2 80.181 20.627 80.364 20.667 ;
      RECT MASK 2 80.938 20.627 81.121 20.667 ;
      RECT MASK 2 81.343 20.627 81.526 20.667 ;
      RECT MASK 2 82.1 20.627 82.283 20.667 ;
      RECT MASK 2 82.505 20.627 82.688 20.667 ;
      RECT MASK 2 85.232 20.627 85.415 20.667 ;
      RECT MASK 2 85.637 20.627 85.82 20.667 ;
      RECT MASK 2 86.394 20.627 86.577 20.667 ;
      RECT MASK 2 86.799 20.627 86.982 20.667 ;
      RECT MASK 2 87.556 20.627 87.739 20.667 ;
      RECT MASK 2 87.961 20.627 88.144 20.667 ;
      RECT MASK 2 88.718 20.627 88.901 20.667 ;
      RECT MASK 2 89.123 20.627 89.306 20.667 ;
      RECT MASK 2 91.85 20.627 92.033 20.667 ;
      RECT MASK 2 92.255 20.627 92.438 20.667 ;
      RECT MASK 2 93.012 20.627 93.195 20.667 ;
      RECT MASK 2 93.417 20.627 93.6 20.667 ;
      RECT MASK 2 94.174 20.627 94.357 20.667 ;
      RECT MASK 2 94.579 20.627 94.762 20.667 ;
      RECT MASK 2 95.336 20.627 95.519 20.667 ;
      RECT MASK 2 95.741 20.627 95.924 20.667 ;
      RECT MASK 2 98.468 20.627 98.651 20.667 ;
      RECT MASK 2 98.873 20.627 99.056 20.667 ;
      RECT MASK 2 99.63 20.627 99.813 20.667 ;
      RECT MASK 2 100.035 20.627 100.218 20.667 ;
      RECT MASK 2 100.792 20.627 100.975 20.667 ;
      RECT MASK 2 101.197 20.627 101.38 20.667 ;
      RECT MASK 2 101.954 20.627 102.137 20.667 ;
      RECT MASK 2 102.359 20.627 102.542 20.667 ;
      RECT MASK 2 105.086 20.627 105.269 20.667 ;
      RECT MASK 2 105.491 20.627 105.674 20.667 ;
      RECT MASK 2 106.248 20.627 106.431 20.667 ;
      RECT MASK 2 106.653 20.627 106.836 20.667 ;
      RECT MASK 2 107.41 20.627 107.593 20.667 ;
      RECT MASK 2 107.815 20.627 107.998 20.667 ;
      RECT MASK 2 108.572 20.627 108.755 20.667 ;
      RECT MASK 2 108.977 20.627 109.16 20.667 ;
      RECT MASK 2 116.291 20.7 116.351 21.75 ;
      RECT MASK 2 116.565 20.7 116.625 21.75 ;
      RECT MASK 2 116.839 20.7 116.899 21.75 ;
      RECT MASK 2 117.113 20.7 117.173 21.75 ;
      RECT MASK 2 117.387 20.7 117.447 21.75 ;
      RECT MASK 2 117.661 20.7 117.721 21.75 ;
      RECT MASK 2 117.935 20.7 117.995 21.75 ;
      RECT MASK 2 118.209 20.7 118.269 21.75 ;
      RECT MASK 2 118.483 20.7 118.543 21.75 ;
      RECT MASK 2 118.757 20.7 118.817 21.75 ;
      RECT MASK 2 119.031 20.7 119.091 21.75 ;
      RECT MASK 2 119.305 20.7 119.365 21.75 ;
      RECT MASK 2 119.579 20.7 119.639 21.75 ;
      RECT MASK 2 119.853 20.7 119.913 21.75 ;
      RECT MASK 2 120.127 20.7 120.187 21.75 ;
      RECT MASK 2 120.401 20.7 120.461 21.75 ;
      RECT MASK 2 120.675 20.7 120.735 21.75 ;
      RECT MASK 2 120.949 20.7 121.009 21.75 ;
      RECT MASK 2 121.223 20.7 121.283 21.75 ;
      RECT MASK 2 121.497 20.7 121.557 21.75 ;
      RECT MASK 2 121.771 20.7 121.831 21.75 ;
      RECT MASK 2 122.045 20.7 122.105 21.75 ;
      RECT MASK 2 122.319 20.7 122.379 21.75 ;
      RECT MASK 2 122.593 20.7 122.653 21.75 ;
      RECT MASK 2 122.867 20.7 122.927 21.75 ;
      RECT MASK 2 123.141 20.7 123.201 21.75 ;
      RECT MASK 2 123.415 20.7 123.475 21.75 ;
      RECT MASK 2 123.689 20.7 123.749 21.75 ;
      RECT MASK 2 123.963 20.7 124.023 21.75 ;
      RECT MASK 2 124.237 20.7 124.297 21.75 ;
      RECT MASK 2 124.511 20.7 124.571 21.75 ;
      RECT MASK 2 124.785 20.7 124.845 21.75 ;
      RECT MASK 2 125.059 20.7 125.119 21.75 ;
      RECT MASK 2 125.333 20.7 125.393 21.75 ;
      RECT MASK 2 125.607 20.7 125.667 21.75 ;
      RECT MASK 2 125.881 20.7 125.941 21.75 ;
      RECT MASK 2 126.155 20.7 126.215 21.75 ;
      RECT MASK 2 126.429 20.7 126.489 21.75 ;
      RECT MASK 2 126.703 20.7 126.763 21.75 ;
      RECT MASK 2 126.977 20.7 127.037 21.75 ;
      RECT MASK 2 127.251 20.7 127.311 21.75 ;
      RECT MASK 2 127.525 20.7 127.585 21.75 ;
      RECT MASK 2 127.799 20.7 127.859 21.75 ;
      RECT MASK 2 128.073 20.7 128.133 21.75 ;
      RECT MASK 2 5.107 20.811 109.869 20.851 ;
      RECT MASK 2 5.107 20.979 109.869 21.019 ;
      RECT MASK 2 5.1135 21.35 109.836 21.39 ;
      RECT MASK 2 2.362 21.48 2.422 22.53 ;
      RECT MASK 2 2.636 21.48 2.696 22.53 ;
      RECT MASK 2 2.91 21.48 2.97 22.53 ;
      RECT MASK 2 3.184 21.48 3.244 22.53 ;
      RECT MASK 2 3.458 21.48 3.518 22.53 ;
      RECT MASK 2 3.732 21.48 3.792 22.53 ;
      RECT MASK 2 5.1135 21.54 109.836 21.58 ;
      RECT MASK 2 5.655 22.098 5.735 22.3285 ;
      RECT MASK 2 5.987 22.098 6.067 22.3285 ;
      RECT MASK 2 6.319 22.098 6.399 22.3285 ;
      RECT MASK 2 6.817 22.098 6.897 22.3285 ;
      RECT MASK 2 7.149 22.098 7.229 22.3285 ;
      RECT MASK 2 7.481 22.098 7.561 22.3285 ;
      RECT MASK 2 7.979 22.098 8.059 22.3285 ;
      RECT MASK 2 8.311 22.098 8.391 22.3285 ;
      RECT MASK 2 8.643 22.098 8.723 22.3285 ;
      RECT MASK 2 9.141 22.098 9.221 22.3285 ;
      RECT MASK 2 9.473 22.098 9.553 22.3285 ;
      RECT MASK 2 9.805 22.098 9.885 22.3285 ;
      RECT MASK 2 12.273 22.098 12.353 22.3285 ;
      RECT MASK 2 12.605 22.098 12.685 22.3285 ;
      RECT MASK 2 12.937 22.098 13.017 22.3285 ;
      RECT MASK 2 13.435 22.098 13.515 22.3285 ;
      RECT MASK 2 13.767 22.098 13.847 22.3285 ;
      RECT MASK 2 14.099 22.098 14.179 22.3285 ;
      RECT MASK 2 14.597 22.098 14.677 22.3285 ;
      RECT MASK 2 14.929 22.098 15.009 22.3285 ;
      RECT MASK 2 15.261 22.098 15.341 22.3285 ;
      RECT MASK 2 15.759 22.098 15.839 22.3285 ;
      RECT MASK 2 16.091 22.098 16.171 22.3285 ;
      RECT MASK 2 16.423 22.098 16.503 22.3285 ;
      RECT MASK 2 18.891 22.098 18.971 22.3285 ;
      RECT MASK 2 19.223 22.098 19.303 22.3285 ;
      RECT MASK 2 19.555 22.098 19.635 22.3285 ;
      RECT MASK 2 20.053 22.098 20.133 22.3285 ;
      RECT MASK 2 20.385 22.098 20.465 22.3285 ;
      RECT MASK 2 20.717 22.098 20.797 22.3285 ;
      RECT MASK 2 21.215 22.098 21.295 22.3285 ;
      RECT MASK 2 21.547 22.098 21.627 22.3285 ;
      RECT MASK 2 21.879 22.098 21.959 22.3285 ;
      RECT MASK 2 22.377 22.098 22.457 22.3285 ;
      RECT MASK 2 22.709 22.098 22.789 22.3285 ;
      RECT MASK 2 23.041 22.098 23.121 22.3285 ;
      RECT MASK 2 25.509 22.098 25.589 22.3285 ;
      RECT MASK 2 25.841 22.098 25.921 22.3285 ;
      RECT MASK 2 26.173 22.098 26.253 22.3285 ;
      RECT MASK 2 26.671 22.098 26.751 22.3285 ;
      RECT MASK 2 27.003 22.098 27.083 22.3285 ;
      RECT MASK 2 27.335 22.098 27.415 22.3285 ;
      RECT MASK 2 27.833 22.098 27.913 22.3285 ;
      RECT MASK 2 28.165 22.098 28.245 22.3285 ;
      RECT MASK 2 28.497 22.098 28.577 22.3285 ;
      RECT MASK 2 28.995 22.098 29.075 22.3285 ;
      RECT MASK 2 29.327 22.098 29.407 22.3285 ;
      RECT MASK 2 29.659 22.098 29.739 22.3285 ;
      RECT MASK 2 32.127 22.098 32.207 22.3285 ;
      RECT MASK 2 32.459 22.098 32.539 22.3285 ;
      RECT MASK 2 32.791 22.098 32.871 22.3285 ;
      RECT MASK 2 33.289 22.098 33.369 22.3285 ;
      RECT MASK 2 33.621 22.098 33.701 22.3285 ;
      RECT MASK 2 33.953 22.098 34.033 22.3285 ;
      RECT MASK 2 34.451 22.098 34.531 22.3285 ;
      RECT MASK 2 34.783 22.098 34.863 22.3285 ;
      RECT MASK 2 35.115 22.098 35.195 22.3285 ;
      RECT MASK 2 35.613 22.098 35.693 22.3285 ;
      RECT MASK 2 35.945 22.098 36.025 22.3285 ;
      RECT MASK 2 36.277 22.098 36.357 22.3285 ;
      RECT MASK 2 38.745 22.098 38.825 22.3285 ;
      RECT MASK 2 39.077 22.098 39.157 22.3285 ;
      RECT MASK 2 39.409 22.098 39.489 22.3285 ;
      RECT MASK 2 39.907 22.098 39.987 22.3285 ;
      RECT MASK 2 40.239 22.098 40.319 22.3285 ;
      RECT MASK 2 40.571 22.098 40.651 22.3285 ;
      RECT MASK 2 41.069 22.098 41.149 22.3285 ;
      RECT MASK 2 41.401 22.098 41.481 22.3285 ;
      RECT MASK 2 41.733 22.098 41.813 22.3285 ;
      RECT MASK 2 42.231 22.098 42.311 22.3285 ;
      RECT MASK 2 42.563 22.098 42.643 22.3285 ;
      RECT MASK 2 42.895 22.098 42.975 22.3285 ;
      RECT MASK 2 45.363 22.098 45.443 22.3285 ;
      RECT MASK 2 45.695 22.098 45.775 22.3285 ;
      RECT MASK 2 46.027 22.098 46.107 22.3285 ;
      RECT MASK 2 46.525 22.098 46.605 22.3285 ;
      RECT MASK 2 46.857 22.098 46.937 22.3285 ;
      RECT MASK 2 47.189 22.098 47.269 22.3285 ;
      RECT MASK 2 47.687 22.098 47.767 22.3285 ;
      RECT MASK 2 48.019 22.098 48.099 22.3285 ;
      RECT MASK 2 48.351 22.098 48.431 22.3285 ;
      RECT MASK 2 48.849 22.098 48.929 22.3285 ;
      RECT MASK 2 49.181 22.098 49.261 22.3285 ;
      RECT MASK 2 49.513 22.098 49.593 22.3285 ;
      RECT MASK 2 51.981 22.098 52.061 22.3285 ;
      RECT MASK 2 52.313 22.098 52.393 22.3285 ;
      RECT MASK 2 52.645 22.098 52.725 22.3285 ;
      RECT MASK 2 53.143 22.098 53.223 22.3285 ;
      RECT MASK 2 53.475 22.098 53.555 22.3285 ;
      RECT MASK 2 53.807 22.098 53.887 22.3285 ;
      RECT MASK 2 54.305 22.098 54.385 22.3285 ;
      RECT MASK 2 54.637 22.098 54.717 22.3285 ;
      RECT MASK 2 54.969 22.098 55.049 22.3285 ;
      RECT MASK 2 55.467 22.098 55.547 22.3285 ;
      RECT MASK 2 55.799 22.098 55.879 22.3285 ;
      RECT MASK 2 56.131 22.098 56.211 22.3285 ;
      RECT MASK 2 58.599 22.098 58.679 22.3285 ;
      RECT MASK 2 58.931 22.098 59.011 22.3285 ;
      RECT MASK 2 59.263 22.098 59.343 22.3285 ;
      RECT MASK 2 59.761 22.098 59.841 22.3285 ;
      RECT MASK 2 60.093 22.098 60.173 22.3285 ;
      RECT MASK 2 60.425 22.098 60.505 22.3285 ;
      RECT MASK 2 60.923 22.098 61.003 22.3285 ;
      RECT MASK 2 61.255 22.098 61.335 22.3285 ;
      RECT MASK 2 61.587 22.098 61.667 22.3285 ;
      RECT MASK 2 62.085 22.098 62.165 22.3285 ;
      RECT MASK 2 62.417 22.098 62.497 22.3285 ;
      RECT MASK 2 62.749 22.098 62.829 22.3285 ;
      RECT MASK 2 65.217 22.098 65.297 22.3285 ;
      RECT MASK 2 65.549 22.098 65.629 22.3285 ;
      RECT MASK 2 65.881 22.098 65.961 22.3285 ;
      RECT MASK 2 66.379 22.098 66.459 22.3285 ;
      RECT MASK 2 66.711 22.098 66.791 22.3285 ;
      RECT MASK 2 67.043 22.098 67.123 22.3285 ;
      RECT MASK 2 67.541 22.098 67.621 22.3285 ;
      RECT MASK 2 67.873 22.098 67.953 22.3285 ;
      RECT MASK 2 68.205 22.098 68.285 22.3285 ;
      RECT MASK 2 68.703 22.098 68.783 22.3285 ;
      RECT MASK 2 69.035 22.098 69.115 22.3285 ;
      RECT MASK 2 69.367 22.098 69.447 22.3285 ;
      RECT MASK 2 71.835 22.098 71.915 22.3285 ;
      RECT MASK 2 72.167 22.098 72.247 22.3285 ;
      RECT MASK 2 72.499 22.098 72.579 22.3285 ;
      RECT MASK 2 72.997 22.098 73.077 22.3285 ;
      RECT MASK 2 73.329 22.098 73.409 22.3285 ;
      RECT MASK 2 73.661 22.098 73.741 22.3285 ;
      RECT MASK 2 74.159 22.098 74.239 22.3285 ;
      RECT MASK 2 74.491 22.098 74.571 22.3285 ;
      RECT MASK 2 74.823 22.098 74.903 22.3285 ;
      RECT MASK 2 75.321 22.098 75.401 22.3285 ;
      RECT MASK 2 75.653 22.098 75.733 22.3285 ;
      RECT MASK 2 75.985 22.098 76.065 22.3285 ;
      RECT MASK 2 78.453 22.098 78.533 22.3285 ;
      RECT MASK 2 78.785 22.098 78.865 22.3285 ;
      RECT MASK 2 79.117 22.098 79.197 22.3285 ;
      RECT MASK 2 79.615 22.098 79.695 22.3285 ;
      RECT MASK 2 79.947 22.098 80.027 22.3285 ;
      RECT MASK 2 80.279 22.098 80.359 22.3285 ;
      RECT MASK 2 80.777 22.098 80.857 22.3285 ;
      RECT MASK 2 81.109 22.098 81.189 22.3285 ;
      RECT MASK 2 81.441 22.098 81.521 22.3285 ;
      RECT MASK 2 81.939 22.098 82.019 22.3285 ;
      RECT MASK 2 82.271 22.098 82.351 22.3285 ;
      RECT MASK 2 82.603 22.098 82.683 22.3285 ;
      RECT MASK 2 85.071 22.098 85.151 22.3285 ;
      RECT MASK 2 85.403 22.098 85.483 22.3285 ;
      RECT MASK 2 85.735 22.098 85.815 22.3285 ;
      RECT MASK 2 86.233 22.098 86.313 22.3285 ;
      RECT MASK 2 86.565 22.098 86.645 22.3285 ;
      RECT MASK 2 86.897 22.098 86.977 22.3285 ;
      RECT MASK 2 87.395 22.098 87.475 22.3285 ;
      RECT MASK 2 87.727 22.098 87.807 22.3285 ;
      RECT MASK 2 88.059 22.098 88.139 22.3285 ;
      RECT MASK 2 88.557 22.098 88.637 22.3285 ;
      RECT MASK 2 88.889 22.098 88.969 22.3285 ;
      RECT MASK 2 89.221 22.098 89.301 22.3285 ;
      RECT MASK 2 91.689 22.098 91.769 22.3285 ;
      RECT MASK 2 92.021 22.098 92.101 22.3285 ;
      RECT MASK 2 92.353 22.098 92.433 22.3285 ;
      RECT MASK 2 92.851 22.098 92.931 22.3285 ;
      RECT MASK 2 93.183 22.098 93.263 22.3285 ;
      RECT MASK 2 93.515 22.098 93.595 22.3285 ;
      RECT MASK 2 94.013 22.098 94.093 22.3285 ;
      RECT MASK 2 94.345 22.098 94.425 22.3285 ;
      RECT MASK 2 94.677 22.098 94.757 22.3285 ;
      RECT MASK 2 95.175 22.098 95.255 22.3285 ;
      RECT MASK 2 95.507 22.098 95.587 22.3285 ;
      RECT MASK 2 95.839 22.098 95.919 22.3285 ;
      RECT MASK 2 98.307 22.098 98.387 22.3285 ;
      RECT MASK 2 98.639 22.098 98.719 22.3285 ;
      RECT MASK 2 98.971 22.098 99.051 22.3285 ;
      RECT MASK 2 99.469 22.098 99.549 22.3285 ;
      RECT MASK 2 99.801 22.098 99.881 22.3285 ;
      RECT MASK 2 100.133 22.098 100.213 22.3285 ;
      RECT MASK 2 100.631 22.098 100.711 22.3285 ;
      RECT MASK 2 100.963 22.098 101.043 22.3285 ;
      RECT MASK 2 101.295 22.098 101.375 22.3285 ;
      RECT MASK 2 101.793 22.098 101.873 22.3285 ;
      RECT MASK 2 102.125 22.098 102.205 22.3285 ;
      RECT MASK 2 102.457 22.098 102.537 22.3285 ;
      RECT MASK 2 104.925 22.098 105.005 22.3285 ;
      RECT MASK 2 105.257 22.098 105.337 22.3285 ;
      RECT MASK 2 105.589 22.098 105.669 22.3285 ;
      RECT MASK 2 106.087 22.098 106.167 22.3285 ;
      RECT MASK 2 106.419 22.098 106.499 22.3285 ;
      RECT MASK 2 106.751 22.098 106.831 22.3285 ;
      RECT MASK 2 107.249 22.098 107.329 22.3285 ;
      RECT MASK 2 107.581 22.098 107.661 22.3285 ;
      RECT MASK 2 107.913 22.098 107.993 22.3285 ;
      RECT MASK 2 108.411 22.098 108.491 22.3285 ;
      RECT MASK 2 108.743 22.098 108.823 22.3285 ;
      RECT MASK 2 109.075 22.098 109.155 22.3285 ;
      RECT MASK 2 116.291 22.41 116.351 23.46 ;
      RECT MASK 2 116.565 22.41 116.625 23.46 ;
      RECT MASK 2 116.839 22.41 116.899 23.46 ;
      RECT MASK 2 117.113 22.41 117.173 23.46 ;
      RECT MASK 2 117.387 22.41 117.447 23.46 ;
      RECT MASK 2 117.661 22.41 117.721 23.46 ;
      RECT MASK 2 117.935 22.41 117.995 23.46 ;
      RECT MASK 2 118.209 22.41 118.269 23.46 ;
      RECT MASK 2 118.483 22.41 118.543 23.46 ;
      RECT MASK 2 118.757 22.41 118.817 23.46 ;
      RECT MASK 2 119.031 22.41 119.091 23.46 ;
      RECT MASK 2 119.305 22.41 119.365 23.46 ;
      RECT MASK 2 119.579 22.41 119.639 23.46 ;
      RECT MASK 2 119.853 22.41 119.913 23.46 ;
      RECT MASK 2 120.127 22.41 120.187 23.46 ;
      RECT MASK 2 120.401 22.41 120.461 23.46 ;
      RECT MASK 2 120.675 22.41 120.735 23.46 ;
      RECT MASK 2 120.949 22.41 121.009 23.46 ;
      RECT MASK 2 121.223 22.41 121.283 23.46 ;
      RECT MASK 2 121.497 22.41 121.557 23.46 ;
      RECT MASK 2 121.771 22.41 121.831 23.46 ;
      RECT MASK 2 122.045 22.41 122.105 23.46 ;
      RECT MASK 2 122.319 22.41 122.379 23.46 ;
      RECT MASK 2 122.593 22.41 122.653 23.46 ;
      RECT MASK 2 122.867 22.41 122.927 23.46 ;
      RECT MASK 2 123.141 22.41 123.201 23.46 ;
      RECT MASK 2 123.415 22.41 123.475 23.46 ;
      RECT MASK 2 123.689 22.41 123.749 23.46 ;
      RECT MASK 2 123.963 22.41 124.023 23.46 ;
      RECT MASK 2 124.237 22.41 124.297 23.46 ;
      RECT MASK 2 124.511 22.41 124.571 23.46 ;
      RECT MASK 2 124.785 22.41 124.845 23.46 ;
      RECT MASK 2 125.059 22.41 125.119 23.46 ;
      RECT MASK 2 125.333 22.41 125.393 23.46 ;
      RECT MASK 2 125.607 22.41 125.667 23.46 ;
      RECT MASK 2 125.881 22.41 125.941 23.46 ;
      RECT MASK 2 126.155 22.41 126.215 23.46 ;
      RECT MASK 2 126.429 22.41 126.489 23.46 ;
      RECT MASK 2 126.703 22.41 126.763 23.46 ;
      RECT MASK 2 126.977 22.41 127.037 23.46 ;
      RECT MASK 2 127.251 22.41 127.311 23.46 ;
      RECT MASK 2 127.525 22.41 127.585 23.46 ;
      RECT MASK 2 127.799 22.41 127.859 23.46 ;
      RECT MASK 2 128.073 22.41 128.133 23.46 ;
      RECT MASK 2 5.655 22.769 5.735 22.994 ;
      RECT MASK 2 5.987 22.769 6.067 22.994 ;
      RECT MASK 2 6.319 22.769 6.399 22.994 ;
      RECT MASK 2 6.817 22.769 6.897 22.994 ;
      RECT MASK 2 7.149 22.769 7.229 22.994 ;
      RECT MASK 2 7.481 22.769 7.561 22.994 ;
      RECT MASK 2 7.979 22.769 8.059 22.994 ;
      RECT MASK 2 8.311 22.769 8.391 22.994 ;
      RECT MASK 2 8.643 22.769 8.723 22.994 ;
      RECT MASK 2 9.141 22.769 9.221 22.994 ;
      RECT MASK 2 9.473 22.769 9.553 22.994 ;
      RECT MASK 2 9.805 22.769 9.885 22.994 ;
      RECT MASK 2 12.273 22.769 12.353 22.994 ;
      RECT MASK 2 12.605 22.769 12.685 22.994 ;
      RECT MASK 2 12.937 22.769 13.017 22.994 ;
      RECT MASK 2 13.435 22.769 13.515 22.994 ;
      RECT MASK 2 13.767 22.769 13.847 22.994 ;
      RECT MASK 2 14.099 22.769 14.179 22.994 ;
      RECT MASK 2 14.597 22.769 14.677 22.994 ;
      RECT MASK 2 14.929 22.769 15.009 22.994 ;
      RECT MASK 2 15.261 22.769 15.341 22.994 ;
      RECT MASK 2 15.759 22.769 15.839 22.994 ;
      RECT MASK 2 16.091 22.769 16.171 22.994 ;
      RECT MASK 2 16.423 22.769 16.503 22.994 ;
      RECT MASK 2 18.891 22.769 18.971 22.994 ;
      RECT MASK 2 19.223 22.769 19.303 22.994 ;
      RECT MASK 2 19.555 22.769 19.635 22.994 ;
      RECT MASK 2 20.053 22.769 20.133 22.994 ;
      RECT MASK 2 20.385 22.769 20.465 22.994 ;
      RECT MASK 2 20.717 22.769 20.797 22.994 ;
      RECT MASK 2 21.215 22.769 21.295 22.994 ;
      RECT MASK 2 21.547 22.769 21.627 22.994 ;
      RECT MASK 2 21.879 22.769 21.959 22.994 ;
      RECT MASK 2 22.377 22.769 22.457 22.994 ;
      RECT MASK 2 22.709 22.769 22.789 22.994 ;
      RECT MASK 2 23.041 22.769 23.121 22.994 ;
      RECT MASK 2 25.509 22.769 25.589 22.994 ;
      RECT MASK 2 25.841 22.769 25.921 22.994 ;
      RECT MASK 2 26.173 22.769 26.253 22.994 ;
      RECT MASK 2 26.671 22.769 26.751 22.994 ;
      RECT MASK 2 27.003 22.769 27.083 22.994 ;
      RECT MASK 2 27.335 22.769 27.415 22.994 ;
      RECT MASK 2 27.833 22.769 27.913 22.994 ;
      RECT MASK 2 28.165 22.769 28.245 22.994 ;
      RECT MASK 2 28.497 22.769 28.577 22.994 ;
      RECT MASK 2 28.995 22.769 29.075 22.994 ;
      RECT MASK 2 29.327 22.769 29.407 22.994 ;
      RECT MASK 2 29.659 22.769 29.739 22.994 ;
      RECT MASK 2 32.127 22.769 32.207 22.994 ;
      RECT MASK 2 32.459 22.769 32.539 22.994 ;
      RECT MASK 2 32.791 22.769 32.871 22.994 ;
      RECT MASK 2 33.289 22.769 33.369 22.994 ;
      RECT MASK 2 33.621 22.769 33.701 22.994 ;
      RECT MASK 2 33.953 22.769 34.033 22.994 ;
      RECT MASK 2 34.451 22.769 34.531 22.994 ;
      RECT MASK 2 34.783 22.769 34.863 22.994 ;
      RECT MASK 2 35.115 22.769 35.195 22.994 ;
      RECT MASK 2 35.613 22.769 35.693 22.994 ;
      RECT MASK 2 35.945 22.769 36.025 22.994 ;
      RECT MASK 2 36.277 22.769 36.357 22.994 ;
      RECT MASK 2 38.745 22.769 38.825 22.994 ;
      RECT MASK 2 39.077 22.769 39.157 22.994 ;
      RECT MASK 2 39.409 22.769 39.489 22.994 ;
      RECT MASK 2 39.907 22.769 39.987 22.994 ;
      RECT MASK 2 40.239 22.769 40.319 22.994 ;
      RECT MASK 2 40.571 22.769 40.651 22.994 ;
      RECT MASK 2 41.069 22.769 41.149 22.994 ;
      RECT MASK 2 41.401 22.769 41.481 22.994 ;
      RECT MASK 2 41.733 22.769 41.813 22.994 ;
      RECT MASK 2 42.231 22.769 42.311 22.994 ;
      RECT MASK 2 42.563 22.769 42.643 22.994 ;
      RECT MASK 2 42.895 22.769 42.975 22.994 ;
      RECT MASK 2 45.363 22.769 45.443 22.994 ;
      RECT MASK 2 45.695 22.769 45.775 22.994 ;
      RECT MASK 2 46.027 22.769 46.107 22.994 ;
      RECT MASK 2 46.525 22.769 46.605 22.994 ;
      RECT MASK 2 46.857 22.769 46.937 22.994 ;
      RECT MASK 2 47.189 22.769 47.269 22.994 ;
      RECT MASK 2 47.687 22.769 47.767 22.994 ;
      RECT MASK 2 48.019 22.769 48.099 22.994 ;
      RECT MASK 2 48.351 22.769 48.431 22.994 ;
      RECT MASK 2 48.849 22.769 48.929 22.994 ;
      RECT MASK 2 49.181 22.769 49.261 22.994 ;
      RECT MASK 2 49.513 22.769 49.593 22.994 ;
      RECT MASK 2 51.981 22.769 52.061 22.994 ;
      RECT MASK 2 52.313 22.769 52.393 22.994 ;
      RECT MASK 2 52.645 22.769 52.725 22.994 ;
      RECT MASK 2 53.143 22.769 53.223 22.994 ;
      RECT MASK 2 53.475 22.769 53.555 22.994 ;
      RECT MASK 2 53.807 22.769 53.887 22.994 ;
      RECT MASK 2 54.305 22.769 54.385 22.994 ;
      RECT MASK 2 54.637 22.769 54.717 22.994 ;
      RECT MASK 2 54.969 22.769 55.049 22.994 ;
      RECT MASK 2 55.467 22.769 55.547 22.994 ;
      RECT MASK 2 55.799 22.769 55.879 22.994 ;
      RECT MASK 2 56.131 22.769 56.211 22.994 ;
      RECT MASK 2 58.599 22.769 58.679 22.994 ;
      RECT MASK 2 58.931 22.769 59.011 22.994 ;
      RECT MASK 2 59.263 22.769 59.343 22.994 ;
      RECT MASK 2 59.761 22.769 59.841 22.994 ;
      RECT MASK 2 60.093 22.769 60.173 22.994 ;
      RECT MASK 2 60.425 22.769 60.505 22.994 ;
      RECT MASK 2 60.923 22.769 61.003 22.994 ;
      RECT MASK 2 61.255 22.769 61.335 22.994 ;
      RECT MASK 2 61.587 22.769 61.667 22.994 ;
      RECT MASK 2 62.085 22.769 62.165 22.994 ;
      RECT MASK 2 62.417 22.769 62.497 22.994 ;
      RECT MASK 2 62.749 22.769 62.829 22.994 ;
      RECT MASK 2 65.217 22.769 65.297 22.994 ;
      RECT MASK 2 65.549 22.769 65.629 22.994 ;
      RECT MASK 2 65.881 22.769 65.961 22.994 ;
      RECT MASK 2 66.379 22.769 66.459 22.994 ;
      RECT MASK 2 66.711 22.769 66.791 22.994 ;
      RECT MASK 2 67.043 22.769 67.123 22.994 ;
      RECT MASK 2 67.541 22.769 67.621 22.994 ;
      RECT MASK 2 67.873 22.769 67.953 22.994 ;
      RECT MASK 2 68.205 22.769 68.285 22.994 ;
      RECT MASK 2 68.703 22.769 68.783 22.994 ;
      RECT MASK 2 69.035 22.769 69.115 22.994 ;
      RECT MASK 2 69.367 22.769 69.447 22.994 ;
      RECT MASK 2 71.835 22.769 71.915 22.994 ;
      RECT MASK 2 72.167 22.769 72.247 22.994 ;
      RECT MASK 2 72.499 22.769 72.579 22.994 ;
      RECT MASK 2 72.997 22.769 73.077 22.994 ;
      RECT MASK 2 73.329 22.769 73.409 22.994 ;
      RECT MASK 2 73.661 22.769 73.741 22.994 ;
      RECT MASK 2 74.159 22.769 74.239 22.994 ;
      RECT MASK 2 74.491 22.769 74.571 22.994 ;
      RECT MASK 2 74.823 22.769 74.903 22.994 ;
      RECT MASK 2 75.321 22.769 75.401 22.994 ;
      RECT MASK 2 75.653 22.769 75.733 22.994 ;
      RECT MASK 2 75.985 22.769 76.065 22.994 ;
      RECT MASK 2 78.453 22.769 78.533 22.994 ;
      RECT MASK 2 78.785 22.769 78.865 22.994 ;
      RECT MASK 2 79.117 22.769 79.197 22.994 ;
      RECT MASK 2 79.615 22.769 79.695 22.994 ;
      RECT MASK 2 79.947 22.769 80.027 22.994 ;
      RECT MASK 2 80.279 22.769 80.359 22.994 ;
      RECT MASK 2 80.777 22.769 80.857 22.994 ;
      RECT MASK 2 81.109 22.769 81.189 22.994 ;
      RECT MASK 2 81.441 22.769 81.521 22.994 ;
      RECT MASK 2 81.939 22.769 82.019 22.994 ;
      RECT MASK 2 82.271 22.769 82.351 22.994 ;
      RECT MASK 2 82.603 22.769 82.683 22.994 ;
      RECT MASK 2 85.071 22.769 85.151 22.994 ;
      RECT MASK 2 85.403 22.769 85.483 22.994 ;
      RECT MASK 2 85.735 22.769 85.815 22.994 ;
      RECT MASK 2 86.233 22.769 86.313 22.994 ;
      RECT MASK 2 86.565 22.769 86.645 22.994 ;
      RECT MASK 2 86.897 22.769 86.977 22.994 ;
      RECT MASK 2 87.395 22.769 87.475 22.994 ;
      RECT MASK 2 87.727 22.769 87.807 22.994 ;
      RECT MASK 2 88.059 22.769 88.139 22.994 ;
      RECT MASK 2 88.557 22.769 88.637 22.994 ;
      RECT MASK 2 88.889 22.769 88.969 22.994 ;
      RECT MASK 2 89.221 22.769 89.301 22.994 ;
      RECT MASK 2 91.689 22.769 91.769 22.994 ;
      RECT MASK 2 92.021 22.769 92.101 22.994 ;
      RECT MASK 2 92.353 22.769 92.433 22.994 ;
      RECT MASK 2 92.851 22.769 92.931 22.994 ;
      RECT MASK 2 93.183 22.769 93.263 22.994 ;
      RECT MASK 2 93.515 22.769 93.595 22.994 ;
      RECT MASK 2 94.013 22.769 94.093 22.994 ;
      RECT MASK 2 94.345 22.769 94.425 22.994 ;
      RECT MASK 2 94.677 22.769 94.757 22.994 ;
      RECT MASK 2 95.175 22.769 95.255 22.994 ;
      RECT MASK 2 95.507 22.769 95.587 22.994 ;
      RECT MASK 2 95.839 22.769 95.919 22.994 ;
      RECT MASK 2 98.307 22.769 98.387 22.994 ;
      RECT MASK 2 98.639 22.769 98.719 22.994 ;
      RECT MASK 2 98.971 22.769 99.051 22.994 ;
      RECT MASK 2 99.469 22.769 99.549 22.994 ;
      RECT MASK 2 99.801 22.769 99.881 22.994 ;
      RECT MASK 2 100.133 22.769 100.213 22.994 ;
      RECT MASK 2 100.631 22.769 100.711 22.994 ;
      RECT MASK 2 100.963 22.769 101.043 22.994 ;
      RECT MASK 2 101.295 22.769 101.375 22.994 ;
      RECT MASK 2 101.793 22.769 101.873 22.994 ;
      RECT MASK 2 102.125 22.769 102.205 22.994 ;
      RECT MASK 2 102.457 22.769 102.537 22.994 ;
      RECT MASK 2 104.925 22.769 105.005 22.994 ;
      RECT MASK 2 105.257 22.769 105.337 22.994 ;
      RECT MASK 2 105.589 22.769 105.669 22.994 ;
      RECT MASK 2 106.087 22.769 106.167 22.994 ;
      RECT MASK 2 106.419 22.769 106.499 22.994 ;
      RECT MASK 2 106.751 22.769 106.831 22.994 ;
      RECT MASK 2 107.249 22.769 107.329 22.994 ;
      RECT MASK 2 107.581 22.769 107.661 22.994 ;
      RECT MASK 2 107.913 22.769 107.993 22.994 ;
      RECT MASK 2 108.411 22.769 108.491 22.994 ;
      RECT MASK 2 108.743 22.769 108.823 22.994 ;
      RECT MASK 2 109.075 22.769 109.155 22.994 ;
      RECT MASK 2 2.362 23.19 2.422 24.24 ;
      RECT MASK 2 2.636 23.19 2.696 24.24 ;
      RECT MASK 2 2.91 23.19 2.97 24.24 ;
      RECT MASK 2 3.184 23.19 3.244 24.24 ;
      RECT MASK 2 3.458 23.19 3.518 24.24 ;
      RECT MASK 2 3.732 23.19 3.792 24.24 ;
      RECT MASK 2 5.1135 23.3 109.836 23.34 ;
      RECT MASK 2 5.1135 23.49 109.836 23.53 ;
      RECT MASK 2 5.1135 23.75 110.065 23.79 ;
      RECT MASK 2 115.425 23.75 129.001 23.79 ;
      RECT MASK 2 5.1135 23.94 110.065 23.98 ;
      RECT MASK 2 115.425 23.94 129.001 23.98 ;
      RECT MASK 2 5.655 24.502 5.735 24.7285 ;
      RECT MASK 2 5.987 24.502 6.067 24.7285 ;
      RECT MASK 2 6.319 24.502 6.399 24.7285 ;
      RECT MASK 2 6.817 24.502 6.897 24.7285 ;
      RECT MASK 2 7.149 24.502 7.229 24.7285 ;
      RECT MASK 2 7.481 24.502 7.561 24.7285 ;
      RECT MASK 2 7.979 24.502 8.059 24.7285 ;
      RECT MASK 2 8.311 24.502 8.391 24.7285 ;
      RECT MASK 2 8.643 24.502 8.723 24.7285 ;
      RECT MASK 2 9.141 24.502 9.221 24.7285 ;
      RECT MASK 2 9.473 24.502 9.553 24.7285 ;
      RECT MASK 2 9.805 24.502 9.885 24.7285 ;
      RECT MASK 2 12.273 24.502 12.353 24.7285 ;
      RECT MASK 2 12.605 24.502 12.685 24.7285 ;
      RECT MASK 2 12.937 24.502 13.017 24.7285 ;
      RECT MASK 2 13.435 24.502 13.515 24.7285 ;
      RECT MASK 2 13.767 24.502 13.847 24.7285 ;
      RECT MASK 2 14.099 24.502 14.179 24.7285 ;
      RECT MASK 2 14.597 24.502 14.677 24.7285 ;
      RECT MASK 2 14.929 24.502 15.009 24.7285 ;
      RECT MASK 2 15.261 24.502 15.341 24.7285 ;
      RECT MASK 2 15.759 24.502 15.839 24.7285 ;
      RECT MASK 2 16.091 24.502 16.171 24.7285 ;
      RECT MASK 2 16.423 24.502 16.503 24.7285 ;
      RECT MASK 2 18.891 24.502 18.971 24.7285 ;
      RECT MASK 2 19.223 24.502 19.303 24.7285 ;
      RECT MASK 2 19.555 24.502 19.635 24.7285 ;
      RECT MASK 2 20.053 24.502 20.133 24.7285 ;
      RECT MASK 2 20.385 24.502 20.465 24.7285 ;
      RECT MASK 2 20.717 24.502 20.797 24.7285 ;
      RECT MASK 2 21.215 24.502 21.295 24.7285 ;
      RECT MASK 2 21.547 24.502 21.627 24.7285 ;
      RECT MASK 2 21.879 24.502 21.959 24.7285 ;
      RECT MASK 2 22.377 24.502 22.457 24.7285 ;
      RECT MASK 2 22.709 24.502 22.789 24.7285 ;
      RECT MASK 2 23.041 24.502 23.121 24.7285 ;
      RECT MASK 2 25.509 24.502 25.589 24.7285 ;
      RECT MASK 2 25.841 24.502 25.921 24.7285 ;
      RECT MASK 2 26.173 24.502 26.253 24.7285 ;
      RECT MASK 2 26.671 24.502 26.751 24.7285 ;
      RECT MASK 2 27.003 24.502 27.083 24.7285 ;
      RECT MASK 2 27.335 24.502 27.415 24.7285 ;
      RECT MASK 2 27.833 24.502 27.913 24.7285 ;
      RECT MASK 2 28.165 24.502 28.245 24.7285 ;
      RECT MASK 2 28.497 24.502 28.577 24.7285 ;
      RECT MASK 2 28.995 24.502 29.075 24.7285 ;
      RECT MASK 2 29.327 24.502 29.407 24.7285 ;
      RECT MASK 2 29.659 24.502 29.739 24.7285 ;
      RECT MASK 2 32.127 24.502 32.207 24.7285 ;
      RECT MASK 2 32.459 24.502 32.539 24.7285 ;
      RECT MASK 2 32.791 24.502 32.871 24.7285 ;
      RECT MASK 2 33.289 24.502 33.369 24.7285 ;
      RECT MASK 2 33.621 24.502 33.701 24.7285 ;
      RECT MASK 2 33.953 24.502 34.033 24.7285 ;
      RECT MASK 2 34.451 24.502 34.531 24.7285 ;
      RECT MASK 2 34.783 24.502 34.863 24.7285 ;
      RECT MASK 2 35.115 24.502 35.195 24.7285 ;
      RECT MASK 2 35.613 24.502 35.693 24.7285 ;
      RECT MASK 2 35.945 24.502 36.025 24.7285 ;
      RECT MASK 2 36.277 24.502 36.357 24.7285 ;
      RECT MASK 2 38.745 24.502 38.825 24.7285 ;
      RECT MASK 2 39.077 24.502 39.157 24.7285 ;
      RECT MASK 2 39.409 24.502 39.489 24.7285 ;
      RECT MASK 2 39.907 24.502 39.987 24.7285 ;
      RECT MASK 2 40.239 24.502 40.319 24.7285 ;
      RECT MASK 2 40.571 24.502 40.651 24.7285 ;
      RECT MASK 2 41.069 24.502 41.149 24.7285 ;
      RECT MASK 2 41.401 24.502 41.481 24.7285 ;
      RECT MASK 2 41.733 24.502 41.813 24.7285 ;
      RECT MASK 2 42.231 24.502 42.311 24.7285 ;
      RECT MASK 2 42.563 24.502 42.643 24.7285 ;
      RECT MASK 2 42.895 24.502 42.975 24.7285 ;
      RECT MASK 2 45.363 24.502 45.443 24.7285 ;
      RECT MASK 2 45.695 24.502 45.775 24.7285 ;
      RECT MASK 2 46.027 24.502 46.107 24.7285 ;
      RECT MASK 2 46.525 24.502 46.605 24.7285 ;
      RECT MASK 2 46.857 24.502 46.937 24.7285 ;
      RECT MASK 2 47.189 24.502 47.269 24.7285 ;
      RECT MASK 2 47.687 24.502 47.767 24.7285 ;
      RECT MASK 2 48.019 24.502 48.099 24.7285 ;
      RECT MASK 2 48.351 24.502 48.431 24.7285 ;
      RECT MASK 2 48.849 24.502 48.929 24.7285 ;
      RECT MASK 2 49.181 24.502 49.261 24.7285 ;
      RECT MASK 2 49.513 24.502 49.593 24.7285 ;
      RECT MASK 2 51.981 24.502 52.061 24.7285 ;
      RECT MASK 2 52.313 24.502 52.393 24.7285 ;
      RECT MASK 2 52.645 24.502 52.725 24.7285 ;
      RECT MASK 2 53.143 24.502 53.223 24.7285 ;
      RECT MASK 2 53.475 24.502 53.555 24.7285 ;
      RECT MASK 2 53.807 24.502 53.887 24.7285 ;
      RECT MASK 2 54.305 24.502 54.385 24.7285 ;
      RECT MASK 2 54.637 24.502 54.717 24.7285 ;
      RECT MASK 2 54.969 24.502 55.049 24.7285 ;
      RECT MASK 2 55.467 24.502 55.547 24.7285 ;
      RECT MASK 2 55.799 24.502 55.879 24.7285 ;
      RECT MASK 2 56.131 24.502 56.211 24.7285 ;
      RECT MASK 2 58.599 24.502 58.679 24.7285 ;
      RECT MASK 2 58.931 24.502 59.011 24.7285 ;
      RECT MASK 2 59.263 24.502 59.343 24.7285 ;
      RECT MASK 2 59.761 24.502 59.841 24.7285 ;
      RECT MASK 2 60.093 24.502 60.173 24.7285 ;
      RECT MASK 2 60.425 24.502 60.505 24.7285 ;
      RECT MASK 2 60.923 24.502 61.003 24.7285 ;
      RECT MASK 2 61.255 24.502 61.335 24.7285 ;
      RECT MASK 2 61.587 24.502 61.667 24.7285 ;
      RECT MASK 2 62.085 24.502 62.165 24.7285 ;
      RECT MASK 2 62.417 24.502 62.497 24.7285 ;
      RECT MASK 2 62.749 24.502 62.829 24.7285 ;
      RECT MASK 2 65.217 24.502 65.297 24.7285 ;
      RECT MASK 2 65.549 24.502 65.629 24.7285 ;
      RECT MASK 2 65.881 24.502 65.961 24.7285 ;
      RECT MASK 2 66.379 24.502 66.459 24.7285 ;
      RECT MASK 2 66.711 24.502 66.791 24.7285 ;
      RECT MASK 2 67.043 24.502 67.123 24.7285 ;
      RECT MASK 2 67.541 24.502 67.621 24.7285 ;
      RECT MASK 2 67.873 24.502 67.953 24.7285 ;
      RECT MASK 2 68.205 24.502 68.285 24.7285 ;
      RECT MASK 2 68.703 24.502 68.783 24.7285 ;
      RECT MASK 2 69.035 24.502 69.115 24.7285 ;
      RECT MASK 2 69.367 24.502 69.447 24.7285 ;
      RECT MASK 2 71.835 24.502 71.915 24.7285 ;
      RECT MASK 2 72.167 24.502 72.247 24.7285 ;
      RECT MASK 2 72.499 24.502 72.579 24.7285 ;
      RECT MASK 2 72.997 24.502 73.077 24.7285 ;
      RECT MASK 2 73.329 24.502 73.409 24.7285 ;
      RECT MASK 2 73.661 24.502 73.741 24.7285 ;
      RECT MASK 2 74.159 24.502 74.239 24.7285 ;
      RECT MASK 2 74.491 24.502 74.571 24.7285 ;
      RECT MASK 2 74.823 24.502 74.903 24.7285 ;
      RECT MASK 2 75.321 24.502 75.401 24.7285 ;
      RECT MASK 2 75.653 24.502 75.733 24.7285 ;
      RECT MASK 2 75.985 24.502 76.065 24.7285 ;
      RECT MASK 2 78.453 24.502 78.533 24.7285 ;
      RECT MASK 2 78.785 24.502 78.865 24.7285 ;
      RECT MASK 2 79.117 24.502 79.197 24.7285 ;
      RECT MASK 2 79.615 24.502 79.695 24.7285 ;
      RECT MASK 2 79.947 24.502 80.027 24.7285 ;
      RECT MASK 2 80.279 24.502 80.359 24.7285 ;
      RECT MASK 2 80.777 24.502 80.857 24.7285 ;
      RECT MASK 2 81.109 24.502 81.189 24.7285 ;
      RECT MASK 2 81.441 24.502 81.521 24.7285 ;
      RECT MASK 2 81.939 24.502 82.019 24.7285 ;
      RECT MASK 2 82.271 24.502 82.351 24.7285 ;
      RECT MASK 2 82.603 24.502 82.683 24.7285 ;
      RECT MASK 2 85.071 24.502 85.151 24.7285 ;
      RECT MASK 2 85.403 24.502 85.483 24.7285 ;
      RECT MASK 2 85.735 24.502 85.815 24.7285 ;
      RECT MASK 2 86.233 24.502 86.313 24.7285 ;
      RECT MASK 2 86.565 24.502 86.645 24.7285 ;
      RECT MASK 2 86.897 24.502 86.977 24.7285 ;
      RECT MASK 2 87.395 24.502 87.475 24.7285 ;
      RECT MASK 2 87.727 24.502 87.807 24.7285 ;
      RECT MASK 2 88.059 24.502 88.139 24.7285 ;
      RECT MASK 2 88.557 24.502 88.637 24.7285 ;
      RECT MASK 2 88.889 24.502 88.969 24.7285 ;
      RECT MASK 2 89.221 24.502 89.301 24.7285 ;
      RECT MASK 2 91.689 24.502 91.769 24.7285 ;
      RECT MASK 2 92.021 24.502 92.101 24.7285 ;
      RECT MASK 2 92.353 24.502 92.433 24.7285 ;
      RECT MASK 2 92.851 24.502 92.931 24.7285 ;
      RECT MASK 2 93.183 24.502 93.263 24.7285 ;
      RECT MASK 2 93.515 24.502 93.595 24.7285 ;
      RECT MASK 2 94.013 24.502 94.093 24.7285 ;
      RECT MASK 2 94.345 24.502 94.425 24.7285 ;
      RECT MASK 2 94.677 24.502 94.757 24.7285 ;
      RECT MASK 2 95.175 24.502 95.255 24.7285 ;
      RECT MASK 2 95.507 24.502 95.587 24.7285 ;
      RECT MASK 2 95.839 24.502 95.919 24.7285 ;
      RECT MASK 2 98.307 24.502 98.387 24.7285 ;
      RECT MASK 2 98.639 24.502 98.719 24.7285 ;
      RECT MASK 2 98.971 24.502 99.051 24.7285 ;
      RECT MASK 2 99.469 24.502 99.549 24.7285 ;
      RECT MASK 2 99.801 24.502 99.881 24.7285 ;
      RECT MASK 2 100.133 24.502 100.213 24.7285 ;
      RECT MASK 2 100.631 24.502 100.711 24.7285 ;
      RECT MASK 2 100.963 24.502 101.043 24.7285 ;
      RECT MASK 2 101.295 24.502 101.375 24.7285 ;
      RECT MASK 2 101.793 24.502 101.873 24.7285 ;
      RECT MASK 2 102.125 24.502 102.205 24.7285 ;
      RECT MASK 2 102.457 24.502 102.537 24.7285 ;
      RECT MASK 2 104.925 24.502 105.005 24.7285 ;
      RECT MASK 2 105.257 24.502 105.337 24.7285 ;
      RECT MASK 2 105.589 24.502 105.669 24.7285 ;
      RECT MASK 2 106.087 24.502 106.167 24.7285 ;
      RECT MASK 2 106.419 24.502 106.499 24.7285 ;
      RECT MASK 2 106.751 24.502 106.831 24.7285 ;
      RECT MASK 2 107.249 24.502 107.329 24.7285 ;
      RECT MASK 2 107.581 24.502 107.661 24.7285 ;
      RECT MASK 2 107.913 24.502 107.993 24.7285 ;
      RECT MASK 2 108.411 24.502 108.491 24.7285 ;
      RECT MASK 2 108.743 24.502 108.823 24.7285 ;
      RECT MASK 2 109.075 24.502 109.155 24.7285 ;
      RECT MASK 2 1.406 24.68 4.69 24.72 ;
      RECT MASK 2 1.406 24.87 4.69 24.91 ;
      RECT MASK 2 5.655 25.167 5.735 25.394 ;
      RECT MASK 2 5.987 25.167 6.067 25.394 ;
      RECT MASK 2 6.319 25.167 6.399 25.394 ;
      RECT MASK 2 6.817 25.167 6.897 25.394 ;
      RECT MASK 2 7.149 25.167 7.229 25.394 ;
      RECT MASK 2 7.481 25.167 7.561 25.394 ;
      RECT MASK 2 7.979 25.167 8.059 25.394 ;
      RECT MASK 2 8.311 25.167 8.391 25.394 ;
      RECT MASK 2 8.643 25.167 8.723 25.394 ;
      RECT MASK 2 9.141 25.167 9.221 25.394 ;
      RECT MASK 2 9.473 25.167 9.553 25.394 ;
      RECT MASK 2 9.805 25.167 9.885 25.394 ;
      RECT MASK 2 12.273 25.167 12.353 25.394 ;
      RECT MASK 2 12.605 25.167 12.685 25.394 ;
      RECT MASK 2 12.937 25.167 13.017 25.394 ;
      RECT MASK 2 13.435 25.167 13.515 25.394 ;
      RECT MASK 2 13.767 25.167 13.847 25.394 ;
      RECT MASK 2 14.099 25.167 14.179 25.394 ;
      RECT MASK 2 14.597 25.167 14.677 25.394 ;
      RECT MASK 2 14.929 25.167 15.009 25.394 ;
      RECT MASK 2 15.261 25.167 15.341 25.394 ;
      RECT MASK 2 15.759 25.167 15.839 25.394 ;
      RECT MASK 2 16.091 25.167 16.171 25.394 ;
      RECT MASK 2 16.423 25.167 16.503 25.394 ;
      RECT MASK 2 18.891 25.167 18.971 25.394 ;
      RECT MASK 2 19.223 25.167 19.303 25.394 ;
      RECT MASK 2 19.555 25.167 19.635 25.394 ;
      RECT MASK 2 20.053 25.167 20.133 25.394 ;
      RECT MASK 2 20.385 25.167 20.465 25.394 ;
      RECT MASK 2 20.717 25.167 20.797 25.394 ;
      RECT MASK 2 21.215 25.167 21.295 25.394 ;
      RECT MASK 2 21.547 25.167 21.627 25.394 ;
      RECT MASK 2 21.879 25.167 21.959 25.394 ;
      RECT MASK 2 22.377 25.167 22.457 25.394 ;
      RECT MASK 2 22.709 25.167 22.789 25.394 ;
      RECT MASK 2 23.041 25.167 23.121 25.394 ;
      RECT MASK 2 25.509 25.167 25.589 25.394 ;
      RECT MASK 2 25.841 25.167 25.921 25.394 ;
      RECT MASK 2 26.173 25.167 26.253 25.394 ;
      RECT MASK 2 26.671 25.167 26.751 25.394 ;
      RECT MASK 2 27.003 25.167 27.083 25.394 ;
      RECT MASK 2 27.335 25.167 27.415 25.394 ;
      RECT MASK 2 27.833 25.167 27.913 25.394 ;
      RECT MASK 2 28.165 25.167 28.245 25.394 ;
      RECT MASK 2 28.497 25.167 28.577 25.394 ;
      RECT MASK 2 28.995 25.167 29.075 25.394 ;
      RECT MASK 2 29.327 25.167 29.407 25.394 ;
      RECT MASK 2 29.659 25.167 29.739 25.394 ;
      RECT MASK 2 32.127 25.167 32.207 25.394 ;
      RECT MASK 2 32.459 25.167 32.539 25.394 ;
      RECT MASK 2 32.791 25.167 32.871 25.394 ;
      RECT MASK 2 33.289 25.167 33.369 25.394 ;
      RECT MASK 2 33.621 25.167 33.701 25.394 ;
      RECT MASK 2 33.953 25.167 34.033 25.394 ;
      RECT MASK 2 34.451 25.167 34.531 25.394 ;
      RECT MASK 2 34.783 25.167 34.863 25.394 ;
      RECT MASK 2 35.115 25.167 35.195 25.394 ;
      RECT MASK 2 35.613 25.167 35.693 25.394 ;
      RECT MASK 2 35.945 25.167 36.025 25.394 ;
      RECT MASK 2 36.277 25.167 36.357 25.394 ;
      RECT MASK 2 38.745 25.167 38.825 25.394 ;
      RECT MASK 2 39.077 25.167 39.157 25.394 ;
      RECT MASK 2 39.409 25.167 39.489 25.394 ;
      RECT MASK 2 39.907 25.167 39.987 25.394 ;
      RECT MASK 2 40.239 25.167 40.319 25.394 ;
      RECT MASK 2 40.571 25.167 40.651 25.394 ;
      RECT MASK 2 41.069 25.167 41.149 25.394 ;
      RECT MASK 2 41.401 25.167 41.481 25.394 ;
      RECT MASK 2 41.733 25.167 41.813 25.394 ;
      RECT MASK 2 42.231 25.167 42.311 25.394 ;
      RECT MASK 2 42.563 25.167 42.643 25.394 ;
      RECT MASK 2 42.895 25.167 42.975 25.394 ;
      RECT MASK 2 45.363 25.167 45.443 25.394 ;
      RECT MASK 2 45.695 25.167 45.775 25.394 ;
      RECT MASK 2 46.027 25.167 46.107 25.394 ;
      RECT MASK 2 46.525 25.167 46.605 25.394 ;
      RECT MASK 2 46.857 25.167 46.937 25.394 ;
      RECT MASK 2 47.189 25.167 47.269 25.394 ;
      RECT MASK 2 47.687 25.167 47.767 25.394 ;
      RECT MASK 2 48.019 25.167 48.099 25.394 ;
      RECT MASK 2 48.351 25.167 48.431 25.394 ;
      RECT MASK 2 48.849 25.167 48.929 25.394 ;
      RECT MASK 2 49.181 25.167 49.261 25.394 ;
      RECT MASK 2 49.513 25.167 49.593 25.394 ;
      RECT MASK 2 51.981 25.167 52.061 25.394 ;
      RECT MASK 2 52.313 25.167 52.393 25.394 ;
      RECT MASK 2 52.645 25.167 52.725 25.394 ;
      RECT MASK 2 53.143 25.167 53.223 25.394 ;
      RECT MASK 2 53.475 25.167 53.555 25.394 ;
      RECT MASK 2 53.807 25.167 53.887 25.394 ;
      RECT MASK 2 54.305 25.167 54.385 25.394 ;
      RECT MASK 2 54.637 25.167 54.717 25.394 ;
      RECT MASK 2 54.969 25.167 55.049 25.394 ;
      RECT MASK 2 55.467 25.167 55.547 25.394 ;
      RECT MASK 2 55.799 25.167 55.879 25.394 ;
      RECT MASK 2 56.131 25.167 56.211 25.394 ;
      RECT MASK 2 58.599 25.167 58.679 25.394 ;
      RECT MASK 2 58.931 25.167 59.011 25.394 ;
      RECT MASK 2 59.263 25.167 59.343 25.394 ;
      RECT MASK 2 59.761 25.167 59.841 25.394 ;
      RECT MASK 2 60.093 25.167 60.173 25.394 ;
      RECT MASK 2 60.425 25.167 60.505 25.394 ;
      RECT MASK 2 60.923 25.167 61.003 25.394 ;
      RECT MASK 2 61.255 25.167 61.335 25.394 ;
      RECT MASK 2 61.587 25.167 61.667 25.394 ;
      RECT MASK 2 62.085 25.167 62.165 25.394 ;
      RECT MASK 2 62.417 25.167 62.497 25.394 ;
      RECT MASK 2 62.749 25.167 62.829 25.394 ;
      RECT MASK 2 65.217 25.167 65.297 25.394 ;
      RECT MASK 2 65.549 25.167 65.629 25.394 ;
      RECT MASK 2 65.881 25.167 65.961 25.394 ;
      RECT MASK 2 66.379 25.167 66.459 25.394 ;
      RECT MASK 2 66.711 25.167 66.791 25.394 ;
      RECT MASK 2 67.043 25.167 67.123 25.394 ;
      RECT MASK 2 67.541 25.167 67.621 25.394 ;
      RECT MASK 2 67.873 25.167 67.953 25.394 ;
      RECT MASK 2 68.205 25.167 68.285 25.394 ;
      RECT MASK 2 68.703 25.167 68.783 25.394 ;
      RECT MASK 2 69.035 25.167 69.115 25.394 ;
      RECT MASK 2 69.367 25.167 69.447 25.394 ;
      RECT MASK 2 71.835 25.167 71.915 25.394 ;
      RECT MASK 2 72.167 25.167 72.247 25.394 ;
      RECT MASK 2 72.499 25.167 72.579 25.394 ;
      RECT MASK 2 72.997 25.167 73.077 25.394 ;
      RECT MASK 2 73.329 25.167 73.409 25.394 ;
      RECT MASK 2 73.661 25.167 73.741 25.394 ;
      RECT MASK 2 74.159 25.167 74.239 25.394 ;
      RECT MASK 2 74.491 25.167 74.571 25.394 ;
      RECT MASK 2 74.823 25.167 74.903 25.394 ;
      RECT MASK 2 75.321 25.167 75.401 25.394 ;
      RECT MASK 2 75.653 25.167 75.733 25.394 ;
      RECT MASK 2 75.985 25.167 76.065 25.394 ;
      RECT MASK 2 78.453 25.167 78.533 25.394 ;
      RECT MASK 2 78.785 25.167 78.865 25.394 ;
      RECT MASK 2 79.117 25.167 79.197 25.394 ;
      RECT MASK 2 79.615 25.167 79.695 25.394 ;
      RECT MASK 2 79.947 25.167 80.027 25.394 ;
      RECT MASK 2 80.279 25.167 80.359 25.394 ;
      RECT MASK 2 80.777 25.167 80.857 25.394 ;
      RECT MASK 2 81.109 25.167 81.189 25.394 ;
      RECT MASK 2 81.441 25.167 81.521 25.394 ;
      RECT MASK 2 81.939 25.167 82.019 25.394 ;
      RECT MASK 2 82.271 25.167 82.351 25.394 ;
      RECT MASK 2 82.603 25.167 82.683 25.394 ;
      RECT MASK 2 85.071 25.167 85.151 25.394 ;
      RECT MASK 2 85.403 25.167 85.483 25.394 ;
      RECT MASK 2 85.735 25.167 85.815 25.394 ;
      RECT MASK 2 86.233 25.167 86.313 25.394 ;
      RECT MASK 2 86.565 25.167 86.645 25.394 ;
      RECT MASK 2 86.897 25.167 86.977 25.394 ;
      RECT MASK 2 87.395 25.167 87.475 25.394 ;
      RECT MASK 2 87.727 25.167 87.807 25.394 ;
      RECT MASK 2 88.059 25.167 88.139 25.394 ;
      RECT MASK 2 88.557 25.167 88.637 25.394 ;
      RECT MASK 2 88.889 25.167 88.969 25.394 ;
      RECT MASK 2 89.221 25.167 89.301 25.394 ;
      RECT MASK 2 91.689 25.167 91.769 25.394 ;
      RECT MASK 2 92.021 25.167 92.101 25.394 ;
      RECT MASK 2 92.353 25.167 92.433 25.394 ;
      RECT MASK 2 92.851 25.167 92.931 25.394 ;
      RECT MASK 2 93.183 25.167 93.263 25.394 ;
      RECT MASK 2 93.515 25.167 93.595 25.394 ;
      RECT MASK 2 94.013 25.167 94.093 25.394 ;
      RECT MASK 2 94.345 25.167 94.425 25.394 ;
      RECT MASK 2 94.677 25.167 94.757 25.394 ;
      RECT MASK 2 95.175 25.167 95.255 25.394 ;
      RECT MASK 2 95.507 25.167 95.587 25.394 ;
      RECT MASK 2 95.839 25.167 95.919 25.394 ;
      RECT MASK 2 98.307 25.167 98.387 25.394 ;
      RECT MASK 2 98.639 25.167 98.719 25.394 ;
      RECT MASK 2 98.971 25.167 99.051 25.394 ;
      RECT MASK 2 99.469 25.167 99.549 25.394 ;
      RECT MASK 2 99.801 25.167 99.881 25.394 ;
      RECT MASK 2 100.133 25.167 100.213 25.394 ;
      RECT MASK 2 100.631 25.167 100.711 25.394 ;
      RECT MASK 2 100.963 25.167 101.043 25.394 ;
      RECT MASK 2 101.295 25.167 101.375 25.394 ;
      RECT MASK 2 101.793 25.167 101.873 25.394 ;
      RECT MASK 2 102.125 25.167 102.205 25.394 ;
      RECT MASK 2 102.457 25.167 102.537 25.394 ;
      RECT MASK 2 104.925 25.167 105.005 25.394 ;
      RECT MASK 2 105.257 25.167 105.337 25.394 ;
      RECT MASK 2 105.589 25.167 105.669 25.394 ;
      RECT MASK 2 106.087 25.167 106.167 25.394 ;
      RECT MASK 2 106.419 25.167 106.499 25.394 ;
      RECT MASK 2 106.751 25.167 106.831 25.394 ;
      RECT MASK 2 107.249 25.167 107.329 25.394 ;
      RECT MASK 2 107.581 25.167 107.661 25.394 ;
      RECT MASK 2 107.913 25.167 107.993 25.394 ;
      RECT MASK 2 108.411 25.167 108.491 25.394 ;
      RECT MASK 2 108.743 25.167 108.823 25.394 ;
      RECT MASK 2 109.075 25.167 109.155 25.394 ;
      RECT MASK 2 5.1135 25.7 110.065 25.74 ;
      RECT MASK 2 5.1135 25.89 110.065 25.93 ;
      RECT MASK 2 1.31 26.21 113.989 26.25 ;
      RECT MASK 2 1.31 26.4 113.989 26.44 ;
      RECT MASK 2 115.539 26.45 126.947 26.49 ;
      RECT MASK 2 115.539 26.64 126.947 26.68 ;
      RECT MASK 2 2.47 26.889 112.442 27.029 ;
      RECT MASK 2 116.08 26.9285 116.3255 26.9685 ;
      RECT MASK 2 126.2895 26.9285 126.487 26.9685 ;
      RECT MASK 2 116.437 27.188 116.497 27.412 ;
      RECT MASK 2 116.769 27.188 116.829 27.412 ;
      RECT MASK 2 117.101 27.188 117.161 27.412 ;
      RECT MASK 2 117.433 27.188 117.493 27.412 ;
      RECT MASK 2 117.765 27.188 117.825 27.412 ;
      RECT MASK 2 118.097 27.188 118.157 27.412 ;
      RECT MASK 2 118.429 27.188 118.489 27.412 ;
      RECT MASK 2 118.761 27.188 118.821 27.412 ;
      RECT MASK 2 119.093 27.188 119.153 27.412 ;
      RECT MASK 2 119.425 27.188 119.485 27.412 ;
      RECT MASK 2 119.757 27.188 119.817 27.412 ;
      RECT MASK 2 120.089 27.188 120.149 27.412 ;
      RECT MASK 2 120.421 27.188 120.481 27.412 ;
      RECT MASK 2 120.753 27.188 120.813 27.412 ;
      RECT MASK 2 121.085 27.188 121.145 27.412 ;
      RECT MASK 2 121.417 27.188 121.477 27.412 ;
      RECT MASK 2 121.749 27.188 121.809 27.412 ;
      RECT MASK 2 122.081 27.188 122.141 27.412 ;
      RECT MASK 2 122.413 27.188 122.473 27.412 ;
      RECT MASK 2 122.745 27.188 122.805 27.412 ;
      RECT MASK 2 123.077 27.188 123.137 27.412 ;
      RECT MASK 2 123.409 27.188 123.469 27.412 ;
      RECT MASK 2 123.741 27.188 123.801 27.412 ;
      RECT MASK 2 124.073 27.188 124.133 27.412 ;
      RECT MASK 2 124.405 27.188 124.465 27.412 ;
      RECT MASK 2 124.737 27.188 124.797 27.412 ;
      RECT MASK 2 125.069 27.188 125.129 27.412 ;
      RECT MASK 2 125.401 27.188 125.461 27.412 ;
      RECT MASK 2 125.733 27.188 125.793 27.412 ;
      RECT MASK 2 126.065 27.188 126.125 27.412 ;
      RECT MASK 2 2.47 27.349 112.442 27.489 ;
      RECT MASK 2 116.08 27.7085 116.356 27.7485 ;
      RECT MASK 2 126.2895 27.7085 126.486 27.7485 ;
      RECT MASK 2 116.437 27.968 116.497 28.192 ;
      RECT MASK 2 116.769 27.968 116.829 28.192 ;
      RECT MASK 2 117.101 27.968 117.161 28.192 ;
      RECT MASK 2 117.433 27.968 117.493 28.192 ;
      RECT MASK 2 117.765 27.968 117.825 28.192 ;
      RECT MASK 2 118.097 27.968 118.157 28.192 ;
      RECT MASK 2 118.429 27.968 118.489 28.192 ;
      RECT MASK 2 118.761 27.968 118.821 28.192 ;
      RECT MASK 2 119.093 27.968 119.153 28.192 ;
      RECT MASK 2 119.425 27.968 119.485 28.192 ;
      RECT MASK 2 119.757 27.968 119.817 28.192 ;
      RECT MASK 2 120.089 27.968 120.149 28.192 ;
      RECT MASK 2 120.421 27.968 120.481 28.192 ;
      RECT MASK 2 120.753 27.968 120.813 28.192 ;
      RECT MASK 2 121.085 27.968 121.145 28.192 ;
      RECT MASK 2 121.417 27.968 121.477 28.192 ;
      RECT MASK 2 121.749 27.968 121.809 28.192 ;
      RECT MASK 2 122.081 27.968 122.141 28.192 ;
      RECT MASK 2 122.413 27.968 122.473 28.192 ;
      RECT MASK 2 122.745 27.968 122.805 28.192 ;
      RECT MASK 2 123.077 27.968 123.137 28.192 ;
      RECT MASK 2 123.409 27.968 123.469 28.192 ;
      RECT MASK 2 123.741 27.968 123.801 28.192 ;
      RECT MASK 2 124.073 27.968 124.133 28.192 ;
      RECT MASK 2 124.405 27.968 124.465 28.192 ;
      RECT MASK 2 124.737 27.968 124.797 28.192 ;
      RECT MASK 2 125.069 27.968 125.129 28.192 ;
      RECT MASK 2 125.401 27.968 125.461 28.192 ;
      RECT MASK 2 125.733 27.968 125.793 28.192 ;
      RECT MASK 2 126.065 27.968 126.125 28.192 ;
      RECT MASK 2 2.47 28.239 4.348 28.379 ;
      RECT MASK 2 4.676 28.239 10.966 28.379 ;
      RECT MASK 2 11.294 28.239 17.584 28.379 ;
      RECT MASK 2 17.912 28.239 24.202 28.379 ;
      RECT MASK 2 24.53 28.239 30.82 28.379 ;
      RECT MASK 2 31.148 28.239 37.438 28.379 ;
      RECT MASK 2 37.766 28.239 44.056 28.379 ;
      RECT MASK 2 44.384 28.239 50.674 28.379 ;
      RECT MASK 2 51.002 28.239 57.292 28.379 ;
      RECT MASK 2 57.62 28.239 63.91 28.379 ;
      RECT MASK 2 64.238 28.239 70.528 28.379 ;
      RECT MASK 2 70.856 28.239 77.146 28.379 ;
      RECT MASK 2 77.474 28.239 83.764 28.379 ;
      RECT MASK 2 84.092 28.239 90.382 28.379 ;
      RECT MASK 2 90.71 28.239 97 28.379 ;
      RECT MASK 2 97.328 28.239 103.618 28.379 ;
      RECT MASK 2 103.946 28.239 110.236 28.379 ;
      RECT MASK 2 110.564 28.239 112.463 28.379 ;
      RECT MASK 2 116.08 28.4885 116.3255 28.5285 ;
      RECT MASK 2 126.2895 28.4885 126.485 28.5285 ;
      RECT MASK 2 2.47 28.699 4.348 28.839 ;
      RECT MASK 2 4.676 28.699 10.966 28.839 ;
      RECT MASK 2 11.294 28.699 17.584 28.839 ;
      RECT MASK 2 17.912 28.699 24.202 28.839 ;
      RECT MASK 2 24.53 28.699 30.82 28.839 ;
      RECT MASK 2 31.148 28.699 37.438 28.839 ;
      RECT MASK 2 37.766 28.699 44.056 28.839 ;
      RECT MASK 2 44.384 28.699 50.674 28.839 ;
      RECT MASK 2 51.002 28.699 57.292 28.839 ;
      RECT MASK 2 57.62 28.699 63.91 28.839 ;
      RECT MASK 2 64.238 28.699 70.528 28.839 ;
      RECT MASK 2 70.856 28.699 77.146 28.839 ;
      RECT MASK 2 77.474 28.699 83.764 28.839 ;
      RECT MASK 2 84.092 28.699 90.382 28.839 ;
      RECT MASK 2 90.71 28.699 97 28.839 ;
      RECT MASK 2 97.328 28.699 103.618 28.839 ;
      RECT MASK 2 103.946 28.699 110.236 28.839 ;
      RECT MASK 2 110.564 28.699 112.463 28.839 ;
      RECT MASK 2 116.437 28.748 116.497 28.972 ;
      RECT MASK 2 116.769 28.748 116.829 28.972 ;
      RECT MASK 2 117.101 28.748 117.161 28.972 ;
      RECT MASK 2 117.433 28.748 117.493 28.972 ;
      RECT MASK 2 117.765 28.748 117.825 28.972 ;
      RECT MASK 2 118.097 28.748 118.157 28.972 ;
      RECT MASK 2 118.429 28.748 118.489 28.972 ;
      RECT MASK 2 118.761 28.748 118.821 28.972 ;
      RECT MASK 2 119.093 28.748 119.153 28.972 ;
      RECT MASK 2 119.425 28.748 119.485 28.972 ;
      RECT MASK 2 119.757 28.748 119.817 28.972 ;
      RECT MASK 2 120.089 28.748 120.149 28.972 ;
      RECT MASK 2 120.421 28.748 120.481 28.972 ;
      RECT MASK 2 120.753 28.748 120.813 28.972 ;
      RECT MASK 2 121.085 28.748 121.145 28.972 ;
      RECT MASK 2 121.417 28.748 121.477 28.972 ;
      RECT MASK 2 121.749 28.748 121.809 28.972 ;
      RECT MASK 2 122.081 28.748 122.141 28.972 ;
      RECT MASK 2 122.413 28.748 122.473 28.972 ;
      RECT MASK 2 122.745 28.748 122.805 28.972 ;
      RECT MASK 2 123.077 28.748 123.137 28.972 ;
      RECT MASK 2 123.409 28.748 123.469 28.972 ;
      RECT MASK 2 123.741 28.748 123.801 28.972 ;
      RECT MASK 2 124.073 28.748 124.133 28.972 ;
      RECT MASK 2 124.405 28.748 124.465 28.972 ;
      RECT MASK 2 124.737 28.748 124.797 28.972 ;
      RECT MASK 2 125.069 28.748 125.129 28.972 ;
      RECT MASK 2 125.401 28.748 125.461 28.972 ;
      RECT MASK 2 125.733 28.748 125.793 28.972 ;
      RECT MASK 2 126.065 28.748 126.125 28.972 ;
      RECT MASK 2 116.08 29.2685 116.3255 29.3085 ;
      RECT MASK 2 126.2895 29.2685 126.483 29.3085 ;
      RECT MASK 2 116.437 29.528 116.497 29.752 ;
      RECT MASK 2 116.769 29.528 116.829 29.752 ;
      RECT MASK 2 117.101 29.528 117.161 29.752 ;
      RECT MASK 2 117.433 29.528 117.493 29.752 ;
      RECT MASK 2 117.765 29.528 117.825 29.752 ;
      RECT MASK 2 118.097 29.528 118.157 29.752 ;
      RECT MASK 2 118.429 29.528 118.489 29.752 ;
      RECT MASK 2 118.761 29.528 118.821 29.752 ;
      RECT MASK 2 119.093 29.528 119.153 29.752 ;
      RECT MASK 2 119.425 29.528 119.485 29.752 ;
      RECT MASK 2 119.757 29.528 119.817 29.752 ;
      RECT MASK 2 120.089 29.528 120.149 29.752 ;
      RECT MASK 2 120.421 29.528 120.481 29.752 ;
      RECT MASK 2 120.753 29.528 120.813 29.752 ;
      RECT MASK 2 121.085 29.528 121.145 29.752 ;
      RECT MASK 2 121.417 29.528 121.477 29.752 ;
      RECT MASK 2 121.749 29.528 121.809 29.752 ;
      RECT MASK 2 122.081 29.528 122.141 29.752 ;
      RECT MASK 2 122.413 29.528 122.473 29.752 ;
      RECT MASK 2 122.745 29.528 122.805 29.752 ;
      RECT MASK 2 123.077 29.528 123.137 29.752 ;
      RECT MASK 2 123.409 29.528 123.469 29.752 ;
      RECT MASK 2 123.741 29.528 123.801 29.752 ;
      RECT MASK 2 124.073 29.528 124.133 29.752 ;
      RECT MASK 2 124.405 29.528 124.465 29.752 ;
      RECT MASK 2 124.737 29.528 124.797 29.752 ;
      RECT MASK 2 125.069 29.528 125.129 29.752 ;
      RECT MASK 2 125.401 29.528 125.461 29.752 ;
      RECT MASK 2 125.733 29.528 125.793 29.752 ;
      RECT MASK 2 126.065 29.528 126.125 29.752 ;
      RECT MASK 2 2.47 29.589 4.348 29.729 ;
      RECT MASK 2 4.676 29.589 10.966 29.729 ;
      RECT MASK 2 11.294 29.589 17.584 29.729 ;
      RECT MASK 2 17.912 29.589 24.202 29.729 ;
      RECT MASK 2 24.53 29.589 30.82 29.729 ;
      RECT MASK 2 31.148 29.589 37.438 29.729 ;
      RECT MASK 2 37.766 29.589 44.056 29.729 ;
      RECT MASK 2 44.384 29.589 50.674 29.729 ;
      RECT MASK 2 51.002 29.589 57.292 29.729 ;
      RECT MASK 2 57.62 29.589 63.91 29.729 ;
      RECT MASK 2 64.238 29.589 70.528 29.729 ;
      RECT MASK 2 70.856 29.589 77.146 29.729 ;
      RECT MASK 2 77.474 29.589 83.764 29.729 ;
      RECT MASK 2 84.092 29.589 90.382 29.729 ;
      RECT MASK 2 90.71 29.589 97 29.729 ;
      RECT MASK 2 97.328 29.589 103.618 29.729 ;
      RECT MASK 2 103.946 29.589 110.236 29.729 ;
      RECT MASK 2 110.564 29.589 112.463 29.729 ;
      RECT MASK 2 2.47 30.049 4.348 30.189 ;
      RECT MASK 2 4.676 30.049 10.966 30.189 ;
      RECT MASK 2 11.294 30.049 17.584 30.189 ;
      RECT MASK 2 17.912 30.049 24.202 30.189 ;
      RECT MASK 2 24.53 30.049 30.82 30.189 ;
      RECT MASK 2 31.148 30.049 37.438 30.189 ;
      RECT MASK 2 37.766 30.049 44.056 30.189 ;
      RECT MASK 2 44.384 30.049 50.674 30.189 ;
      RECT MASK 2 51.002 30.049 57.292 30.189 ;
      RECT MASK 2 57.62 30.049 63.91 30.189 ;
      RECT MASK 2 64.238 30.049 70.528 30.189 ;
      RECT MASK 2 70.856 30.049 77.146 30.189 ;
      RECT MASK 2 77.474 30.049 83.764 30.189 ;
      RECT MASK 2 84.092 30.049 90.382 30.189 ;
      RECT MASK 2 90.71 30.049 97 30.189 ;
      RECT MASK 2 97.328 30.049 103.618 30.189 ;
      RECT MASK 2 103.946 30.049 110.236 30.189 ;
      RECT MASK 2 110.564 30.049 112.463 30.189 ;
      RECT MASK 2 115.539 30.26 126.947 30.3 ;
      RECT MASK 2 115.539 30.45 126.947 30.49 ;
      RECT MASK 2 2.47 30.939 4.348 31.079 ;
      RECT MASK 2 4.676 30.939 10.966 31.079 ;
      RECT MASK 2 11.294 30.939 17.584 31.079 ;
      RECT MASK 2 17.912 30.939 24.202 31.079 ;
      RECT MASK 2 24.53 30.939 30.82 31.079 ;
      RECT MASK 2 31.148 30.939 37.438 31.079 ;
      RECT MASK 2 37.766 30.939 44.056 31.079 ;
      RECT MASK 2 44.384 30.939 50.674 31.079 ;
      RECT MASK 2 51.002 30.939 57.292 31.079 ;
      RECT MASK 2 57.62 30.939 63.91 31.079 ;
      RECT MASK 2 64.238 30.939 70.528 31.079 ;
      RECT MASK 2 70.856 30.939 77.146 31.079 ;
      RECT MASK 2 77.474 30.939 83.764 31.079 ;
      RECT MASK 2 84.092 30.939 90.382 31.079 ;
      RECT MASK 2 90.71 30.939 97 31.079 ;
      RECT MASK 2 97.328 30.939 103.618 31.079 ;
      RECT MASK 2 103.946 30.939 110.236 31.079 ;
      RECT MASK 2 110.564 30.939 112.463 31.079 ;
      RECT MASK 2 113.869 31.19 129.1075 31.23 ;
      RECT MASK 2 113.869 31.38 129.1075 31.42 ;
      RECT MASK 2 2.47 31.399 4.348 31.539 ;
      RECT MASK 2 4.676 31.399 10.966 31.539 ;
      RECT MASK 2 11.294 31.399 17.584 31.539 ;
      RECT MASK 2 17.912 31.399 24.202 31.539 ;
      RECT MASK 2 24.53 31.399 30.82 31.539 ;
      RECT MASK 2 31.148 31.399 37.438 31.539 ;
      RECT MASK 2 37.766 31.399 44.056 31.539 ;
      RECT MASK 2 44.384 31.399 50.674 31.539 ;
      RECT MASK 2 51.002 31.399 57.292 31.539 ;
      RECT MASK 2 57.62 31.399 63.91 31.539 ;
      RECT MASK 2 64.238 31.399 70.528 31.539 ;
      RECT MASK 2 70.856 31.399 77.146 31.539 ;
      RECT MASK 2 77.474 31.399 83.764 31.539 ;
      RECT MASK 2 84.092 31.399 90.382 31.539 ;
      RECT MASK 2 90.71 31.399 97 31.539 ;
      RECT MASK 2 97.328 31.399 103.618 31.539 ;
      RECT MASK 2 103.946 31.399 110.236 31.539 ;
      RECT MASK 2 110.564 31.399 112.463 31.539 ;
      RECT MASK 2 2.47 32.289 4.348 32.429 ;
      RECT MASK 2 4.676 32.289 10.966 32.429 ;
      RECT MASK 2 11.294 32.289 17.584 32.429 ;
      RECT MASK 2 17.912 32.289 24.202 32.429 ;
      RECT MASK 2 24.53 32.289 30.82 32.429 ;
      RECT MASK 2 31.148 32.289 37.438 32.429 ;
      RECT MASK 2 37.766 32.289 44.056 32.429 ;
      RECT MASK 2 44.384 32.289 50.674 32.429 ;
      RECT MASK 2 51.002 32.289 57.292 32.429 ;
      RECT MASK 2 57.62 32.289 63.91 32.429 ;
      RECT MASK 2 64.238 32.289 70.528 32.429 ;
      RECT MASK 2 70.856 32.289 77.146 32.429 ;
      RECT MASK 2 77.474 32.289 83.764 32.429 ;
      RECT MASK 2 84.092 32.289 90.382 32.429 ;
      RECT MASK 2 90.71 32.289 97 32.429 ;
      RECT MASK 2 97.328 32.289 103.618 32.429 ;
      RECT MASK 2 103.946 32.289 110.236 32.429 ;
      RECT MASK 2 110.564 32.289 116.854 32.429 ;
      RECT MASK 2 117.182 32.289 127.884 32.429 ;
      RECT MASK 2 2.47 32.749 4.348 32.889 ;
      RECT MASK 2 4.676 32.749 10.966 32.889 ;
      RECT MASK 2 11.294 32.749 17.584 32.889 ;
      RECT MASK 2 17.912 32.749 24.202 32.889 ;
      RECT MASK 2 24.53 32.749 30.82 32.889 ;
      RECT MASK 2 31.148 32.749 37.438 32.889 ;
      RECT MASK 2 37.766 32.749 44.056 32.889 ;
      RECT MASK 2 44.384 32.749 50.674 32.889 ;
      RECT MASK 2 51.002 32.749 57.292 32.889 ;
      RECT MASK 2 57.62 32.749 63.91 32.889 ;
      RECT MASK 2 64.238 32.749 70.528 32.889 ;
      RECT MASK 2 70.856 32.749 77.146 32.889 ;
      RECT MASK 2 77.474 32.749 83.764 32.889 ;
      RECT MASK 2 84.092 32.749 90.382 32.889 ;
      RECT MASK 2 90.71 32.749 97 32.889 ;
      RECT MASK 2 97.328 32.749 103.618 32.889 ;
      RECT MASK 2 103.946 32.749 110.236 32.889 ;
      RECT MASK 2 110.564 32.749 116.854 32.889 ;
      RECT MASK 2 117.182 32.749 127.884 32.889 ;
      RECT MASK 2 1.9425 33.29 41.8765 33.33 ;
      RECT MASK 2 42.6605 33.29 82.5945 33.33 ;
      RECT MASK 2 83.4005 33.29 128.3145 33.33 ;
      RECT MASK 2 1.9425 33.45 41.8765 33.49 ;
      RECT MASK 2 42.6605 33.45 82.5945 33.49 ;
      RECT MASK 2 83.4005 33.45 128.3145 33.49 ;
      RECT MASK 2 1.9425 33.71 41.8765 33.75 ;
      RECT MASK 2 42.6605 33.71 82.5945 33.75 ;
      RECT MASK 2 83.4005 33.71 128.3145 33.75 ;
      RECT MASK 2 1.9425 33.87 41.8765 33.91 ;
      RECT MASK 2 42.6605 33.87 82.5945 33.91 ;
      RECT MASK 2 83.4005 33.87 128.3145 33.91 ;
      RECT MASK 2 2.47 34.329 4.348 34.469 ;
      RECT MASK 2 4.676 34.329 10.966 34.469 ;
      RECT MASK 2 11.294 34.329 17.584 34.469 ;
      RECT MASK 2 17.912 34.329 24.202 34.469 ;
      RECT MASK 2 24.53 34.329 30.82 34.469 ;
      RECT MASK 2 31.148 34.329 37.438 34.469 ;
      RECT MASK 2 37.766 34.329 44.056 34.469 ;
      RECT MASK 2 44.384 34.329 50.674 34.469 ;
      RECT MASK 2 51.002 34.329 57.292 34.469 ;
      RECT MASK 2 57.62 34.329 63.91 34.469 ;
      RECT MASK 2 64.238 34.329 70.528 34.469 ;
      RECT MASK 2 70.856 34.329 77.146 34.469 ;
      RECT MASK 2 77.474 34.329 83.764 34.469 ;
      RECT MASK 2 84.092 34.329 90.382 34.469 ;
      RECT MASK 2 90.71 34.329 97 34.469 ;
      RECT MASK 2 97.328 34.329 103.618 34.469 ;
      RECT MASK 2 103.946 34.329 110.236 34.469 ;
      RECT MASK 2 110.564 34.329 116.854 34.469 ;
      RECT MASK 2 117.182 34.329 127.884 34.469 ;
      RECT MASK 2 2.47 34.789 4.348 34.929 ;
      RECT MASK 2 4.676 34.789 10.966 34.929 ;
      RECT MASK 2 11.294 34.789 17.584 34.929 ;
      RECT MASK 2 17.912 34.789 24.202 34.929 ;
      RECT MASK 2 24.53 34.789 30.82 34.929 ;
      RECT MASK 2 31.148 34.789 37.438 34.929 ;
      RECT MASK 2 37.766 34.789 44.056 34.929 ;
      RECT MASK 2 44.384 34.789 50.674 34.929 ;
      RECT MASK 2 51.002 34.789 57.292 34.929 ;
      RECT MASK 2 57.62 34.789 63.91 34.929 ;
      RECT MASK 2 64.238 34.789 70.528 34.929 ;
      RECT MASK 2 70.856 34.789 77.146 34.929 ;
      RECT MASK 2 77.474 34.789 83.764 34.929 ;
      RECT MASK 2 84.092 34.789 90.382 34.929 ;
      RECT MASK 2 90.71 34.789 97 34.929 ;
      RECT MASK 2 97.328 34.789 103.618 34.929 ;
      RECT MASK 2 103.946 34.789 110.236 34.929 ;
      RECT MASK 2 110.564 34.789 116.854 34.929 ;
      RECT MASK 2 117.182 34.789 127.884 34.929 ;
      RECT MASK 2 2.47 35.679 4.348 35.819 ;
      RECT MASK 2 4.676 35.679 10.966 35.819 ;
      RECT MASK 2 11.294 35.679 17.584 35.819 ;
      RECT MASK 2 17.912 35.679 24.202 35.819 ;
      RECT MASK 2 24.53 35.679 30.82 35.819 ;
      RECT MASK 2 31.148 35.679 37.438 35.819 ;
      RECT MASK 2 37.766 35.679 44.056 35.819 ;
      RECT MASK 2 44.384 35.679 50.674 35.819 ;
      RECT MASK 2 51.002 35.679 57.292 35.819 ;
      RECT MASK 2 57.62 35.679 63.91 35.819 ;
      RECT MASK 2 64.238 35.679 70.528 35.819 ;
      RECT MASK 2 70.856 35.679 77.146 35.819 ;
      RECT MASK 2 77.474 35.679 83.764 35.819 ;
      RECT MASK 2 84.092 35.679 90.382 35.819 ;
      RECT MASK 2 90.71 35.679 97 35.819 ;
      RECT MASK 2 97.328 35.679 103.618 35.819 ;
      RECT MASK 2 103.946 35.679 110.236 35.819 ;
      RECT MASK 2 110.564 35.679 116.854 35.819 ;
      RECT MASK 2 117.182 35.679 127.884 35.819 ;
      RECT MASK 2 2.47 36.139 4.348 36.279 ;
      RECT MASK 2 4.676 36.139 10.966 36.279 ;
      RECT MASK 2 11.294 36.139 17.584 36.279 ;
      RECT MASK 2 17.912 36.139 24.202 36.279 ;
      RECT MASK 2 24.53 36.139 30.82 36.279 ;
      RECT MASK 2 31.148 36.139 37.438 36.279 ;
      RECT MASK 2 37.766 36.139 44.056 36.279 ;
      RECT MASK 2 44.384 36.139 50.674 36.279 ;
      RECT MASK 2 51.002 36.139 57.292 36.279 ;
      RECT MASK 2 57.62 36.139 63.91 36.279 ;
      RECT MASK 2 64.238 36.139 70.528 36.279 ;
      RECT MASK 2 70.856 36.139 77.146 36.279 ;
      RECT MASK 2 77.474 36.139 83.764 36.279 ;
      RECT MASK 2 84.092 36.139 90.382 36.279 ;
      RECT MASK 2 90.71 36.139 97 36.279 ;
      RECT MASK 2 97.328 36.139 103.618 36.279 ;
      RECT MASK 2 103.946 36.139 110.236 36.279 ;
      RECT MASK 2 110.564 36.139 116.854 36.279 ;
      RECT MASK 2 117.182 36.139 127.884 36.279 ;
      RECT MASK 2 2.47 37.029 4.348 37.169 ;
      RECT MASK 2 4.676 37.029 10.966 37.169 ;
      RECT MASK 2 11.294 37.029 17.584 37.169 ;
      RECT MASK 2 17.912 37.029 24.202 37.169 ;
      RECT MASK 2 24.53 37.029 30.82 37.169 ;
      RECT MASK 2 31.148 37.029 37.438 37.169 ;
      RECT MASK 2 37.766 37.029 44.056 37.169 ;
      RECT MASK 2 44.384 37.029 50.674 37.169 ;
      RECT MASK 2 51.002 37.029 57.292 37.169 ;
      RECT MASK 2 57.62 37.029 63.91 37.169 ;
      RECT MASK 2 64.238 37.029 70.528 37.169 ;
      RECT MASK 2 70.856 37.029 77.146 37.169 ;
      RECT MASK 2 77.474 37.029 83.764 37.169 ;
      RECT MASK 2 84.092 37.029 90.382 37.169 ;
      RECT MASK 2 90.71 37.029 97 37.169 ;
      RECT MASK 2 97.328 37.029 103.618 37.169 ;
      RECT MASK 2 103.946 37.029 110.236 37.169 ;
      RECT MASK 2 110.564 37.029 116.854 37.169 ;
      RECT MASK 2 117.182 37.029 127.884 37.169 ;
      RECT MASK 2 2.47 37.489 4.348 37.629 ;
      RECT MASK 2 4.676 37.489 10.966 37.629 ;
      RECT MASK 2 11.294 37.489 17.584 37.629 ;
      RECT MASK 2 17.912 37.489 24.202 37.629 ;
      RECT MASK 2 24.53 37.489 30.82 37.629 ;
      RECT MASK 2 31.148 37.489 37.438 37.629 ;
      RECT MASK 2 37.766 37.489 44.056 37.629 ;
      RECT MASK 2 44.384 37.489 50.674 37.629 ;
      RECT MASK 2 51.002 37.489 57.292 37.629 ;
      RECT MASK 2 57.62 37.489 63.91 37.629 ;
      RECT MASK 2 64.238 37.489 70.528 37.629 ;
      RECT MASK 2 70.856 37.489 77.146 37.629 ;
      RECT MASK 2 77.474 37.489 83.764 37.629 ;
      RECT MASK 2 84.092 37.489 90.382 37.629 ;
      RECT MASK 2 90.71 37.489 97 37.629 ;
      RECT MASK 2 97.328 37.489 103.618 37.629 ;
      RECT MASK 2 103.946 37.489 110.236 37.629 ;
      RECT MASK 2 110.564 37.489 116.854 37.629 ;
      RECT MASK 2 117.182 37.489 127.884 37.629 ;
      RECT MASK 2 2.47 38.379 4.348 38.519 ;
      RECT MASK 2 4.676 38.379 10.966 38.519 ;
      RECT MASK 2 11.294 38.379 17.584 38.519 ;
      RECT MASK 2 17.912 38.379 24.202 38.519 ;
      RECT MASK 2 24.53 38.379 30.82 38.519 ;
      RECT MASK 2 31.148 38.379 37.438 38.519 ;
      RECT MASK 2 37.766 38.379 44.056 38.519 ;
      RECT MASK 2 44.384 38.379 50.674 38.519 ;
      RECT MASK 2 51.002 38.379 57.292 38.519 ;
      RECT MASK 2 57.62 38.379 63.91 38.519 ;
      RECT MASK 2 64.238 38.379 70.528 38.519 ;
      RECT MASK 2 70.856 38.379 77.146 38.519 ;
      RECT MASK 2 77.474 38.379 83.764 38.519 ;
      RECT MASK 2 84.092 38.379 90.382 38.519 ;
      RECT MASK 2 90.71 38.379 97 38.519 ;
      RECT MASK 2 97.328 38.379 103.618 38.519 ;
      RECT MASK 2 103.946 38.379 110.236 38.519 ;
      RECT MASK 2 110.564 38.379 116.854 38.519 ;
      RECT MASK 2 117.182 38.379 127.884 38.519 ;
      RECT MASK 2 2.47 38.839 4.348 38.979 ;
      RECT MASK 2 4.676 38.839 10.966 38.979 ;
      RECT MASK 2 11.294 38.839 17.584 38.979 ;
      RECT MASK 2 17.912 38.839 24.202 38.979 ;
      RECT MASK 2 24.53 38.839 30.82 38.979 ;
      RECT MASK 2 31.148 38.839 37.438 38.979 ;
      RECT MASK 2 37.766 38.839 44.056 38.979 ;
      RECT MASK 2 44.384 38.839 50.674 38.979 ;
      RECT MASK 2 51.002 38.839 57.292 38.979 ;
      RECT MASK 2 57.62 38.839 63.91 38.979 ;
      RECT MASK 2 64.238 38.839 70.528 38.979 ;
      RECT MASK 2 70.856 38.839 77.146 38.979 ;
      RECT MASK 2 77.474 38.839 83.764 38.979 ;
      RECT MASK 2 84.092 38.839 90.382 38.979 ;
      RECT MASK 2 90.71 38.839 97 38.979 ;
      RECT MASK 2 97.328 38.839 103.618 38.979 ;
      RECT MASK 2 103.946 38.839 110.236 38.979 ;
      RECT MASK 2 110.564 38.839 116.854 38.979 ;
      RECT MASK 2 117.182 38.839 127.884 38.979 ;
      RECT MASK 2 1.9425 39.38 41.8765 39.42 ;
      RECT MASK 2 42.6605 39.38 82.5945 39.42 ;
      RECT MASK 2 83.4005 39.38 128.3145 39.42 ;
      RECT MASK 2 1.9425 39.54 41.8765 39.58 ;
      RECT MASK 2 42.6605 39.54 82.5945 39.58 ;
      RECT MASK 2 83.4005 39.54 128.3145 39.58 ;
      RECT MASK 2 1.9425 39.8 41.8765 39.84 ;
      RECT MASK 2 42.6605 39.8 82.5945 39.84 ;
      RECT MASK 2 83.4005 39.8 128.3145 39.84 ;
      RECT MASK 2 1.9425 39.96 41.8765 40 ;
      RECT MASK 2 42.6605 39.96 82.5945 40 ;
      RECT MASK 2 83.4005 39.96 128.3145 40 ;
      RECT MASK 2 2.47 40.449 4.348 40.589 ;
      RECT MASK 2 4.676 40.449 10.966 40.589 ;
      RECT MASK 2 11.294 40.449 17.584 40.589 ;
      RECT MASK 2 17.912 40.449 24.202 40.589 ;
      RECT MASK 2 24.53 40.449 30.82 40.589 ;
      RECT MASK 2 31.148 40.449 37.438 40.589 ;
      RECT MASK 2 37.766 40.449 44.056 40.589 ;
      RECT MASK 2 44.384 40.449 50.674 40.589 ;
      RECT MASK 2 51.002 40.449 57.292 40.589 ;
      RECT MASK 2 57.62 40.449 63.91 40.589 ;
      RECT MASK 2 64.238 40.449 70.528 40.589 ;
      RECT MASK 2 70.856 40.449 77.146 40.589 ;
      RECT MASK 2 77.474 40.449 83.764 40.589 ;
      RECT MASK 2 84.092 40.449 90.382 40.589 ;
      RECT MASK 2 90.71 40.449 97 40.589 ;
      RECT MASK 2 97.328 40.449 103.618 40.589 ;
      RECT MASK 2 103.946 40.449 110.236 40.589 ;
      RECT MASK 2 110.564 40.449 116.854 40.589 ;
      RECT MASK 2 117.182 40.449 127.884 40.589 ;
      RECT MASK 2 2.47 40.909 4.348 41.049 ;
      RECT MASK 2 4.676 40.909 10.966 41.049 ;
      RECT MASK 2 11.294 40.909 17.584 41.049 ;
      RECT MASK 2 17.912 40.909 24.202 41.049 ;
      RECT MASK 2 24.53 40.909 30.82 41.049 ;
      RECT MASK 2 31.148 40.909 37.438 41.049 ;
      RECT MASK 2 37.766 40.909 44.056 41.049 ;
      RECT MASK 2 44.384 40.909 50.674 41.049 ;
      RECT MASK 2 51.002 40.909 57.292 41.049 ;
      RECT MASK 2 57.62 40.909 63.91 41.049 ;
      RECT MASK 2 64.238 40.909 70.528 41.049 ;
      RECT MASK 2 70.856 40.909 77.146 41.049 ;
      RECT MASK 2 77.474 40.909 83.764 41.049 ;
      RECT MASK 2 84.092 40.909 90.382 41.049 ;
      RECT MASK 2 90.71 40.909 97 41.049 ;
      RECT MASK 2 97.328 40.909 103.618 41.049 ;
      RECT MASK 2 103.946 40.909 110.236 41.049 ;
      RECT MASK 2 110.564 40.909 116.854 41.049 ;
      RECT MASK 2 117.182 40.909 127.884 41.049 ;
      RECT MASK 2 2.47 41.799 4.348 41.939 ;
      RECT MASK 2 4.676 41.799 10.966 41.939 ;
      RECT MASK 2 11.294 41.799 17.584 41.939 ;
      RECT MASK 2 17.912 41.799 24.202 41.939 ;
      RECT MASK 2 24.53 41.799 30.82 41.939 ;
      RECT MASK 2 31.148 41.799 37.438 41.939 ;
      RECT MASK 2 37.766 41.799 44.056 41.939 ;
      RECT MASK 2 44.384 41.799 50.674 41.939 ;
      RECT MASK 2 51.002 41.799 57.292 41.939 ;
      RECT MASK 2 57.62 41.799 63.91 41.939 ;
      RECT MASK 2 64.238 41.799 70.528 41.939 ;
      RECT MASK 2 70.856 41.799 77.146 41.939 ;
      RECT MASK 2 77.474 41.799 83.764 41.939 ;
      RECT MASK 2 84.092 41.799 90.382 41.939 ;
      RECT MASK 2 90.71 41.799 97 41.939 ;
      RECT MASK 2 97.328 41.799 103.618 41.939 ;
      RECT MASK 2 103.946 41.799 110.236 41.939 ;
      RECT MASK 2 110.564 41.799 116.854 41.939 ;
      RECT MASK 2 117.182 41.799 127.884 41.939 ;
      RECT MASK 2 2.47 42.259 4.348 42.399 ;
      RECT MASK 2 4.676 42.259 10.966 42.399 ;
      RECT MASK 2 11.294 42.259 17.584 42.399 ;
      RECT MASK 2 17.912 42.259 24.202 42.399 ;
      RECT MASK 2 24.53 42.259 30.82 42.399 ;
      RECT MASK 2 31.148 42.259 37.438 42.399 ;
      RECT MASK 2 37.766 42.259 44.056 42.399 ;
      RECT MASK 2 44.384 42.259 50.674 42.399 ;
      RECT MASK 2 51.002 42.259 57.292 42.399 ;
      RECT MASK 2 57.62 42.259 63.91 42.399 ;
      RECT MASK 2 64.238 42.259 70.528 42.399 ;
      RECT MASK 2 70.856 42.259 77.146 42.399 ;
      RECT MASK 2 77.474 42.259 83.764 42.399 ;
      RECT MASK 2 84.092 42.259 90.382 42.399 ;
      RECT MASK 2 90.71 42.259 97 42.399 ;
      RECT MASK 2 97.328 42.259 103.618 42.399 ;
      RECT MASK 2 103.946 42.259 110.236 42.399 ;
      RECT MASK 2 110.564 42.259 116.854 42.399 ;
      RECT MASK 2 117.182 42.259 127.884 42.399 ;
      RECT MASK 2 2.47 43.149 4.348 43.289 ;
      RECT MASK 2 4.676 43.149 10.966 43.289 ;
      RECT MASK 2 11.294 43.149 17.584 43.289 ;
      RECT MASK 2 17.912 43.149 24.202 43.289 ;
      RECT MASK 2 24.53 43.149 30.82 43.289 ;
      RECT MASK 2 31.148 43.149 37.438 43.289 ;
      RECT MASK 2 37.766 43.149 44.056 43.289 ;
      RECT MASK 2 44.384 43.149 50.674 43.289 ;
      RECT MASK 2 51.002 43.149 57.292 43.289 ;
      RECT MASK 2 57.62 43.149 63.91 43.289 ;
      RECT MASK 2 64.238 43.149 70.528 43.289 ;
      RECT MASK 2 70.856 43.149 77.146 43.289 ;
      RECT MASK 2 77.474 43.149 83.764 43.289 ;
      RECT MASK 2 84.092 43.149 90.382 43.289 ;
      RECT MASK 2 90.71 43.149 97 43.289 ;
      RECT MASK 2 97.328 43.149 103.618 43.289 ;
      RECT MASK 2 103.946 43.149 110.236 43.289 ;
      RECT MASK 2 110.564 43.149 116.854 43.289 ;
      RECT MASK 2 117.182 43.149 127.884 43.289 ;
      RECT MASK 2 2.47 43.609 4.348 43.749 ;
      RECT MASK 2 4.676 43.609 10.966 43.749 ;
      RECT MASK 2 11.294 43.609 17.584 43.749 ;
      RECT MASK 2 17.912 43.609 24.202 43.749 ;
      RECT MASK 2 24.53 43.609 30.82 43.749 ;
      RECT MASK 2 31.148 43.609 37.438 43.749 ;
      RECT MASK 2 37.766 43.609 44.056 43.749 ;
      RECT MASK 2 44.384 43.609 50.674 43.749 ;
      RECT MASK 2 51.002 43.609 57.292 43.749 ;
      RECT MASK 2 57.62 43.609 63.91 43.749 ;
      RECT MASK 2 64.238 43.609 70.528 43.749 ;
      RECT MASK 2 70.856 43.609 77.146 43.749 ;
      RECT MASK 2 77.474 43.609 83.764 43.749 ;
      RECT MASK 2 84.092 43.609 90.382 43.749 ;
      RECT MASK 2 90.71 43.609 97 43.749 ;
      RECT MASK 2 97.328 43.609 103.618 43.749 ;
      RECT MASK 2 103.946 43.609 110.236 43.749 ;
      RECT MASK 2 110.564 43.609 116.854 43.749 ;
      RECT MASK 2 117.182 43.609 127.884 43.749 ;
      RECT MASK 2 2.47 44.499 4.348 44.639 ;
      RECT MASK 2 4.676 44.499 10.966 44.639 ;
      RECT MASK 2 11.294 44.499 17.584 44.639 ;
      RECT MASK 2 17.912 44.499 24.202 44.639 ;
      RECT MASK 2 24.53 44.499 30.82 44.639 ;
      RECT MASK 2 31.148 44.499 37.438 44.639 ;
      RECT MASK 2 37.766 44.499 44.056 44.639 ;
      RECT MASK 2 44.384 44.499 50.674 44.639 ;
      RECT MASK 2 51.002 44.499 57.292 44.639 ;
      RECT MASK 2 57.62 44.499 63.91 44.639 ;
      RECT MASK 2 64.238 44.499 70.528 44.639 ;
      RECT MASK 2 70.856 44.499 77.146 44.639 ;
      RECT MASK 2 77.474 44.499 83.764 44.639 ;
      RECT MASK 2 84.092 44.499 90.382 44.639 ;
      RECT MASK 2 90.71 44.499 97 44.639 ;
      RECT MASK 2 97.328 44.499 103.618 44.639 ;
      RECT MASK 2 103.946 44.499 110.236 44.639 ;
      RECT MASK 2 110.564 44.499 116.854 44.639 ;
      RECT MASK 2 117.182 44.499 127.884 44.639 ;
      RECT MASK 2 2.47 44.959 4.348 45.099 ;
      RECT MASK 2 4.676 44.959 10.966 45.099 ;
      RECT MASK 2 11.294 44.959 17.584 45.099 ;
      RECT MASK 2 17.912 44.959 24.202 45.099 ;
      RECT MASK 2 24.53 44.959 30.82 45.099 ;
      RECT MASK 2 31.148 44.959 37.438 45.099 ;
      RECT MASK 2 37.766 44.959 44.056 45.099 ;
      RECT MASK 2 44.384 44.959 50.674 45.099 ;
      RECT MASK 2 51.002 44.959 57.292 45.099 ;
      RECT MASK 2 57.62 44.959 63.91 45.099 ;
      RECT MASK 2 64.238 44.959 70.528 45.099 ;
      RECT MASK 2 70.856 44.959 77.146 45.099 ;
      RECT MASK 2 77.474 44.959 83.764 45.099 ;
      RECT MASK 2 84.092 44.959 90.382 45.099 ;
      RECT MASK 2 90.71 44.959 97 45.099 ;
      RECT MASK 2 97.328 44.959 103.618 45.099 ;
      RECT MASK 2 103.946 44.959 110.236 45.099 ;
      RECT MASK 2 110.564 44.959 116.854 45.099 ;
      RECT MASK 2 117.182 44.959 127.884 45.099 ;
      RECT MASK 2 1.9425 45.5 41.8765 45.54 ;
      RECT MASK 2 42.6605 45.5 82.5945 45.54 ;
      RECT MASK 2 83.4005 45.5 128.3145 45.54 ;
      RECT MASK 2 1.9425 45.66 41.8765 45.7 ;
      RECT MASK 2 42.6605 45.66 82.5945 45.7 ;
      RECT MASK 2 83.4005 45.66 128.3145 45.7 ;
      RECT MASK 2 1.9425 45.92 41.8765 45.96 ;
      RECT MASK 2 42.6605 45.92 82.5945 45.96 ;
      RECT MASK 2 83.4005 45.92 128.3145 45.96 ;
      RECT MASK 2 1.9425 46.08 41.8765 46.12 ;
      RECT MASK 2 42.6605 46.08 82.5945 46.12 ;
      RECT MASK 2 83.4005 46.08 128.3145 46.12 ;
      RECT MASK 2 2.47 46.569 4.348 46.709 ;
      RECT MASK 2 4.676 46.569 10.966 46.709 ;
      RECT MASK 2 11.294 46.569 17.584 46.709 ;
      RECT MASK 2 17.912 46.569 24.202 46.709 ;
      RECT MASK 2 24.53 46.569 30.82 46.709 ;
      RECT MASK 2 31.148 46.569 37.438 46.709 ;
      RECT MASK 2 37.766 46.569 44.056 46.709 ;
      RECT MASK 2 44.384 46.569 50.674 46.709 ;
      RECT MASK 2 51.002 46.569 57.292 46.709 ;
      RECT MASK 2 57.62 46.569 63.91 46.709 ;
      RECT MASK 2 64.238 46.569 70.528 46.709 ;
      RECT MASK 2 70.856 46.569 77.146 46.709 ;
      RECT MASK 2 77.474 46.569 83.764 46.709 ;
      RECT MASK 2 84.092 46.569 90.382 46.709 ;
      RECT MASK 2 90.71 46.569 97 46.709 ;
      RECT MASK 2 97.328 46.569 103.618 46.709 ;
      RECT MASK 2 103.946 46.569 110.236 46.709 ;
      RECT MASK 2 110.564 46.569 116.854 46.709 ;
      RECT MASK 2 117.182 46.569 127.884 46.709 ;
      RECT MASK 2 2.47 47.029 4.348 47.169 ;
      RECT MASK 2 4.676 47.029 10.966 47.169 ;
      RECT MASK 2 11.294 47.029 17.584 47.169 ;
      RECT MASK 2 17.912 47.029 24.202 47.169 ;
      RECT MASK 2 24.53 47.029 30.82 47.169 ;
      RECT MASK 2 31.148 47.029 37.438 47.169 ;
      RECT MASK 2 37.766 47.029 44.056 47.169 ;
      RECT MASK 2 44.384 47.029 50.674 47.169 ;
      RECT MASK 2 51.002 47.029 57.292 47.169 ;
      RECT MASK 2 57.62 47.029 63.91 47.169 ;
      RECT MASK 2 64.238 47.029 70.528 47.169 ;
      RECT MASK 2 70.856 47.029 77.146 47.169 ;
      RECT MASK 2 77.474 47.029 83.764 47.169 ;
      RECT MASK 2 84.092 47.029 90.382 47.169 ;
      RECT MASK 2 90.71 47.029 97 47.169 ;
      RECT MASK 2 97.328 47.029 103.618 47.169 ;
      RECT MASK 2 103.946 47.029 110.236 47.169 ;
      RECT MASK 2 110.564 47.029 116.854 47.169 ;
      RECT MASK 2 117.182 47.029 127.884 47.169 ;
      RECT MASK 2 2.47 47.919 4.348 48.059 ;
      RECT MASK 2 4.676 47.919 10.966 48.059 ;
      RECT MASK 2 11.294 47.919 17.584 48.059 ;
      RECT MASK 2 17.912 47.919 24.202 48.059 ;
      RECT MASK 2 24.53 47.919 30.82 48.059 ;
      RECT MASK 2 31.148 47.919 37.438 48.059 ;
      RECT MASK 2 37.766 47.919 44.056 48.059 ;
      RECT MASK 2 44.384 47.919 50.674 48.059 ;
      RECT MASK 2 51.002 47.919 57.292 48.059 ;
      RECT MASK 2 57.62 47.919 63.91 48.059 ;
      RECT MASK 2 64.238 47.919 70.528 48.059 ;
      RECT MASK 2 70.856 47.919 77.146 48.059 ;
      RECT MASK 2 77.474 47.919 83.764 48.059 ;
      RECT MASK 2 84.092 47.919 90.382 48.059 ;
      RECT MASK 2 90.71 47.919 97 48.059 ;
      RECT MASK 2 97.328 47.919 103.618 48.059 ;
      RECT MASK 2 103.946 47.919 110.236 48.059 ;
      RECT MASK 2 110.564 47.919 116.854 48.059 ;
      RECT MASK 2 117.182 47.919 127.884 48.059 ;
      RECT MASK 2 2.47 48.379 4.348 48.519 ;
      RECT MASK 2 4.676 48.379 10.966 48.519 ;
      RECT MASK 2 11.294 48.379 17.584 48.519 ;
      RECT MASK 2 17.912 48.379 24.202 48.519 ;
      RECT MASK 2 24.53 48.379 30.82 48.519 ;
      RECT MASK 2 31.148 48.379 37.438 48.519 ;
      RECT MASK 2 37.766 48.379 44.056 48.519 ;
      RECT MASK 2 44.384 48.379 50.674 48.519 ;
      RECT MASK 2 51.002 48.379 57.292 48.519 ;
      RECT MASK 2 57.62 48.379 63.91 48.519 ;
      RECT MASK 2 64.238 48.379 70.528 48.519 ;
      RECT MASK 2 70.856 48.379 77.146 48.519 ;
      RECT MASK 2 77.474 48.379 83.764 48.519 ;
      RECT MASK 2 84.092 48.379 90.382 48.519 ;
      RECT MASK 2 90.71 48.379 97 48.519 ;
      RECT MASK 2 97.328 48.379 103.618 48.519 ;
      RECT MASK 2 103.946 48.379 110.236 48.519 ;
      RECT MASK 2 110.564 48.379 116.854 48.519 ;
      RECT MASK 2 117.182 48.379 127.884 48.519 ;
      RECT MASK 2 2.47 49.269 4.348 49.409 ;
      RECT MASK 2 4.676 49.269 10.966 49.409 ;
      RECT MASK 2 11.294 49.269 17.584 49.409 ;
      RECT MASK 2 17.912 49.269 24.202 49.409 ;
      RECT MASK 2 24.53 49.269 30.82 49.409 ;
      RECT MASK 2 31.148 49.269 37.438 49.409 ;
      RECT MASK 2 37.766 49.269 44.056 49.409 ;
      RECT MASK 2 44.384 49.269 50.674 49.409 ;
      RECT MASK 2 51.002 49.269 57.292 49.409 ;
      RECT MASK 2 57.62 49.269 63.91 49.409 ;
      RECT MASK 2 64.238 49.269 70.528 49.409 ;
      RECT MASK 2 70.856 49.269 77.146 49.409 ;
      RECT MASK 2 77.474 49.269 83.764 49.409 ;
      RECT MASK 2 84.092 49.269 90.382 49.409 ;
      RECT MASK 2 90.71 49.269 97 49.409 ;
      RECT MASK 2 97.328 49.269 103.618 49.409 ;
      RECT MASK 2 103.946 49.269 110.236 49.409 ;
      RECT MASK 2 110.564 49.269 116.854 49.409 ;
      RECT MASK 2 117.182 49.269 123.472 49.409 ;
      RECT MASK 2 123.8 49.269 127.884 49.409 ;
      RECT MASK 2 2.47 49.729 4.348 49.869 ;
      RECT MASK 2 4.676 49.729 10.966 49.869 ;
      RECT MASK 2 11.294 49.729 17.584 49.869 ;
      RECT MASK 2 17.912 49.729 24.202 49.869 ;
      RECT MASK 2 24.53 49.729 30.82 49.869 ;
      RECT MASK 2 31.148 49.729 37.438 49.869 ;
      RECT MASK 2 37.766 49.729 44.056 49.869 ;
      RECT MASK 2 44.384 49.729 50.674 49.869 ;
      RECT MASK 2 51.002 49.729 57.292 49.869 ;
      RECT MASK 2 57.62 49.729 63.91 49.869 ;
      RECT MASK 2 64.238 49.729 70.528 49.869 ;
      RECT MASK 2 70.856 49.729 77.146 49.869 ;
      RECT MASK 2 77.474 49.729 83.764 49.869 ;
      RECT MASK 2 84.092 49.729 90.382 49.869 ;
      RECT MASK 2 90.71 49.729 97 49.869 ;
      RECT MASK 2 97.328 49.729 103.618 49.869 ;
      RECT MASK 2 103.946 49.729 110.236 49.869 ;
      RECT MASK 2 110.564 49.729 116.854 49.869 ;
      RECT MASK 2 117.182 49.729 123.472 49.869 ;
      RECT MASK 2 123.8 49.729 127.884 49.869 ;
      RECT MASK 2 2.47 50.619 4.348 50.759 ;
      RECT MASK 2 4.676 50.619 10.966 50.759 ;
      RECT MASK 2 11.294 50.619 17.584 50.759 ;
      RECT MASK 2 17.912 50.619 24.202 50.759 ;
      RECT MASK 2 24.53 50.619 30.82 50.759 ;
      RECT MASK 2 31.148 50.619 37.438 50.759 ;
      RECT MASK 2 37.766 50.619 44.056 50.759 ;
      RECT MASK 2 44.384 50.619 50.674 50.759 ;
      RECT MASK 2 51.002 50.619 57.292 50.759 ;
      RECT MASK 2 57.62 50.619 63.91 50.759 ;
      RECT MASK 2 64.238 50.619 70.528 50.759 ;
      RECT MASK 2 70.856 50.619 77.146 50.759 ;
      RECT MASK 2 77.474 50.619 83.764 50.759 ;
      RECT MASK 2 84.092 50.619 90.382 50.759 ;
      RECT MASK 2 90.71 50.619 97 50.759 ;
      RECT MASK 2 97.328 50.619 103.618 50.759 ;
      RECT MASK 2 103.946 50.619 110.236 50.759 ;
      RECT MASK 2 110.564 50.619 116.854 50.759 ;
      RECT MASK 2 117.182 50.619 123.472 50.759 ;
      RECT MASK 2 123.8 50.619 127.884 50.759 ;
      RECT MASK 2 110.564 51.059 123.472 51.239 ;
      RECT MASK 2 2.47 51.079 4.348 51.219 ;
      RECT MASK 2 4.676 51.079 10.966 51.219 ;
      RECT MASK 2 11.294 51.079 17.584 51.219 ;
      RECT MASK 2 17.912 51.079 24.202 51.219 ;
      RECT MASK 2 24.53 51.079 30.82 51.219 ;
      RECT MASK 2 31.148 51.079 37.438 51.219 ;
      RECT MASK 2 37.766 51.079 44.056 51.219 ;
      RECT MASK 2 44.384 51.079 50.674 51.219 ;
      RECT MASK 2 51.002 51.079 57.292 51.219 ;
      RECT MASK 2 57.62 51.079 63.91 51.219 ;
      RECT MASK 2 64.238 51.079 70.528 51.219 ;
      RECT MASK 2 70.856 51.079 77.146 51.219 ;
      RECT MASK 2 77.474 51.079 83.764 51.219 ;
      RECT MASK 2 84.092 51.079 90.382 51.219 ;
      RECT MASK 2 90.71 51.079 97 51.219 ;
      RECT MASK 2 97.328 51.079 103.618 51.219 ;
      RECT MASK 2 103.946 51.079 110.236 51.219 ;
      RECT MASK 2 123.8 51.079 127.884 51.219 ;
      RECT MASK 2 1.9425 51.62 41.8765 51.66 ;
      RECT MASK 2 42.6605 51.62 82.5945 51.66 ;
      RECT MASK 2 83.4005 51.62 128.3145 51.66 ;
      RECT MASK 2 1.9425 51.78 41.8765 51.82 ;
      RECT MASK 2 42.6605 51.78 82.5945 51.82 ;
      RECT MASK 2 83.4005 51.78 128.3145 51.82 ;
      RECT MASK 2 1.9425 52.04 41.8765 52.08 ;
      RECT MASK 2 42.6605 52.04 82.5945 52.08 ;
      RECT MASK 2 83.4005 52.04 128.3145 52.08 ;
      RECT MASK 2 1.9425 52.2 41.8765 52.24 ;
      RECT MASK 2 42.6605 52.2 82.5945 52.24 ;
      RECT MASK 2 83.4005 52.2 128.3145 52.24 ;
      RECT MASK 2 2.46 52.689 4.348 52.829 ;
      RECT MASK 2 4.676 52.689 10.966 52.829 ;
      RECT MASK 2 11.294 52.689 17.584 52.829 ;
      RECT MASK 2 17.912 52.689 24.202 52.829 ;
      RECT MASK 2 24.53 52.689 30.82 52.829 ;
      RECT MASK 2 31.148 52.689 37.438 52.829 ;
      RECT MASK 2 37.766 52.689 44.056 52.829 ;
      RECT MASK 2 44.384 52.689 50.674 52.829 ;
      RECT MASK 2 51.002 52.689 57.292 52.829 ;
      RECT MASK 2 57.62 52.689 63.91 52.829 ;
      RECT MASK 2 64.238 52.689 70.528 52.829 ;
      RECT MASK 2 70.856 52.689 77.146 52.829 ;
      RECT MASK 2 77.474 52.689 83.764 52.829 ;
      RECT MASK 2 84.092 52.689 90.382 52.829 ;
      RECT MASK 2 90.71 52.689 97 52.829 ;
      RECT MASK 2 97.328 52.689 103.618 52.829 ;
      RECT MASK 2 103.946 52.689 110.236 52.829 ;
      RECT MASK 2 110.564 52.689 123.472 52.829 ;
      RECT MASK 2 123.8 52.689 127.884 52.829 ;
      RECT MASK 2 2.46 53.149 4.348 53.289 ;
      RECT MASK 2 4.676 53.149 10.966 53.289 ;
      RECT MASK 2 11.294 53.149 17.584 53.289 ;
      RECT MASK 2 17.912 53.149 24.202 53.289 ;
      RECT MASK 2 24.53 53.149 30.82 53.289 ;
      RECT MASK 2 31.148 53.149 37.438 53.289 ;
      RECT MASK 2 37.766 53.149 44.056 53.289 ;
      RECT MASK 2 44.384 53.149 50.674 53.289 ;
      RECT MASK 2 51.002 53.149 57.292 53.289 ;
      RECT MASK 2 57.62 53.149 63.91 53.289 ;
      RECT MASK 2 64.238 53.149 70.528 53.289 ;
      RECT MASK 2 70.856 53.149 77.146 53.289 ;
      RECT MASK 2 77.474 53.149 83.764 53.289 ;
      RECT MASK 2 84.092 53.149 90.382 53.289 ;
      RECT MASK 2 90.71 53.149 97 53.289 ;
      RECT MASK 2 97.328 53.149 103.618 53.289 ;
      RECT MASK 2 103.946 53.149 110.236 53.289 ;
      RECT MASK 2 110.564 53.149 116.854 53.289 ;
      RECT MASK 2 117.182 53.149 123.472 53.289 ;
      RECT MASK 2 123.8 53.149 127.884 53.289 ;
      RECT MASK 2 2.46 54.039 4.348 54.179 ;
      RECT MASK 2 4.676 54.039 10.966 54.179 ;
      RECT MASK 2 11.294 54.039 17.584 54.179 ;
      RECT MASK 2 17.912 54.039 24.202 54.179 ;
      RECT MASK 2 24.53 54.039 30.82 54.179 ;
      RECT MASK 2 31.148 54.039 37.438 54.179 ;
      RECT MASK 2 37.766 54.039 44.056 54.179 ;
      RECT MASK 2 44.384 54.039 50.674 54.179 ;
      RECT MASK 2 51.002 54.039 57.292 54.179 ;
      RECT MASK 2 57.62 54.039 63.91 54.179 ;
      RECT MASK 2 64.238 54.039 70.528 54.179 ;
      RECT MASK 2 70.856 54.039 77.146 54.179 ;
      RECT MASK 2 77.474 54.039 83.764 54.179 ;
      RECT MASK 2 84.092 54.039 90.382 54.179 ;
      RECT MASK 2 90.71 54.039 97 54.179 ;
      RECT MASK 2 97.328 54.039 103.618 54.179 ;
      RECT MASK 2 103.946 54.039 110.236 54.179 ;
      RECT MASK 2 110.564 54.039 116.854 54.179 ;
      RECT MASK 2 117.182 54.039 123.472 54.179 ;
      RECT MASK 2 123.8 54.039 127.884 54.179 ;
      RECT MASK 2 2.46 54.499 4.348 54.639 ;
      RECT MASK 2 4.676 54.499 10.966 54.639 ;
      RECT MASK 2 11.294 54.499 17.584 54.639 ;
      RECT MASK 2 17.912 54.499 24.202 54.639 ;
      RECT MASK 2 24.53 54.499 30.82 54.639 ;
      RECT MASK 2 31.148 54.499 37.438 54.639 ;
      RECT MASK 2 37.766 54.499 44.056 54.639 ;
      RECT MASK 2 44.384 54.499 50.674 54.639 ;
      RECT MASK 2 51.002 54.499 57.292 54.639 ;
      RECT MASK 2 57.62 54.499 63.91 54.639 ;
      RECT MASK 2 64.238 54.499 70.528 54.639 ;
      RECT MASK 2 70.856 54.499 77.146 54.639 ;
      RECT MASK 2 77.474 54.499 83.764 54.639 ;
      RECT MASK 2 84.092 54.499 90.382 54.639 ;
      RECT MASK 2 90.71 54.499 97 54.639 ;
      RECT MASK 2 97.328 54.499 103.618 54.639 ;
      RECT MASK 2 103.946 54.499 110.236 54.639 ;
      RECT MASK 2 110.564 54.499 116.854 54.639 ;
      RECT MASK 2 117.182 54.499 123.472 54.639 ;
      RECT MASK 2 123.8 54.499 127.884 54.639 ;
      RECT MASK 2 2.46 55.389 4.348 55.529 ;
      RECT MASK 2 4.676 55.389 10.966 55.529 ;
      RECT MASK 2 11.294 55.389 17.584 55.529 ;
      RECT MASK 2 17.912 55.389 24.202 55.529 ;
      RECT MASK 2 24.53 55.389 30.82 55.529 ;
      RECT MASK 2 31.148 55.389 37.438 55.529 ;
      RECT MASK 2 37.766 55.389 44.056 55.529 ;
      RECT MASK 2 44.384 55.389 50.674 55.529 ;
      RECT MASK 2 51.002 55.389 57.292 55.529 ;
      RECT MASK 2 57.62 55.389 63.91 55.529 ;
      RECT MASK 2 64.238 55.389 70.528 55.529 ;
      RECT MASK 2 70.856 55.389 77.146 55.529 ;
      RECT MASK 2 77.474 55.389 83.764 55.529 ;
      RECT MASK 2 84.092 55.389 90.382 55.529 ;
      RECT MASK 2 90.71 55.389 97 55.529 ;
      RECT MASK 2 97.328 55.389 103.618 55.529 ;
      RECT MASK 2 103.946 55.389 110.236 55.529 ;
      RECT MASK 2 110.564 55.389 116.854 55.529 ;
      RECT MASK 2 117.182 55.389 127.884 55.529 ;
      RECT MASK 2 2.46 55.849 4.348 55.989 ;
      RECT MASK 2 4.676 55.849 10.966 55.989 ;
      RECT MASK 2 11.294 55.849 17.584 55.989 ;
      RECT MASK 2 17.912 55.849 24.202 55.989 ;
      RECT MASK 2 24.53 55.849 30.82 55.989 ;
      RECT MASK 2 31.148 55.849 37.438 55.989 ;
      RECT MASK 2 37.766 55.849 44.056 55.989 ;
      RECT MASK 2 44.384 55.849 50.674 55.989 ;
      RECT MASK 2 51.002 55.849 57.292 55.989 ;
      RECT MASK 2 57.62 55.849 63.91 55.989 ;
      RECT MASK 2 64.238 55.849 70.528 55.989 ;
      RECT MASK 2 70.856 55.849 77.146 55.989 ;
      RECT MASK 2 77.474 55.849 83.764 55.989 ;
      RECT MASK 2 84.092 55.849 90.382 55.989 ;
      RECT MASK 2 90.71 55.849 97 55.989 ;
      RECT MASK 2 97.328 55.849 103.618 55.989 ;
      RECT MASK 2 103.946 55.849 110.236 55.989 ;
      RECT MASK 2 110.564 55.849 116.854 55.989 ;
      RECT MASK 2 117.182 55.849 127.884 55.989 ;
      RECT MASK 2 2.46 56.739 4.348 56.879 ;
      RECT MASK 2 4.676 56.739 10.966 56.879 ;
      RECT MASK 2 11.294 56.739 17.584 56.879 ;
      RECT MASK 2 17.912 56.739 24.202 56.879 ;
      RECT MASK 2 24.53 56.739 30.82 56.879 ;
      RECT MASK 2 31.148 56.739 37.438 56.879 ;
      RECT MASK 2 37.766 56.739 44.056 56.879 ;
      RECT MASK 2 44.384 56.739 50.674 56.879 ;
      RECT MASK 2 51.002 56.739 57.292 56.879 ;
      RECT MASK 2 57.62 56.739 63.91 56.879 ;
      RECT MASK 2 64.238 56.739 70.528 56.879 ;
      RECT MASK 2 70.856 56.739 77.146 56.879 ;
      RECT MASK 2 77.474 56.739 83.764 56.879 ;
      RECT MASK 2 84.092 56.739 90.382 56.879 ;
      RECT MASK 2 90.71 56.739 97 56.879 ;
      RECT MASK 2 97.328 56.739 103.618 56.879 ;
      RECT MASK 2 103.946 56.739 110.236 56.879 ;
      RECT MASK 2 110.564 56.739 116.854 56.879 ;
      RECT MASK 2 117.182 56.739 127.884 56.879 ;
      RECT MASK 2 2.46 57.199 4.348 57.339 ;
      RECT MASK 2 4.676 57.199 10.966 57.339 ;
      RECT MASK 2 11.294 57.199 17.584 57.339 ;
      RECT MASK 2 17.912 57.199 24.202 57.339 ;
      RECT MASK 2 24.53 57.199 30.82 57.339 ;
      RECT MASK 2 31.148 57.199 37.438 57.339 ;
      RECT MASK 2 37.766 57.199 44.056 57.339 ;
      RECT MASK 2 44.384 57.199 50.674 57.339 ;
      RECT MASK 2 51.002 57.199 57.292 57.339 ;
      RECT MASK 2 57.62 57.199 63.91 57.339 ;
      RECT MASK 2 64.238 57.199 70.528 57.339 ;
      RECT MASK 2 70.856 57.199 77.146 57.339 ;
      RECT MASK 2 77.474 57.199 83.764 57.339 ;
      RECT MASK 2 84.092 57.199 90.382 57.339 ;
      RECT MASK 2 90.71 57.199 97 57.339 ;
      RECT MASK 2 97.328 57.199 103.618 57.339 ;
      RECT MASK 2 103.946 57.199 110.236 57.339 ;
      RECT MASK 2 110.564 57.199 116.854 57.339 ;
      RECT MASK 2 117.182 57.199 127.884 57.339 ;
      RECT MASK 2 1.9425 57.74 41.8765 57.78 ;
      RECT MASK 2 42.6605 57.74 82.5945 57.78 ;
      RECT MASK 2 83.4005 57.74 128.3145 57.78 ;
      RECT MASK 2 1.9425 57.9 41.8765 57.94 ;
      RECT MASK 2 42.6605 57.9 82.5945 57.94 ;
      RECT MASK 2 83.4005 57.9 128.3145 57.94 ;
      RECT MASK 2 1.9425 58.16 41.8765 58.2 ;
      RECT MASK 2 42.6605 58.16 82.5945 58.2 ;
      RECT MASK 2 83.4005 58.16 128.3145 58.2 ;
      RECT MASK 2 1.9425 58.32 41.8765 58.36 ;
      RECT MASK 2 42.6605 58.32 82.5945 58.36 ;
      RECT MASK 2 83.4005 58.32 128.3145 58.36 ;
      RECT MASK 2 2.46 58.809 4.348 58.949 ;
      RECT MASK 2 4.676 58.809 10.966 58.949 ;
      RECT MASK 2 11.294 58.809 17.584 58.949 ;
      RECT MASK 2 17.912 58.809 24.202 58.949 ;
      RECT MASK 2 24.53 58.809 30.82 58.949 ;
      RECT MASK 2 31.148 58.809 37.438 58.949 ;
      RECT MASK 2 37.766 58.809 44.056 58.949 ;
      RECT MASK 2 44.384 58.809 50.674 58.949 ;
      RECT MASK 2 51.002 58.809 57.292 58.949 ;
      RECT MASK 2 57.62 58.809 63.91 58.949 ;
      RECT MASK 2 64.238 58.809 70.528 58.949 ;
      RECT MASK 2 70.856 58.809 77.146 58.949 ;
      RECT MASK 2 77.474 58.809 83.764 58.949 ;
      RECT MASK 2 84.092 58.809 90.382 58.949 ;
      RECT MASK 2 90.71 58.809 97 58.949 ;
      RECT MASK 2 97.328 58.809 103.618 58.949 ;
      RECT MASK 2 103.946 58.809 110.236 58.949 ;
      RECT MASK 2 110.564 58.809 116.854 58.949 ;
      RECT MASK 2 117.182 58.809 127.884 58.949 ;
      RECT MASK 2 2.46 59.269 4.348 59.409 ;
      RECT MASK 2 4.676 59.269 10.966 59.409 ;
      RECT MASK 2 11.294 59.269 17.584 59.409 ;
      RECT MASK 2 17.912 59.269 24.202 59.409 ;
      RECT MASK 2 24.53 59.269 30.82 59.409 ;
      RECT MASK 2 31.148 59.269 37.438 59.409 ;
      RECT MASK 2 37.766 59.269 44.056 59.409 ;
      RECT MASK 2 44.384 59.269 50.674 59.409 ;
      RECT MASK 2 51.002 59.269 57.292 59.409 ;
      RECT MASK 2 57.62 59.269 63.91 59.409 ;
      RECT MASK 2 64.238 59.269 70.528 59.409 ;
      RECT MASK 2 70.856 59.269 77.146 59.409 ;
      RECT MASK 2 77.474 59.269 83.764 59.409 ;
      RECT MASK 2 84.092 59.269 90.382 59.409 ;
      RECT MASK 2 90.71 59.269 97 59.409 ;
      RECT MASK 2 97.328 59.269 103.618 59.409 ;
      RECT MASK 2 103.946 59.269 110.236 59.409 ;
      RECT MASK 2 110.564 59.269 116.854 59.409 ;
      RECT MASK 2 117.182 59.269 127.884 59.409 ;
      RECT MASK 2 2.46 60.159 4.348 60.299 ;
      RECT MASK 2 4.676 60.159 10.966 60.299 ;
      RECT MASK 2 11.294 60.159 17.584 60.299 ;
      RECT MASK 2 17.912 60.159 24.202 60.299 ;
      RECT MASK 2 24.53 60.159 30.82 60.299 ;
      RECT MASK 2 31.148 60.159 37.438 60.299 ;
      RECT MASK 2 37.766 60.159 44.056 60.299 ;
      RECT MASK 2 44.384 60.159 50.674 60.299 ;
      RECT MASK 2 51.002 60.159 57.292 60.299 ;
      RECT MASK 2 57.62 60.159 63.91 60.299 ;
      RECT MASK 2 64.238 60.159 70.528 60.299 ;
      RECT MASK 2 70.856 60.159 77.146 60.299 ;
      RECT MASK 2 77.474 60.159 83.764 60.299 ;
      RECT MASK 2 84.092 60.159 90.382 60.299 ;
      RECT MASK 2 90.71 60.159 97 60.299 ;
      RECT MASK 2 97.328 60.159 103.618 60.299 ;
      RECT MASK 2 103.946 60.159 110.236 60.299 ;
      RECT MASK 2 110.564 60.159 116.854 60.299 ;
      RECT MASK 2 117.182 60.159 127.884 60.299 ;
      RECT MASK 2 2.46 60.619 4.348 60.759 ;
      RECT MASK 2 4.676 60.619 10.966 60.759 ;
      RECT MASK 2 11.294 60.619 17.584 60.759 ;
      RECT MASK 2 17.912 60.619 24.202 60.759 ;
      RECT MASK 2 24.53 60.619 30.82 60.759 ;
      RECT MASK 2 31.148 60.619 37.438 60.759 ;
      RECT MASK 2 37.766 60.619 44.056 60.759 ;
      RECT MASK 2 44.384 60.619 50.674 60.759 ;
      RECT MASK 2 51.002 60.619 57.292 60.759 ;
      RECT MASK 2 57.62 60.619 63.91 60.759 ;
      RECT MASK 2 64.238 60.619 70.528 60.759 ;
      RECT MASK 2 70.856 60.619 77.146 60.759 ;
      RECT MASK 2 77.474 60.619 83.764 60.759 ;
      RECT MASK 2 84.092 60.619 90.382 60.759 ;
      RECT MASK 2 90.71 60.619 97 60.759 ;
      RECT MASK 2 97.328 60.619 103.618 60.759 ;
      RECT MASK 2 103.946 60.619 110.236 60.759 ;
      RECT MASK 2 110.564 60.619 116.854 60.759 ;
      RECT MASK 2 117.182 60.619 127.884 60.759 ;
      RECT MASK 2 2.46 61.509 4.348 61.649 ;
      RECT MASK 2 4.676 61.509 10.966 61.649 ;
      RECT MASK 2 11.294 61.509 17.584 61.649 ;
      RECT MASK 2 17.912 61.509 24.202 61.649 ;
      RECT MASK 2 24.53 61.509 30.82 61.649 ;
      RECT MASK 2 31.148 61.509 37.438 61.649 ;
      RECT MASK 2 37.766 61.509 44.056 61.649 ;
      RECT MASK 2 44.384 61.509 50.674 61.649 ;
      RECT MASK 2 51.002 61.509 57.292 61.649 ;
      RECT MASK 2 57.62 61.509 63.91 61.649 ;
      RECT MASK 2 64.238 61.509 70.528 61.649 ;
      RECT MASK 2 70.856 61.509 77.146 61.649 ;
      RECT MASK 2 77.474 61.509 83.764 61.649 ;
      RECT MASK 2 84.092 61.509 90.382 61.649 ;
      RECT MASK 2 90.71 61.509 97 61.649 ;
      RECT MASK 2 97.328 61.509 103.618 61.649 ;
      RECT MASK 2 103.946 61.509 110.236 61.649 ;
      RECT MASK 2 110.564 61.509 116.854 61.649 ;
      RECT MASK 2 117.182 61.509 127.884 61.649 ;
      RECT MASK 2 2.46 61.969 4.348 62.109 ;
      RECT MASK 2 4.676 61.969 10.966 62.109 ;
      RECT MASK 2 11.294 61.969 17.584 62.109 ;
      RECT MASK 2 17.912 61.969 24.202 62.109 ;
      RECT MASK 2 24.53 61.969 30.82 62.109 ;
      RECT MASK 2 31.148 61.969 37.438 62.109 ;
      RECT MASK 2 37.766 61.969 44.056 62.109 ;
      RECT MASK 2 44.384 61.969 50.674 62.109 ;
      RECT MASK 2 51.002 61.969 57.292 62.109 ;
      RECT MASK 2 57.62 61.969 63.91 62.109 ;
      RECT MASK 2 64.238 61.969 70.528 62.109 ;
      RECT MASK 2 70.856 61.969 77.146 62.109 ;
      RECT MASK 2 77.474 61.969 83.764 62.109 ;
      RECT MASK 2 84.092 61.969 90.382 62.109 ;
      RECT MASK 2 90.71 61.969 97 62.109 ;
      RECT MASK 2 97.328 61.969 103.618 62.109 ;
      RECT MASK 2 103.946 61.969 110.236 62.109 ;
      RECT MASK 2 110.564 61.969 116.854 62.109 ;
      RECT MASK 2 117.182 61.969 127.884 62.109 ;
      RECT MASK 2 2.46 62.859 4.348 62.999 ;
      RECT MASK 2 4.676 62.859 10.966 62.999 ;
      RECT MASK 2 11.294 62.859 17.584 62.999 ;
      RECT MASK 2 17.912 62.859 24.202 62.999 ;
      RECT MASK 2 24.53 62.859 30.82 62.999 ;
      RECT MASK 2 31.148 62.859 37.438 62.999 ;
      RECT MASK 2 37.766 62.859 44.056 62.999 ;
      RECT MASK 2 44.384 62.859 50.674 62.999 ;
      RECT MASK 2 51.002 62.859 57.292 62.999 ;
      RECT MASK 2 57.62 62.859 63.91 62.999 ;
      RECT MASK 2 64.238 62.859 70.528 62.999 ;
      RECT MASK 2 70.856 62.859 77.146 62.999 ;
      RECT MASK 2 77.474 62.859 83.764 62.999 ;
      RECT MASK 2 84.092 62.859 90.382 62.999 ;
      RECT MASK 2 90.71 62.859 97 62.999 ;
      RECT MASK 2 97.328 62.859 103.618 62.999 ;
      RECT MASK 2 103.946 62.859 110.236 62.999 ;
      RECT MASK 2 110.564 62.859 116.854 62.999 ;
      RECT MASK 2 117.182 62.859 127.884 62.999 ;
      RECT MASK 2 2.46 63.319 4.348 63.459 ;
      RECT MASK 2 4.676 63.319 10.966 63.459 ;
      RECT MASK 2 11.294 63.319 17.584 63.459 ;
      RECT MASK 2 17.912 63.319 24.202 63.459 ;
      RECT MASK 2 24.53 63.319 30.82 63.459 ;
      RECT MASK 2 31.148 63.319 37.438 63.459 ;
      RECT MASK 2 37.766 63.319 44.056 63.459 ;
      RECT MASK 2 44.384 63.319 50.674 63.459 ;
      RECT MASK 2 51.002 63.319 57.292 63.459 ;
      RECT MASK 2 57.62 63.319 63.91 63.459 ;
      RECT MASK 2 64.238 63.319 70.528 63.459 ;
      RECT MASK 2 70.856 63.319 77.146 63.459 ;
      RECT MASK 2 77.474 63.319 83.764 63.459 ;
      RECT MASK 2 84.092 63.319 90.382 63.459 ;
      RECT MASK 2 90.71 63.319 97 63.459 ;
      RECT MASK 2 97.328 63.319 103.618 63.459 ;
      RECT MASK 2 103.946 63.319 110.236 63.459 ;
      RECT MASK 2 110.564 63.319 116.854 63.459 ;
      RECT MASK 2 117.182 63.319 127.884 63.459 ;
      RECT MASK 2 1.9425 63.86 41.8765 63.9 ;
      RECT MASK 2 42.6605 63.86 82.5945 63.9 ;
      RECT MASK 2 83.4005 63.86 128.3145 63.9 ;
      RECT MASK 2 1.9425 64.02 41.8765 64.06 ;
      RECT MASK 2 42.6605 64.02 82.5945 64.06 ;
      RECT MASK 2 83.4005 64.02 128.3145 64.06 ;
      RECT MASK 2 1.9425 64.28 41.8765 64.32 ;
      RECT MASK 2 42.6605 64.28 82.5945 64.32 ;
      RECT MASK 2 83.4005 64.28 128.3145 64.32 ;
      RECT MASK 2 1.9425 64.44 41.8765 64.48 ;
      RECT MASK 2 42.6605 64.44 82.5945 64.48 ;
      RECT MASK 2 83.4005 64.44 128.3145 64.48 ;
      RECT MASK 2 2.46 64.929 4.348 65.069 ;
      RECT MASK 2 4.676 64.929 10.966 65.069 ;
      RECT MASK 2 11.294 64.929 17.584 65.069 ;
      RECT MASK 2 17.912 64.929 24.202 65.069 ;
      RECT MASK 2 24.53 64.929 30.82 65.069 ;
      RECT MASK 2 31.148 64.929 37.438 65.069 ;
      RECT MASK 2 37.766 64.929 44.056 65.069 ;
      RECT MASK 2 44.384 64.929 50.674 65.069 ;
      RECT MASK 2 51.002 64.929 57.292 65.069 ;
      RECT MASK 2 57.62 64.929 63.91 65.069 ;
      RECT MASK 2 64.238 64.929 70.528 65.069 ;
      RECT MASK 2 70.856 64.929 77.146 65.069 ;
      RECT MASK 2 77.474 64.929 83.764 65.069 ;
      RECT MASK 2 84.092 64.929 90.382 65.069 ;
      RECT MASK 2 90.71 64.929 97 65.069 ;
      RECT MASK 2 97.328 64.929 103.618 65.069 ;
      RECT MASK 2 103.946 64.929 110.236 65.069 ;
      RECT MASK 2 110.564 64.929 116.854 65.069 ;
      RECT MASK 2 117.182 64.929 127.884 65.069 ;
      RECT MASK 2 2.46 65.389 4.348 65.529 ;
      RECT MASK 2 4.676 65.389 10.966 65.529 ;
      RECT MASK 2 11.294 65.389 17.584 65.529 ;
      RECT MASK 2 17.912 65.389 24.202 65.529 ;
      RECT MASK 2 24.53 65.389 30.82 65.529 ;
      RECT MASK 2 31.148 65.389 37.438 65.529 ;
      RECT MASK 2 37.766 65.389 44.056 65.529 ;
      RECT MASK 2 44.384 65.389 50.674 65.529 ;
      RECT MASK 2 51.002 65.389 57.292 65.529 ;
      RECT MASK 2 57.62 65.389 63.91 65.529 ;
      RECT MASK 2 64.238 65.389 70.528 65.529 ;
      RECT MASK 2 70.856 65.389 77.146 65.529 ;
      RECT MASK 2 77.474 65.389 83.764 65.529 ;
      RECT MASK 2 84.092 65.389 90.382 65.529 ;
      RECT MASK 2 90.71 65.389 97 65.529 ;
      RECT MASK 2 97.328 65.389 103.618 65.529 ;
      RECT MASK 2 103.946 65.389 110.236 65.529 ;
      RECT MASK 2 110.564 65.389 116.854 65.529 ;
      RECT MASK 2 117.182 65.389 127.884 65.529 ;
      RECT MASK 2 2.46 66.279 4.348 66.419 ;
      RECT MASK 2 4.676 66.279 10.966 66.419 ;
      RECT MASK 2 11.294 66.279 17.584 66.419 ;
      RECT MASK 2 17.912 66.279 24.202 66.419 ;
      RECT MASK 2 24.53 66.279 30.82 66.419 ;
      RECT MASK 2 31.148 66.279 37.438 66.419 ;
      RECT MASK 2 37.766 66.279 44.056 66.419 ;
      RECT MASK 2 44.384 66.279 50.674 66.419 ;
      RECT MASK 2 51.002 66.279 57.292 66.419 ;
      RECT MASK 2 57.62 66.279 63.91 66.419 ;
      RECT MASK 2 64.238 66.279 70.528 66.419 ;
      RECT MASK 2 70.856 66.279 77.146 66.419 ;
      RECT MASK 2 77.474 66.279 83.764 66.419 ;
      RECT MASK 2 84.092 66.279 90.382 66.419 ;
      RECT MASK 2 90.71 66.279 97 66.419 ;
      RECT MASK 2 97.328 66.279 103.618 66.419 ;
      RECT MASK 2 103.946 66.279 110.236 66.419 ;
      RECT MASK 2 110.564 66.279 116.854 66.419 ;
      RECT MASK 2 117.182 66.279 127.884 66.419 ;
      RECT MASK 2 2.46 66.739 4.348 66.879 ;
      RECT MASK 2 4.676 66.739 10.966 66.879 ;
      RECT MASK 2 11.294 66.739 17.584 66.879 ;
      RECT MASK 2 17.912 66.739 24.202 66.879 ;
      RECT MASK 2 24.53 66.739 30.82 66.879 ;
      RECT MASK 2 31.148 66.739 37.438 66.879 ;
      RECT MASK 2 37.766 66.739 44.056 66.879 ;
      RECT MASK 2 44.384 66.739 50.674 66.879 ;
      RECT MASK 2 51.002 66.739 57.292 66.879 ;
      RECT MASK 2 57.62 66.739 63.91 66.879 ;
      RECT MASK 2 64.238 66.739 70.528 66.879 ;
      RECT MASK 2 70.856 66.739 77.146 66.879 ;
      RECT MASK 2 77.474 66.739 83.764 66.879 ;
      RECT MASK 2 84.092 66.739 90.382 66.879 ;
      RECT MASK 2 90.71 66.739 97 66.879 ;
      RECT MASK 2 97.328 66.739 103.618 66.879 ;
      RECT MASK 2 103.946 66.739 110.236 66.879 ;
      RECT MASK 2 110.564 66.739 116.854 66.879 ;
      RECT MASK 2 117.182 66.739 127.884 66.879 ;
      RECT MASK 2 2.46 67.629 4.348 67.769 ;
      RECT MASK 2 4.676 67.629 10.966 67.769 ;
      RECT MASK 2 11.294 67.629 17.584 67.769 ;
      RECT MASK 2 17.912 67.629 24.202 67.769 ;
      RECT MASK 2 24.53 67.629 30.82 67.769 ;
      RECT MASK 2 31.148 67.629 37.438 67.769 ;
      RECT MASK 2 37.766 67.629 44.056 67.769 ;
      RECT MASK 2 44.384 67.629 50.674 67.769 ;
      RECT MASK 2 51.002 67.629 57.292 67.769 ;
      RECT MASK 2 57.62 67.629 63.91 67.769 ;
      RECT MASK 2 64.238 67.629 70.528 67.769 ;
      RECT MASK 2 70.856 67.629 77.146 67.769 ;
      RECT MASK 2 77.474 67.629 83.764 67.769 ;
      RECT MASK 2 84.092 67.629 90.382 67.769 ;
      RECT MASK 2 90.71 67.629 97 67.769 ;
      RECT MASK 2 97.328 67.629 103.618 67.769 ;
      RECT MASK 2 103.946 67.629 110.236 67.769 ;
      RECT MASK 2 110.564 67.629 116.854 67.769 ;
      RECT MASK 2 117.182 67.629 127.884 67.769 ;
      RECT MASK 2 2.46 68.089 4.348 68.229 ;
      RECT MASK 2 4.676 68.089 10.966 68.229 ;
      RECT MASK 2 11.294 68.089 17.584 68.229 ;
      RECT MASK 2 17.912 68.089 24.202 68.229 ;
      RECT MASK 2 24.53 68.089 30.82 68.229 ;
      RECT MASK 2 31.148 68.089 37.438 68.229 ;
      RECT MASK 2 37.766 68.089 44.056 68.229 ;
      RECT MASK 2 44.384 68.089 50.674 68.229 ;
      RECT MASK 2 51.002 68.089 57.292 68.229 ;
      RECT MASK 2 57.62 68.089 63.91 68.229 ;
      RECT MASK 2 64.238 68.089 70.528 68.229 ;
      RECT MASK 2 70.856 68.089 77.146 68.229 ;
      RECT MASK 2 77.474 68.089 83.764 68.229 ;
      RECT MASK 2 84.092 68.089 90.382 68.229 ;
      RECT MASK 2 90.71 68.089 97 68.229 ;
      RECT MASK 2 97.328 68.089 103.618 68.229 ;
      RECT MASK 2 103.946 68.089 110.236 68.229 ;
      RECT MASK 2 110.564 68.089 116.854 68.229 ;
      RECT MASK 2 117.182 68.089 127.884 68.229 ;
      RECT MASK 2 2.46 68.979 4.348 69.119 ;
      RECT MASK 2 4.676 68.979 10.966 69.119 ;
      RECT MASK 2 11.294 68.979 17.584 69.119 ;
      RECT MASK 2 17.912 68.979 24.202 69.119 ;
      RECT MASK 2 24.53 68.979 30.82 69.119 ;
      RECT MASK 2 31.148 68.979 37.438 69.119 ;
      RECT MASK 2 37.766 68.979 44.056 69.119 ;
      RECT MASK 2 44.384 68.979 50.674 69.119 ;
      RECT MASK 2 51.002 68.979 57.292 69.119 ;
      RECT MASK 2 57.62 68.979 63.91 69.119 ;
      RECT MASK 2 64.238 68.979 70.528 69.119 ;
      RECT MASK 2 70.856 68.979 77.146 69.119 ;
      RECT MASK 2 77.474 68.979 83.764 69.119 ;
      RECT MASK 2 84.092 68.979 90.382 69.119 ;
      RECT MASK 2 90.71 68.979 97 69.119 ;
      RECT MASK 2 97.328 68.979 103.618 69.119 ;
      RECT MASK 2 103.946 68.979 110.236 69.119 ;
      RECT MASK 2 110.564 68.979 116.854 69.119 ;
      RECT MASK 2 117.182 68.979 127.884 69.119 ;
      RECT MASK 2 2.46 69.439 4.348 69.579 ;
      RECT MASK 2 4.676 69.439 10.966 69.579 ;
      RECT MASK 2 11.294 69.439 17.584 69.579 ;
      RECT MASK 2 17.912 69.439 24.202 69.579 ;
      RECT MASK 2 24.53 69.439 30.82 69.579 ;
      RECT MASK 2 31.148 69.439 37.438 69.579 ;
      RECT MASK 2 37.766 69.439 44.056 69.579 ;
      RECT MASK 2 44.384 69.439 50.674 69.579 ;
      RECT MASK 2 51.002 69.439 57.292 69.579 ;
      RECT MASK 2 57.62 69.439 63.91 69.579 ;
      RECT MASK 2 64.238 69.439 70.528 69.579 ;
      RECT MASK 2 70.856 69.439 77.146 69.579 ;
      RECT MASK 2 77.474 69.439 83.764 69.579 ;
      RECT MASK 2 84.092 69.439 90.382 69.579 ;
      RECT MASK 2 90.71 69.439 97 69.579 ;
      RECT MASK 2 97.328 69.439 103.618 69.579 ;
      RECT MASK 2 103.946 69.439 110.236 69.579 ;
      RECT MASK 2 110.564 69.439 116.854 69.579 ;
      RECT MASK 2 117.182 69.439 127.884 69.579 ;
      RECT MASK 2 1.9425 69.98 41.8765 70.02 ;
      RECT MASK 2 42.6605 69.98 82.5945 70.02 ;
      RECT MASK 2 83.4005 69.98 128.3145 70.02 ;
      RECT MASK 2 1.9425 70.14 41.8765 70.18 ;
      RECT MASK 2 42.6605 70.14 82.5945 70.18 ;
      RECT MASK 2 83.4005 70.14 128.3145 70.18 ;
      RECT MASK 2 1.9425 70.4 41.8765 70.44 ;
      RECT MASK 2 42.6605 70.4 82.5945 70.44 ;
      RECT MASK 2 83.4005 70.4 128.3145 70.44 ;
      RECT MASK 2 1.9425 70.56 41.8765 70.6 ;
      RECT MASK 2 42.6605 70.56 82.5945 70.6 ;
      RECT MASK 2 83.4005 70.56 128.3145 70.6 ;
      RECT MASK 2 2.46 71.049 4.348 71.189 ;
      RECT MASK 2 4.676 71.049 10.966 71.189 ;
      RECT MASK 2 11.294 71.049 17.584 71.189 ;
      RECT MASK 2 17.912 71.049 24.202 71.189 ;
      RECT MASK 2 24.53 71.049 30.82 71.189 ;
      RECT MASK 2 31.148 71.049 37.438 71.189 ;
      RECT MASK 2 37.766 71.049 44.056 71.189 ;
      RECT MASK 2 44.384 71.049 50.674 71.189 ;
      RECT MASK 2 51.002 71.049 57.292 71.189 ;
      RECT MASK 2 57.62 71.049 63.91 71.189 ;
      RECT MASK 2 64.238 71.049 70.528 71.189 ;
      RECT MASK 2 70.856 71.049 77.146 71.189 ;
      RECT MASK 2 77.474 71.049 83.764 71.189 ;
      RECT MASK 2 84.092 71.049 90.382 71.189 ;
      RECT MASK 2 90.71 71.049 97 71.189 ;
      RECT MASK 2 97.328 71.049 103.618 71.189 ;
      RECT MASK 2 103.946 71.049 110.236 71.189 ;
      RECT MASK 2 110.564 71.049 116.854 71.189 ;
      RECT MASK 2 117.182 71.049 127.884 71.189 ;
      RECT MASK 2 2.46 71.509 4.348 71.649 ;
      RECT MASK 2 4.676 71.509 10.966 71.649 ;
      RECT MASK 2 11.294 71.509 17.584 71.649 ;
      RECT MASK 2 17.912 71.509 24.202 71.649 ;
      RECT MASK 2 24.53 71.509 30.82 71.649 ;
      RECT MASK 2 31.148 71.509 37.438 71.649 ;
      RECT MASK 2 37.766 71.509 44.056 71.649 ;
      RECT MASK 2 44.384 71.509 50.674 71.649 ;
      RECT MASK 2 51.002 71.509 57.292 71.649 ;
      RECT MASK 2 57.62 71.509 63.91 71.649 ;
      RECT MASK 2 64.238 71.509 70.528 71.649 ;
      RECT MASK 2 70.856 71.509 77.146 71.649 ;
      RECT MASK 2 77.474 71.509 83.764 71.649 ;
      RECT MASK 2 84.092 71.509 90.382 71.649 ;
      RECT MASK 2 90.71 71.509 97 71.649 ;
      RECT MASK 2 97.328 71.509 103.618 71.649 ;
      RECT MASK 2 103.946 71.509 110.236 71.649 ;
      RECT MASK 2 110.564 71.509 116.854 71.649 ;
      RECT MASK 2 117.182 71.509 127.884 71.649 ;
      RECT MASK 2 113.869 72.29 129.095 72.33 ;
      RECT MASK 2 2.46 72.399 4.348 72.539 ;
      RECT MASK 2 4.676 72.399 10.966 72.539 ;
      RECT MASK 2 11.294 72.399 17.584 72.539 ;
      RECT MASK 2 17.912 72.399 24.202 72.539 ;
      RECT MASK 2 24.53 72.399 30.82 72.539 ;
      RECT MASK 2 31.148 72.399 37.438 72.539 ;
      RECT MASK 2 37.766 72.399 44.056 72.539 ;
      RECT MASK 2 44.384 72.399 50.674 72.539 ;
      RECT MASK 2 51.002 72.399 57.292 72.539 ;
      RECT MASK 2 57.62 72.399 63.91 72.539 ;
      RECT MASK 2 64.238 72.399 70.528 72.539 ;
      RECT MASK 2 70.856 72.399 77.146 72.539 ;
      RECT MASK 2 77.474 72.399 83.764 72.539 ;
      RECT MASK 2 84.092 72.399 90.382 72.539 ;
      RECT MASK 2 90.71 72.399 97 72.539 ;
      RECT MASK 2 97.328 72.399 103.618 72.539 ;
      RECT MASK 2 103.946 72.399 110.236 72.539 ;
      RECT MASK 2 110.564 72.399 112.463 72.539 ;
      RECT MASK 2 113.869 72.48 129.095 72.52 ;
      RECT MASK 2 114.345 72.77 129.322 72.81 ;
      RECT MASK 2 2.46 72.859 4.348 72.999 ;
      RECT MASK 2 4.676 72.859 10.966 72.999 ;
      RECT MASK 2 11.294 72.859 17.584 72.999 ;
      RECT MASK 2 17.912 72.859 24.202 72.999 ;
      RECT MASK 2 24.53 72.859 30.82 72.999 ;
      RECT MASK 2 31.148 72.859 37.438 72.999 ;
      RECT MASK 2 37.766 72.859 44.056 72.999 ;
      RECT MASK 2 44.384 72.859 50.674 72.999 ;
      RECT MASK 2 51.002 72.859 57.292 72.999 ;
      RECT MASK 2 57.62 72.859 63.91 72.999 ;
      RECT MASK 2 64.238 72.859 70.528 72.999 ;
      RECT MASK 2 70.856 72.859 77.146 72.999 ;
      RECT MASK 2 77.474 72.859 83.764 72.999 ;
      RECT MASK 2 84.092 72.859 90.382 72.999 ;
      RECT MASK 2 90.71 72.859 97 72.999 ;
      RECT MASK 2 97.328 72.859 103.618 72.999 ;
      RECT MASK 2 103.946 72.859 110.236 72.999 ;
      RECT MASK 2 110.564 72.859 112.463 72.999 ;
      RECT MASK 2 114.345 72.96 129.322 73 ;
      RECT MASK 2 115.539 73.25 126.947 73.29 ;
      RECT MASK 2 115.539 73.44 126.947 73.48 ;
      RECT MASK 2 2.46 73.749 4.348 73.889 ;
      RECT MASK 2 4.676 73.749 10.966 73.889 ;
      RECT MASK 2 11.294 73.749 17.584 73.889 ;
      RECT MASK 2 17.912 73.749 24.202 73.889 ;
      RECT MASK 2 24.53 73.749 30.82 73.889 ;
      RECT MASK 2 31.148 73.749 37.438 73.889 ;
      RECT MASK 2 37.766 73.749 44.056 73.889 ;
      RECT MASK 2 44.384 73.749 50.674 73.889 ;
      RECT MASK 2 51.002 73.749 57.292 73.889 ;
      RECT MASK 2 57.62 73.749 63.91 73.889 ;
      RECT MASK 2 64.238 73.749 70.528 73.889 ;
      RECT MASK 2 70.856 73.749 77.146 73.889 ;
      RECT MASK 2 77.474 73.749 83.764 73.889 ;
      RECT MASK 2 84.092 73.749 90.382 73.889 ;
      RECT MASK 2 90.71 73.749 97 73.889 ;
      RECT MASK 2 97.328 73.749 103.618 73.889 ;
      RECT MASK 2 103.946 73.749 110.236 73.889 ;
      RECT MASK 2 110.564 73.749 112.463 73.889 ;
      RECT MASK 2 116.437 73.988 116.497 74.212 ;
      RECT MASK 2 116.769 73.988 116.829 74.212 ;
      RECT MASK 2 117.101 73.988 117.161 74.212 ;
      RECT MASK 2 117.433 73.988 117.493 74.212 ;
      RECT MASK 2 117.765 73.988 117.825 74.212 ;
      RECT MASK 2 118.097 73.988 118.157 74.212 ;
      RECT MASK 2 118.429 73.988 118.489 74.212 ;
      RECT MASK 2 118.761 73.988 118.821 74.212 ;
      RECT MASK 2 119.093 73.988 119.153 74.212 ;
      RECT MASK 2 119.425 73.988 119.485 74.212 ;
      RECT MASK 2 119.757 73.988 119.817 74.212 ;
      RECT MASK 2 120.089 73.988 120.149 74.212 ;
      RECT MASK 2 120.421 73.988 120.481 74.212 ;
      RECT MASK 2 120.753 73.988 120.813 74.212 ;
      RECT MASK 2 121.085 73.988 121.145 74.212 ;
      RECT MASK 2 121.417 73.988 121.477 74.212 ;
      RECT MASK 2 121.749 73.988 121.809 74.212 ;
      RECT MASK 2 122.081 73.988 122.141 74.212 ;
      RECT MASK 2 122.413 73.988 122.473 74.212 ;
      RECT MASK 2 122.745 73.988 122.805 74.212 ;
      RECT MASK 2 123.077 73.988 123.137 74.212 ;
      RECT MASK 2 123.409 73.988 123.469 74.212 ;
      RECT MASK 2 123.741 73.988 123.801 74.212 ;
      RECT MASK 2 124.073 73.988 124.133 74.212 ;
      RECT MASK 2 124.405 73.988 124.465 74.212 ;
      RECT MASK 2 124.737 73.988 124.797 74.212 ;
      RECT MASK 2 125.069 73.988 125.129 74.212 ;
      RECT MASK 2 125.401 73.988 125.461 74.212 ;
      RECT MASK 2 125.733 73.988 125.793 74.212 ;
      RECT MASK 2 126.065 73.988 126.125 74.212 ;
      RECT MASK 2 2.46 74.209 4.348 74.349 ;
      RECT MASK 2 4.676 74.209 10.966 74.349 ;
      RECT MASK 2 11.294 74.209 17.584 74.349 ;
      RECT MASK 2 17.912 74.209 24.202 74.349 ;
      RECT MASK 2 24.53 74.209 30.82 74.349 ;
      RECT MASK 2 31.148 74.209 37.438 74.349 ;
      RECT MASK 2 37.766 74.209 44.056 74.349 ;
      RECT MASK 2 44.384 74.209 50.674 74.349 ;
      RECT MASK 2 51.002 74.209 57.292 74.349 ;
      RECT MASK 2 57.62 74.209 63.91 74.349 ;
      RECT MASK 2 64.238 74.209 70.528 74.349 ;
      RECT MASK 2 70.856 74.209 77.146 74.349 ;
      RECT MASK 2 77.474 74.209 83.764 74.349 ;
      RECT MASK 2 84.092 74.209 90.382 74.349 ;
      RECT MASK 2 90.71 74.209 97 74.349 ;
      RECT MASK 2 97.328 74.209 103.618 74.349 ;
      RECT MASK 2 103.946 74.209 110.236 74.349 ;
      RECT MASK 2 110.564 74.209 112.463 74.349 ;
      RECT MASK 2 116.079 74.4325 116.2725 74.4725 ;
      RECT MASK 2 126.2895 74.4325 126.483 74.4725 ;
      RECT MASK 2 116.437 74.768 116.497 74.992 ;
      RECT MASK 2 116.769 74.768 116.829 74.992 ;
      RECT MASK 2 117.101 74.768 117.161 74.992 ;
      RECT MASK 2 117.433 74.768 117.493 74.992 ;
      RECT MASK 2 117.765 74.768 117.825 74.992 ;
      RECT MASK 2 118.097 74.768 118.157 74.992 ;
      RECT MASK 2 118.429 74.768 118.489 74.992 ;
      RECT MASK 2 118.761 74.768 118.821 74.992 ;
      RECT MASK 2 119.093 74.768 119.153 74.992 ;
      RECT MASK 2 119.425 74.768 119.485 74.992 ;
      RECT MASK 2 119.757 74.768 119.817 74.992 ;
      RECT MASK 2 120.089 74.768 120.149 74.992 ;
      RECT MASK 2 120.421 74.768 120.481 74.992 ;
      RECT MASK 2 120.753 74.768 120.813 74.992 ;
      RECT MASK 2 121.085 74.768 121.145 74.992 ;
      RECT MASK 2 121.417 74.768 121.477 74.992 ;
      RECT MASK 2 121.749 74.768 121.809 74.992 ;
      RECT MASK 2 122.081 74.768 122.141 74.992 ;
      RECT MASK 2 122.413 74.768 122.473 74.992 ;
      RECT MASK 2 122.745 74.768 122.805 74.992 ;
      RECT MASK 2 123.077 74.768 123.137 74.992 ;
      RECT MASK 2 123.409 74.768 123.469 74.992 ;
      RECT MASK 2 123.741 74.768 123.801 74.992 ;
      RECT MASK 2 124.073 74.768 124.133 74.992 ;
      RECT MASK 2 124.405 74.768 124.465 74.992 ;
      RECT MASK 2 124.737 74.768 124.797 74.992 ;
      RECT MASK 2 125.069 74.768 125.129 74.992 ;
      RECT MASK 2 125.401 74.768 125.461 74.992 ;
      RECT MASK 2 125.733 74.768 125.793 74.992 ;
      RECT MASK 2 126.065 74.768 126.125 74.992 ;
      RECT MASK 2 2.46 75.099 4.348 75.239 ;
      RECT MASK 2 4.676 75.099 10.966 75.239 ;
      RECT MASK 2 11.294 75.099 17.584 75.239 ;
      RECT MASK 2 17.912 75.099 24.202 75.239 ;
      RECT MASK 2 24.53 75.099 30.82 75.239 ;
      RECT MASK 2 31.148 75.099 37.438 75.239 ;
      RECT MASK 2 37.766 75.099 44.056 75.239 ;
      RECT MASK 2 44.384 75.099 50.674 75.239 ;
      RECT MASK 2 51.002 75.099 57.292 75.239 ;
      RECT MASK 2 57.62 75.099 63.91 75.239 ;
      RECT MASK 2 64.238 75.099 70.528 75.239 ;
      RECT MASK 2 70.856 75.099 77.146 75.239 ;
      RECT MASK 2 77.474 75.099 83.764 75.239 ;
      RECT MASK 2 84.092 75.099 90.382 75.239 ;
      RECT MASK 2 90.71 75.099 97 75.239 ;
      RECT MASK 2 97.328 75.099 103.618 75.239 ;
      RECT MASK 2 103.946 75.099 110.236 75.239 ;
      RECT MASK 2 110.564 75.099 112.463 75.239 ;
      RECT MASK 2 116.079 75.2125 116.2725 75.2525 ;
      RECT MASK 2 126.2895 75.2125 126.483 75.2525 ;
      RECT MASK 2 116.437 75.548 116.497 75.772 ;
      RECT MASK 2 116.769 75.548 116.829 75.772 ;
      RECT MASK 2 117.101 75.548 117.161 75.772 ;
      RECT MASK 2 117.433 75.548 117.493 75.772 ;
      RECT MASK 2 117.765 75.548 117.825 75.772 ;
      RECT MASK 2 118.097 75.548 118.157 75.772 ;
      RECT MASK 2 118.429 75.548 118.489 75.772 ;
      RECT MASK 2 118.761 75.548 118.821 75.772 ;
      RECT MASK 2 119.093 75.548 119.153 75.772 ;
      RECT MASK 2 119.425 75.548 119.485 75.772 ;
      RECT MASK 2 119.757 75.548 119.817 75.772 ;
      RECT MASK 2 120.089 75.548 120.149 75.772 ;
      RECT MASK 2 120.421 75.548 120.481 75.772 ;
      RECT MASK 2 120.753 75.548 120.813 75.772 ;
      RECT MASK 2 121.085 75.548 121.145 75.772 ;
      RECT MASK 2 121.417 75.548 121.477 75.772 ;
      RECT MASK 2 121.749 75.548 121.809 75.772 ;
      RECT MASK 2 122.081 75.548 122.141 75.772 ;
      RECT MASK 2 122.413 75.548 122.473 75.772 ;
      RECT MASK 2 122.745 75.548 122.805 75.772 ;
      RECT MASK 2 123.077 75.548 123.137 75.772 ;
      RECT MASK 2 123.409 75.548 123.469 75.772 ;
      RECT MASK 2 123.741 75.548 123.801 75.772 ;
      RECT MASK 2 124.073 75.548 124.133 75.772 ;
      RECT MASK 2 124.405 75.548 124.465 75.772 ;
      RECT MASK 2 124.737 75.548 124.797 75.772 ;
      RECT MASK 2 125.069 75.548 125.129 75.772 ;
      RECT MASK 2 125.401 75.548 125.461 75.772 ;
      RECT MASK 2 125.733 75.548 125.793 75.772 ;
      RECT MASK 2 126.065 75.548 126.125 75.772 ;
      RECT MASK 2 2.46 75.559 4.348 75.699 ;
      RECT MASK 2 4.676 75.559 10.966 75.699 ;
      RECT MASK 2 11.294 75.559 17.584 75.699 ;
      RECT MASK 2 17.912 75.559 24.202 75.699 ;
      RECT MASK 2 24.53 75.559 30.82 75.699 ;
      RECT MASK 2 31.148 75.559 37.438 75.699 ;
      RECT MASK 2 37.766 75.559 44.056 75.699 ;
      RECT MASK 2 44.384 75.559 50.674 75.699 ;
      RECT MASK 2 51.002 75.559 57.292 75.699 ;
      RECT MASK 2 57.62 75.559 63.91 75.699 ;
      RECT MASK 2 64.238 75.559 70.528 75.699 ;
      RECT MASK 2 70.856 75.559 77.146 75.699 ;
      RECT MASK 2 77.474 75.559 83.764 75.699 ;
      RECT MASK 2 84.092 75.559 90.382 75.699 ;
      RECT MASK 2 90.71 75.559 97 75.699 ;
      RECT MASK 2 97.328 75.559 103.618 75.699 ;
      RECT MASK 2 103.946 75.559 110.236 75.699 ;
      RECT MASK 2 110.564 75.559 112.463 75.699 ;
      RECT MASK 2 116.079 75.9925 116.2725 76.0325 ;
      RECT MASK 2 126.2895 75.9925 126.483 76.0325 ;
      RECT MASK 2 116.437 76.328 116.497 76.552 ;
      RECT MASK 2 116.769 76.328 116.829 76.552 ;
      RECT MASK 2 117.101 76.328 117.161 76.552 ;
      RECT MASK 2 117.433 76.328 117.493 76.552 ;
      RECT MASK 2 117.765 76.328 117.825 76.552 ;
      RECT MASK 2 118.097 76.328 118.157 76.552 ;
      RECT MASK 2 118.429 76.328 118.489 76.552 ;
      RECT MASK 2 118.761 76.328 118.821 76.552 ;
      RECT MASK 2 119.093 76.328 119.153 76.552 ;
      RECT MASK 2 119.425 76.328 119.485 76.552 ;
      RECT MASK 2 119.757 76.328 119.817 76.552 ;
      RECT MASK 2 120.089 76.328 120.149 76.552 ;
      RECT MASK 2 120.421 76.328 120.481 76.552 ;
      RECT MASK 2 120.753 76.328 120.813 76.552 ;
      RECT MASK 2 121.085 76.328 121.145 76.552 ;
      RECT MASK 2 121.417 76.328 121.477 76.552 ;
      RECT MASK 2 121.749 76.328 121.809 76.552 ;
      RECT MASK 2 122.081 76.328 122.141 76.552 ;
      RECT MASK 2 122.413 76.328 122.473 76.552 ;
      RECT MASK 2 122.745 76.328 122.805 76.552 ;
      RECT MASK 2 123.077 76.328 123.137 76.552 ;
      RECT MASK 2 123.409 76.328 123.469 76.552 ;
      RECT MASK 2 123.741 76.328 123.801 76.552 ;
      RECT MASK 2 124.073 76.328 124.133 76.552 ;
      RECT MASK 2 124.405 76.328 124.465 76.552 ;
      RECT MASK 2 124.737 76.328 124.797 76.552 ;
      RECT MASK 2 125.069 76.328 125.129 76.552 ;
      RECT MASK 2 125.401 76.328 125.461 76.552 ;
      RECT MASK 2 125.733 76.328 125.793 76.552 ;
      RECT MASK 2 126.065 76.328 126.125 76.552 ;
      RECT MASK 2 2.47 76.449 112.442 76.589 ;
      RECT MASK 2 116.079 76.7725 116.2725 76.8125 ;
      RECT MASK 2 126.2895 76.7725 126.483 76.8125 ;
      RECT MASK 2 2.47 76.909 112.442 77.049 ;
      RECT MASK 2 116.437 77.108 116.497 77.332 ;
      RECT MASK 2 116.769 77.108 116.829 77.332 ;
      RECT MASK 2 117.101 77.108 117.161 77.332 ;
      RECT MASK 2 117.433 77.108 117.493 77.332 ;
      RECT MASK 2 117.765 77.108 117.825 77.332 ;
      RECT MASK 2 118.097 77.108 118.157 77.332 ;
      RECT MASK 2 118.429 77.108 118.489 77.332 ;
      RECT MASK 2 118.761 77.108 118.821 77.332 ;
      RECT MASK 2 119.093 77.108 119.153 77.332 ;
      RECT MASK 2 119.425 77.108 119.485 77.332 ;
      RECT MASK 2 119.757 77.108 119.817 77.332 ;
      RECT MASK 2 120.089 77.108 120.149 77.332 ;
      RECT MASK 2 120.421 77.108 120.481 77.332 ;
      RECT MASK 2 120.753 77.108 120.813 77.332 ;
      RECT MASK 2 121.085 77.108 121.145 77.332 ;
      RECT MASK 2 121.417 77.108 121.477 77.332 ;
      RECT MASK 2 121.749 77.108 121.809 77.332 ;
      RECT MASK 2 122.081 77.108 122.141 77.332 ;
      RECT MASK 2 122.413 77.108 122.473 77.332 ;
      RECT MASK 2 122.745 77.108 122.805 77.332 ;
      RECT MASK 2 123.077 77.108 123.137 77.332 ;
      RECT MASK 2 123.409 77.108 123.469 77.332 ;
      RECT MASK 2 123.741 77.108 123.801 77.332 ;
      RECT MASK 2 124.073 77.108 124.133 77.332 ;
      RECT MASK 2 124.405 77.108 124.465 77.332 ;
      RECT MASK 2 124.737 77.108 124.797 77.332 ;
      RECT MASK 2 125.069 77.108 125.129 77.332 ;
      RECT MASK 2 125.401 77.108 125.461 77.332 ;
      RECT MASK 2 125.733 77.108 125.793 77.332 ;
      RECT MASK 2 126.065 77.108 126.125 77.332 ;
      RECT MASK 2 1.31 77.54 113.984 77.58 ;
      RECT MASK 2 116.079 77.5525 116.2725 77.5925 ;
      RECT MASK 2 126.2895 77.5525 126.483 77.5925 ;
      RECT MASK 2 1.31 77.73 113.984 77.77 ;
      RECT MASK 2 116.437 77.888 116.497 78.112 ;
      RECT MASK 2 116.769 77.888 116.829 78.112 ;
      RECT MASK 2 117.101 77.888 117.161 78.112 ;
      RECT MASK 2 117.433 77.888 117.493 78.112 ;
      RECT MASK 2 117.765 77.888 117.825 78.112 ;
      RECT MASK 2 118.097 77.888 118.157 78.112 ;
      RECT MASK 2 118.429 77.888 118.489 78.112 ;
      RECT MASK 2 118.761 77.888 118.821 78.112 ;
      RECT MASK 2 119.093 77.888 119.153 78.112 ;
      RECT MASK 2 119.425 77.888 119.485 78.112 ;
      RECT MASK 2 119.757 77.888 119.817 78.112 ;
      RECT MASK 2 120.089 77.888 120.149 78.112 ;
      RECT MASK 2 120.421 77.888 120.481 78.112 ;
      RECT MASK 2 120.753 77.888 120.813 78.112 ;
      RECT MASK 2 121.085 77.888 121.145 78.112 ;
      RECT MASK 2 121.417 77.888 121.477 78.112 ;
      RECT MASK 2 121.749 77.888 121.809 78.112 ;
      RECT MASK 2 122.081 77.888 122.141 78.112 ;
      RECT MASK 2 122.413 77.888 122.473 78.112 ;
      RECT MASK 2 122.745 77.888 122.805 78.112 ;
      RECT MASK 2 123.077 77.888 123.137 78.112 ;
      RECT MASK 2 123.409 77.888 123.469 78.112 ;
      RECT MASK 2 123.741 77.888 123.801 78.112 ;
      RECT MASK 2 124.073 77.888 124.133 78.112 ;
      RECT MASK 2 124.405 77.888 124.465 78.112 ;
      RECT MASK 2 124.737 77.888 124.797 78.112 ;
      RECT MASK 2 125.069 77.888 125.129 78.112 ;
      RECT MASK 2 125.401 77.888 125.461 78.112 ;
      RECT MASK 2 125.733 77.888 125.793 78.112 ;
      RECT MASK 2 126.065 77.888 126.125 78.112 ;
      RECT MASK 2 6.224 78.05 110.065 78.09 ;
      RECT MASK 2 6.224 78.24 110.065 78.28 ;
      RECT MASK 2 116.079 78.3325 116.2725 78.3725 ;
      RECT MASK 2 126.2895 78.3325 126.483 78.3725 ;
      RECT MASK 2 11.941 78.4895 12.021 79.4645 ;
      RECT MASK 2 16.921 78.4895 17.001 79.4645 ;
      RECT MASK 2 18.559 78.4895 18.639 79.4645 ;
      RECT MASK 2 23.539 78.4895 23.619 79.4645 ;
      RECT MASK 2 25.177 78.4895 25.257 79.4645 ;
      RECT MASK 2 30.157 78.4895 30.237 79.4645 ;
      RECT MASK 2 31.795 78.4895 31.875 79.4645 ;
      RECT MASK 2 36.775 78.4895 36.855 79.4645 ;
      RECT MASK 2 38.413 78.4895 38.493 79.4645 ;
      RECT MASK 2 43.393 78.4895 43.473 79.4645 ;
      RECT MASK 2 45.031 78.4895 45.111 79.4645 ;
      RECT MASK 2 50.011 78.4895 50.091 79.4645 ;
      RECT MASK 2 51.649 78.4895 51.729 79.4645 ;
      RECT MASK 2 56.629 78.4895 56.709 79.4645 ;
      RECT MASK 2 58.267 78.4895 58.347 79.4645 ;
      RECT MASK 2 63.247 78.4895 63.327 79.4645 ;
      RECT MASK 2 64.885 78.4895 64.965 79.4645 ;
      RECT MASK 2 69.865 78.4895 69.945 79.4645 ;
      RECT MASK 2 71.503 78.4895 71.583 79.4645 ;
      RECT MASK 2 76.483 78.4895 76.563 79.4645 ;
      RECT MASK 2 78.121 78.4895 78.201 79.4645 ;
      RECT MASK 2 83.101 78.4895 83.181 79.4645 ;
      RECT MASK 2 84.739 78.4895 84.819 79.4645 ;
      RECT MASK 2 89.719 78.4895 89.799 79.4645 ;
      RECT MASK 2 91.357 78.4895 91.437 79.4645 ;
      RECT MASK 2 96.337 78.4895 96.417 79.4645 ;
      RECT MASK 2 97.975 78.4895 98.055 79.4645 ;
      RECT MASK 2 102.955 78.4895 103.035 79.4645 ;
      RECT MASK 2 104.593 78.4895 104.673 79.4645 ;
      RECT MASK 2 109.573 78.4895 109.653 79.4645 ;
      RECT MASK 2 1.248 78.56 5.362 78.6 ;
      RECT MASK 2 6.817 78.586 6.897 78.813 ;
      RECT MASK 2 7.149 78.586 7.229 78.813 ;
      RECT MASK 2 7.481 78.586 7.561 78.813 ;
      RECT MASK 2 7.979 78.586 8.059 78.813 ;
      RECT MASK 2 8.311 78.586 8.391 78.813 ;
      RECT MASK 2 8.643 78.586 8.723 78.813 ;
      RECT MASK 2 9.141 78.586 9.221 78.813 ;
      RECT MASK 2 9.473 78.586 9.553 78.813 ;
      RECT MASK 2 9.805 78.586 9.885 78.813 ;
      RECT MASK 2 12.273 78.586 12.353 78.813 ;
      RECT MASK 2 12.605 78.586 12.685 78.813 ;
      RECT MASK 2 12.937 78.586 13.017 78.813 ;
      RECT MASK 2 13.435 78.586 13.515 78.813 ;
      RECT MASK 2 13.767 78.586 13.847 78.813 ;
      RECT MASK 2 14.099 78.586 14.179 78.813 ;
      RECT MASK 2 14.597 78.586 14.677 78.813 ;
      RECT MASK 2 14.929 78.586 15.009 78.813 ;
      RECT MASK 2 15.261 78.586 15.341 78.813 ;
      RECT MASK 2 15.759 78.586 15.839 78.813 ;
      RECT MASK 2 16.091 78.586 16.171 78.813 ;
      RECT MASK 2 16.423 78.586 16.503 78.813 ;
      RECT MASK 2 18.891 78.586 18.971 78.813 ;
      RECT MASK 2 19.223 78.586 19.303 78.813 ;
      RECT MASK 2 19.555 78.586 19.635 78.813 ;
      RECT MASK 2 20.053 78.586 20.133 78.813 ;
      RECT MASK 2 20.385 78.586 20.465 78.813 ;
      RECT MASK 2 20.717 78.586 20.797 78.813 ;
      RECT MASK 2 21.215 78.586 21.295 78.813 ;
      RECT MASK 2 21.547 78.586 21.627 78.813 ;
      RECT MASK 2 21.879 78.586 21.959 78.813 ;
      RECT MASK 2 22.377 78.586 22.457 78.813 ;
      RECT MASK 2 22.709 78.586 22.789 78.813 ;
      RECT MASK 2 23.041 78.586 23.121 78.813 ;
      RECT MASK 2 25.509 78.586 25.589 78.813 ;
      RECT MASK 2 25.841 78.586 25.921 78.813 ;
      RECT MASK 2 26.173 78.586 26.253 78.813 ;
      RECT MASK 2 26.671 78.586 26.751 78.813 ;
      RECT MASK 2 27.003 78.586 27.083 78.813 ;
      RECT MASK 2 27.335 78.586 27.415 78.813 ;
      RECT MASK 2 27.833 78.586 27.913 78.813 ;
      RECT MASK 2 28.165 78.586 28.245 78.813 ;
      RECT MASK 2 28.497 78.586 28.577 78.813 ;
      RECT MASK 2 28.995 78.586 29.075 78.813 ;
      RECT MASK 2 29.327 78.586 29.407 78.813 ;
      RECT MASK 2 29.659 78.586 29.739 78.813 ;
      RECT MASK 2 32.127 78.586 32.207 78.813 ;
      RECT MASK 2 32.459 78.586 32.539 78.813 ;
      RECT MASK 2 32.791 78.586 32.871 78.813 ;
      RECT MASK 2 33.289 78.586 33.369 78.813 ;
      RECT MASK 2 33.621 78.586 33.701 78.813 ;
      RECT MASK 2 33.953 78.586 34.033 78.813 ;
      RECT MASK 2 34.451 78.586 34.531 78.813 ;
      RECT MASK 2 34.783 78.586 34.863 78.813 ;
      RECT MASK 2 35.115 78.586 35.195 78.813 ;
      RECT MASK 2 35.613 78.586 35.693 78.813 ;
      RECT MASK 2 35.945 78.586 36.025 78.813 ;
      RECT MASK 2 36.277 78.586 36.357 78.813 ;
      RECT MASK 2 38.745 78.586 38.825 78.813 ;
      RECT MASK 2 39.077 78.586 39.157 78.813 ;
      RECT MASK 2 39.409 78.586 39.489 78.813 ;
      RECT MASK 2 39.907 78.586 39.987 78.813 ;
      RECT MASK 2 40.239 78.586 40.319 78.813 ;
      RECT MASK 2 40.571 78.586 40.651 78.813 ;
      RECT MASK 2 41.069 78.586 41.149 78.813 ;
      RECT MASK 2 41.401 78.586 41.481 78.813 ;
      RECT MASK 2 41.733 78.586 41.813 78.813 ;
      RECT MASK 2 42.231 78.586 42.311 78.813 ;
      RECT MASK 2 42.563 78.586 42.643 78.813 ;
      RECT MASK 2 42.895 78.586 42.975 78.813 ;
      RECT MASK 2 45.363 78.586 45.443 78.813 ;
      RECT MASK 2 45.695 78.586 45.775 78.813 ;
      RECT MASK 2 46.027 78.586 46.107 78.813 ;
      RECT MASK 2 46.525 78.586 46.605 78.813 ;
      RECT MASK 2 46.857 78.586 46.937 78.813 ;
      RECT MASK 2 47.189 78.586 47.269 78.813 ;
      RECT MASK 2 47.687 78.586 47.767 78.813 ;
      RECT MASK 2 48.019 78.586 48.099 78.813 ;
      RECT MASK 2 48.351 78.586 48.431 78.813 ;
      RECT MASK 2 48.849 78.586 48.929 78.813 ;
      RECT MASK 2 49.181 78.586 49.261 78.813 ;
      RECT MASK 2 49.513 78.586 49.593 78.813 ;
      RECT MASK 2 51.981 78.586 52.061 78.813 ;
      RECT MASK 2 52.313 78.586 52.393 78.813 ;
      RECT MASK 2 52.645 78.586 52.725 78.813 ;
      RECT MASK 2 53.143 78.586 53.223 78.813 ;
      RECT MASK 2 53.475 78.586 53.555 78.813 ;
      RECT MASK 2 53.807 78.586 53.887 78.813 ;
      RECT MASK 2 54.305 78.586 54.385 78.813 ;
      RECT MASK 2 54.637 78.586 54.717 78.813 ;
      RECT MASK 2 54.969 78.586 55.049 78.813 ;
      RECT MASK 2 55.467 78.586 55.547 78.813 ;
      RECT MASK 2 55.799 78.586 55.879 78.813 ;
      RECT MASK 2 56.131 78.586 56.211 78.813 ;
      RECT MASK 2 58.599 78.586 58.679 78.813 ;
      RECT MASK 2 58.931 78.586 59.011 78.813 ;
      RECT MASK 2 59.263 78.586 59.343 78.813 ;
      RECT MASK 2 59.761 78.586 59.841 78.813 ;
      RECT MASK 2 60.093 78.586 60.173 78.813 ;
      RECT MASK 2 60.425 78.586 60.505 78.813 ;
      RECT MASK 2 60.923 78.586 61.003 78.813 ;
      RECT MASK 2 61.255 78.586 61.335 78.813 ;
      RECT MASK 2 61.587 78.586 61.667 78.813 ;
      RECT MASK 2 62.085 78.586 62.165 78.813 ;
      RECT MASK 2 62.417 78.586 62.497 78.813 ;
      RECT MASK 2 62.749 78.586 62.829 78.813 ;
      RECT MASK 2 65.217 78.586 65.297 78.813 ;
      RECT MASK 2 65.549 78.586 65.629 78.813 ;
      RECT MASK 2 65.881 78.586 65.961 78.813 ;
      RECT MASK 2 66.379 78.586 66.459 78.813 ;
      RECT MASK 2 66.711 78.586 66.791 78.813 ;
      RECT MASK 2 67.043 78.586 67.123 78.813 ;
      RECT MASK 2 67.541 78.586 67.621 78.813 ;
      RECT MASK 2 67.873 78.586 67.953 78.813 ;
      RECT MASK 2 68.205 78.586 68.285 78.813 ;
      RECT MASK 2 68.703 78.586 68.783 78.813 ;
      RECT MASK 2 69.035 78.586 69.115 78.813 ;
      RECT MASK 2 69.367 78.586 69.447 78.813 ;
      RECT MASK 2 71.835 78.586 71.915 78.813 ;
      RECT MASK 2 72.167 78.586 72.247 78.813 ;
      RECT MASK 2 72.499 78.586 72.579 78.813 ;
      RECT MASK 2 72.997 78.586 73.077 78.813 ;
      RECT MASK 2 73.329 78.586 73.409 78.813 ;
      RECT MASK 2 73.661 78.586 73.741 78.813 ;
      RECT MASK 2 74.159 78.586 74.239 78.813 ;
      RECT MASK 2 74.491 78.586 74.571 78.813 ;
      RECT MASK 2 74.823 78.586 74.903 78.813 ;
      RECT MASK 2 75.321 78.586 75.401 78.813 ;
      RECT MASK 2 75.653 78.586 75.733 78.813 ;
      RECT MASK 2 75.985 78.586 76.065 78.813 ;
      RECT MASK 2 78.453 78.586 78.533 78.813 ;
      RECT MASK 2 78.785 78.586 78.865 78.813 ;
      RECT MASK 2 79.117 78.586 79.197 78.813 ;
      RECT MASK 2 79.615 78.586 79.695 78.813 ;
      RECT MASK 2 79.947 78.586 80.027 78.813 ;
      RECT MASK 2 80.279 78.586 80.359 78.813 ;
      RECT MASK 2 80.777 78.586 80.857 78.813 ;
      RECT MASK 2 81.109 78.586 81.189 78.813 ;
      RECT MASK 2 81.441 78.586 81.521 78.813 ;
      RECT MASK 2 81.939 78.586 82.019 78.813 ;
      RECT MASK 2 82.271 78.586 82.351 78.813 ;
      RECT MASK 2 82.603 78.586 82.683 78.813 ;
      RECT MASK 2 85.071 78.586 85.151 78.813 ;
      RECT MASK 2 85.403 78.586 85.483 78.813 ;
      RECT MASK 2 85.735 78.586 85.815 78.813 ;
      RECT MASK 2 86.233 78.586 86.313 78.813 ;
      RECT MASK 2 86.565 78.586 86.645 78.813 ;
      RECT MASK 2 86.897 78.586 86.977 78.813 ;
      RECT MASK 2 87.395 78.586 87.475 78.813 ;
      RECT MASK 2 87.727 78.586 87.807 78.813 ;
      RECT MASK 2 88.059 78.586 88.139 78.813 ;
      RECT MASK 2 88.557 78.586 88.637 78.813 ;
      RECT MASK 2 88.889 78.586 88.969 78.813 ;
      RECT MASK 2 89.221 78.586 89.301 78.813 ;
      RECT MASK 2 91.689 78.586 91.769 78.813 ;
      RECT MASK 2 92.021 78.586 92.101 78.813 ;
      RECT MASK 2 92.353 78.586 92.433 78.813 ;
      RECT MASK 2 92.851 78.586 92.931 78.813 ;
      RECT MASK 2 93.183 78.586 93.263 78.813 ;
      RECT MASK 2 93.515 78.586 93.595 78.813 ;
      RECT MASK 2 94.013 78.586 94.093 78.813 ;
      RECT MASK 2 94.345 78.586 94.425 78.813 ;
      RECT MASK 2 94.677 78.586 94.757 78.813 ;
      RECT MASK 2 95.175 78.586 95.255 78.813 ;
      RECT MASK 2 95.507 78.586 95.587 78.813 ;
      RECT MASK 2 95.839 78.586 95.919 78.813 ;
      RECT MASK 2 98.307 78.586 98.387 78.813 ;
      RECT MASK 2 98.639 78.586 98.719 78.813 ;
      RECT MASK 2 98.971 78.586 99.051 78.813 ;
      RECT MASK 2 99.469 78.586 99.549 78.813 ;
      RECT MASK 2 99.801 78.586 99.881 78.813 ;
      RECT MASK 2 100.133 78.586 100.213 78.813 ;
      RECT MASK 2 100.631 78.586 100.711 78.813 ;
      RECT MASK 2 100.963 78.586 101.043 78.813 ;
      RECT MASK 2 101.295 78.586 101.375 78.813 ;
      RECT MASK 2 101.793 78.586 101.873 78.813 ;
      RECT MASK 2 102.125 78.586 102.205 78.813 ;
      RECT MASK 2 102.457 78.586 102.537 78.813 ;
      RECT MASK 2 104.925 78.586 105.005 78.813 ;
      RECT MASK 2 105.257 78.586 105.337 78.813 ;
      RECT MASK 2 105.589 78.586 105.669 78.813 ;
      RECT MASK 2 106.087 78.586 106.167 78.813 ;
      RECT MASK 2 106.419 78.586 106.499 78.813 ;
      RECT MASK 2 106.751 78.586 106.831 78.813 ;
      RECT MASK 2 107.249 78.586 107.329 78.813 ;
      RECT MASK 2 107.581 78.586 107.661 78.813 ;
      RECT MASK 2 107.913 78.586 107.993 78.813 ;
      RECT MASK 2 108.411 78.586 108.491 78.813 ;
      RECT MASK 2 108.743 78.586 108.823 78.813 ;
      RECT MASK 2 109.075 78.586 109.155 78.813 ;
      RECT MASK 2 116.437 78.668 116.497 78.892 ;
      RECT MASK 2 116.769 78.668 116.829 78.892 ;
      RECT MASK 2 117.101 78.668 117.161 78.892 ;
      RECT MASK 2 117.433 78.668 117.493 78.892 ;
      RECT MASK 2 117.765 78.668 117.825 78.892 ;
      RECT MASK 2 118.097 78.668 118.157 78.892 ;
      RECT MASK 2 118.429 78.668 118.489 78.892 ;
      RECT MASK 2 118.761 78.668 118.821 78.892 ;
      RECT MASK 2 119.093 78.668 119.153 78.892 ;
      RECT MASK 2 119.425 78.668 119.485 78.892 ;
      RECT MASK 2 119.757 78.668 119.817 78.892 ;
      RECT MASK 2 120.089 78.668 120.149 78.892 ;
      RECT MASK 2 120.421 78.668 120.481 78.892 ;
      RECT MASK 2 120.753 78.668 120.813 78.892 ;
      RECT MASK 2 121.085 78.668 121.145 78.892 ;
      RECT MASK 2 121.417 78.668 121.477 78.892 ;
      RECT MASK 2 121.749 78.668 121.809 78.892 ;
      RECT MASK 2 122.081 78.668 122.141 78.892 ;
      RECT MASK 2 122.413 78.668 122.473 78.892 ;
      RECT MASK 2 122.745 78.668 122.805 78.892 ;
      RECT MASK 2 123.077 78.668 123.137 78.892 ;
      RECT MASK 2 123.409 78.668 123.469 78.892 ;
      RECT MASK 2 123.741 78.668 123.801 78.892 ;
      RECT MASK 2 124.073 78.668 124.133 78.892 ;
      RECT MASK 2 124.405 78.668 124.465 78.892 ;
      RECT MASK 2 124.737 78.668 124.797 78.892 ;
      RECT MASK 2 125.069 78.668 125.129 78.892 ;
      RECT MASK 2 125.401 78.668 125.461 78.892 ;
      RECT MASK 2 125.733 78.668 125.793 78.892 ;
      RECT MASK 2 126.065 78.668 126.125 78.892 ;
      RECT MASK 2 1.248 78.75 5.362 78.79 ;
      RECT MASK 2 111.186 78.8 113.288 78.84 ;
      RECT MASK 2 10.873 78.9455 10.953 79.217 ;
      RECT MASK 2 11.205 78.9455 11.285 79.217 ;
      RECT MASK 2 17.491 78.9455 17.571 79.217 ;
      RECT MASK 2 17.823 78.9455 17.903 79.217 ;
      RECT MASK 2 24.109 78.9455 24.189 79.217 ;
      RECT MASK 2 24.441 78.9455 24.521 79.217 ;
      RECT MASK 2 30.727 78.9455 30.807 79.217 ;
      RECT MASK 2 31.059 78.9455 31.139 79.217 ;
      RECT MASK 2 37.345 78.9455 37.425 79.217 ;
      RECT MASK 2 37.677 78.9455 37.757 79.217 ;
      RECT MASK 2 43.963 78.9455 44.043 79.217 ;
      RECT MASK 2 44.295 78.9455 44.375 79.217 ;
      RECT MASK 2 50.581 78.9455 50.661 79.217 ;
      RECT MASK 2 50.913 78.9455 50.993 79.217 ;
      RECT MASK 2 57.199 78.9455 57.279 79.217 ;
      RECT MASK 2 57.531 78.9455 57.611 79.217 ;
      RECT MASK 2 63.817 78.9455 63.897 79.217 ;
      RECT MASK 2 64.149 78.9455 64.229 79.217 ;
      RECT MASK 2 70.435 78.9455 70.515 79.217 ;
      RECT MASK 2 70.767 78.9455 70.847 79.217 ;
      RECT MASK 2 77.053 78.9455 77.133 79.217 ;
      RECT MASK 2 77.385 78.9455 77.465 79.217 ;
      RECT MASK 2 83.671 78.9455 83.751 79.217 ;
      RECT MASK 2 84.003 78.9455 84.083 79.217 ;
      RECT MASK 2 90.289 78.9455 90.369 79.217 ;
      RECT MASK 2 90.621 78.9455 90.701 79.217 ;
      RECT MASK 2 96.907 78.9455 96.987 79.217 ;
      RECT MASK 2 97.239 78.9455 97.319 79.217 ;
      RECT MASK 2 103.525 78.9455 103.605 79.217 ;
      RECT MASK 2 103.857 78.9455 103.937 79.217 ;
      RECT MASK 2 111.186 78.99 113.288 79.03 ;
      RECT MASK 2 116.079 79.1125 116.2725 79.1525 ;
      RECT MASK 2 126.2895 79.1125 126.483 79.1525 ;
      RECT MASK 2 6.817 79.2515 6.897 79.478 ;
      RECT MASK 2 7.149 79.2515 7.229 79.478 ;
      RECT MASK 2 7.481 79.2515 7.561 79.478 ;
      RECT MASK 2 7.979 79.2515 8.059 79.478 ;
      RECT MASK 2 8.311 79.2515 8.391 79.478 ;
      RECT MASK 2 8.643 79.2515 8.723 79.478 ;
      RECT MASK 2 9.141 79.2515 9.221 79.478 ;
      RECT MASK 2 9.473 79.2515 9.553 79.478 ;
      RECT MASK 2 9.805 79.2515 9.885 79.478 ;
      RECT MASK 2 12.273 79.2515 12.353 79.478 ;
      RECT MASK 2 12.605 79.2515 12.685 79.478 ;
      RECT MASK 2 12.937 79.2515 13.017 79.478 ;
      RECT MASK 2 13.435 79.2515 13.515 79.478 ;
      RECT MASK 2 13.767 79.2515 13.847 79.478 ;
      RECT MASK 2 14.099 79.2515 14.179 79.478 ;
      RECT MASK 2 14.597 79.2515 14.677 79.478 ;
      RECT MASK 2 14.929 79.2515 15.009 79.478 ;
      RECT MASK 2 15.261 79.2515 15.341 79.478 ;
      RECT MASK 2 15.759 79.2515 15.839 79.478 ;
      RECT MASK 2 16.091 79.2515 16.171 79.478 ;
      RECT MASK 2 16.423 79.2515 16.503 79.478 ;
      RECT MASK 2 18.891 79.2515 18.971 79.478 ;
      RECT MASK 2 19.223 79.2515 19.303 79.478 ;
      RECT MASK 2 19.555 79.2515 19.635 79.478 ;
      RECT MASK 2 20.053 79.2515 20.133 79.478 ;
      RECT MASK 2 20.385 79.2515 20.465 79.478 ;
      RECT MASK 2 20.717 79.2515 20.797 79.478 ;
      RECT MASK 2 21.215 79.2515 21.295 79.478 ;
      RECT MASK 2 21.547 79.2515 21.627 79.478 ;
      RECT MASK 2 21.879 79.2515 21.959 79.478 ;
      RECT MASK 2 22.377 79.2515 22.457 79.478 ;
      RECT MASK 2 22.709 79.2515 22.789 79.478 ;
      RECT MASK 2 23.041 79.2515 23.121 79.478 ;
      RECT MASK 2 25.509 79.2515 25.589 79.478 ;
      RECT MASK 2 25.841 79.2515 25.921 79.478 ;
      RECT MASK 2 26.173 79.2515 26.253 79.478 ;
      RECT MASK 2 26.671 79.2515 26.751 79.478 ;
      RECT MASK 2 27.003 79.2515 27.083 79.478 ;
      RECT MASK 2 27.335 79.2515 27.415 79.478 ;
      RECT MASK 2 27.833 79.2515 27.913 79.478 ;
      RECT MASK 2 28.165 79.2515 28.245 79.478 ;
      RECT MASK 2 28.497 79.2515 28.577 79.478 ;
      RECT MASK 2 28.995 79.2515 29.075 79.478 ;
      RECT MASK 2 29.327 79.2515 29.407 79.478 ;
      RECT MASK 2 29.659 79.2515 29.739 79.478 ;
      RECT MASK 2 32.127 79.2515 32.207 79.478 ;
      RECT MASK 2 32.459 79.2515 32.539 79.478 ;
      RECT MASK 2 32.791 79.2515 32.871 79.478 ;
      RECT MASK 2 33.289 79.2515 33.369 79.478 ;
      RECT MASK 2 33.621 79.2515 33.701 79.478 ;
      RECT MASK 2 33.953 79.2515 34.033 79.478 ;
      RECT MASK 2 34.451 79.2515 34.531 79.478 ;
      RECT MASK 2 34.783 79.2515 34.863 79.478 ;
      RECT MASK 2 35.115 79.2515 35.195 79.478 ;
      RECT MASK 2 35.613 79.2515 35.693 79.478 ;
      RECT MASK 2 35.945 79.2515 36.025 79.478 ;
      RECT MASK 2 36.277 79.2515 36.357 79.478 ;
      RECT MASK 2 38.745 79.2515 38.825 79.478 ;
      RECT MASK 2 39.077 79.2515 39.157 79.478 ;
      RECT MASK 2 39.409 79.2515 39.489 79.478 ;
      RECT MASK 2 39.907 79.2515 39.987 79.478 ;
      RECT MASK 2 40.239 79.2515 40.319 79.478 ;
      RECT MASK 2 40.571 79.2515 40.651 79.478 ;
      RECT MASK 2 41.069 79.2515 41.149 79.478 ;
      RECT MASK 2 41.401 79.2515 41.481 79.478 ;
      RECT MASK 2 41.733 79.2515 41.813 79.478 ;
      RECT MASK 2 42.231 79.2515 42.311 79.478 ;
      RECT MASK 2 42.563 79.2515 42.643 79.478 ;
      RECT MASK 2 42.895 79.2515 42.975 79.478 ;
      RECT MASK 2 45.363 79.2515 45.443 79.478 ;
      RECT MASK 2 45.695 79.2515 45.775 79.478 ;
      RECT MASK 2 46.027 79.2515 46.107 79.478 ;
      RECT MASK 2 46.525 79.2515 46.605 79.478 ;
      RECT MASK 2 46.857 79.2515 46.937 79.478 ;
      RECT MASK 2 47.189 79.2515 47.269 79.478 ;
      RECT MASK 2 47.687 79.2515 47.767 79.478 ;
      RECT MASK 2 48.019 79.2515 48.099 79.478 ;
      RECT MASK 2 48.351 79.2515 48.431 79.478 ;
      RECT MASK 2 48.849 79.2515 48.929 79.478 ;
      RECT MASK 2 49.181 79.2515 49.261 79.478 ;
      RECT MASK 2 49.513 79.2515 49.593 79.478 ;
      RECT MASK 2 51.981 79.2515 52.061 79.478 ;
      RECT MASK 2 52.313 79.2515 52.393 79.478 ;
      RECT MASK 2 52.645 79.2515 52.725 79.478 ;
      RECT MASK 2 53.143 79.2515 53.223 79.478 ;
      RECT MASK 2 53.475 79.2515 53.555 79.478 ;
      RECT MASK 2 53.807 79.2515 53.887 79.478 ;
      RECT MASK 2 54.305 79.2515 54.385 79.478 ;
      RECT MASK 2 54.637 79.2515 54.717 79.478 ;
      RECT MASK 2 54.969 79.2515 55.049 79.478 ;
      RECT MASK 2 55.467 79.2515 55.547 79.478 ;
      RECT MASK 2 55.799 79.2515 55.879 79.478 ;
      RECT MASK 2 56.131 79.2515 56.211 79.478 ;
      RECT MASK 2 58.599 79.2515 58.679 79.478 ;
      RECT MASK 2 58.931 79.2515 59.011 79.478 ;
      RECT MASK 2 59.263 79.2515 59.343 79.478 ;
      RECT MASK 2 59.761 79.2515 59.841 79.478 ;
      RECT MASK 2 60.093 79.2515 60.173 79.478 ;
      RECT MASK 2 60.425 79.2515 60.505 79.478 ;
      RECT MASK 2 60.923 79.2515 61.003 79.478 ;
      RECT MASK 2 61.255 79.2515 61.335 79.478 ;
      RECT MASK 2 61.587 79.2515 61.667 79.478 ;
      RECT MASK 2 62.085 79.2515 62.165 79.478 ;
      RECT MASK 2 62.417 79.2515 62.497 79.478 ;
      RECT MASK 2 62.749 79.2515 62.829 79.478 ;
      RECT MASK 2 65.217 79.2515 65.297 79.478 ;
      RECT MASK 2 65.549 79.2515 65.629 79.478 ;
      RECT MASK 2 65.881 79.2515 65.961 79.478 ;
      RECT MASK 2 66.379 79.2515 66.459 79.478 ;
      RECT MASK 2 66.711 79.2515 66.791 79.478 ;
      RECT MASK 2 67.043 79.2515 67.123 79.478 ;
      RECT MASK 2 67.541 79.2515 67.621 79.478 ;
      RECT MASK 2 67.873 79.2515 67.953 79.478 ;
      RECT MASK 2 68.205 79.2515 68.285 79.478 ;
      RECT MASK 2 68.703 79.2515 68.783 79.478 ;
      RECT MASK 2 69.035 79.2515 69.115 79.478 ;
      RECT MASK 2 69.367 79.2515 69.447 79.478 ;
      RECT MASK 2 71.835 79.2515 71.915 79.478 ;
      RECT MASK 2 72.167 79.2515 72.247 79.478 ;
      RECT MASK 2 72.499 79.2515 72.579 79.478 ;
      RECT MASK 2 72.997 79.2515 73.077 79.478 ;
      RECT MASK 2 73.329 79.2515 73.409 79.478 ;
      RECT MASK 2 73.661 79.2515 73.741 79.478 ;
      RECT MASK 2 74.159 79.2515 74.239 79.478 ;
      RECT MASK 2 74.491 79.2515 74.571 79.478 ;
      RECT MASK 2 74.823 79.2515 74.903 79.478 ;
      RECT MASK 2 75.321 79.2515 75.401 79.478 ;
      RECT MASK 2 75.653 79.2515 75.733 79.478 ;
      RECT MASK 2 75.985 79.2515 76.065 79.478 ;
      RECT MASK 2 78.453 79.2515 78.533 79.478 ;
      RECT MASK 2 78.785 79.2515 78.865 79.478 ;
      RECT MASK 2 79.117 79.2515 79.197 79.478 ;
      RECT MASK 2 79.615 79.2515 79.695 79.478 ;
      RECT MASK 2 79.947 79.2515 80.027 79.478 ;
      RECT MASK 2 80.279 79.2515 80.359 79.478 ;
      RECT MASK 2 80.777 79.2515 80.857 79.478 ;
      RECT MASK 2 81.109 79.2515 81.189 79.478 ;
      RECT MASK 2 81.441 79.2515 81.521 79.478 ;
      RECT MASK 2 81.939 79.2515 82.019 79.478 ;
      RECT MASK 2 82.271 79.2515 82.351 79.478 ;
      RECT MASK 2 82.603 79.2515 82.683 79.478 ;
      RECT MASK 2 85.071 79.2515 85.151 79.478 ;
      RECT MASK 2 85.403 79.2515 85.483 79.478 ;
      RECT MASK 2 85.735 79.2515 85.815 79.478 ;
      RECT MASK 2 86.233 79.2515 86.313 79.478 ;
      RECT MASK 2 86.565 79.2515 86.645 79.478 ;
      RECT MASK 2 86.897 79.2515 86.977 79.478 ;
      RECT MASK 2 87.395 79.2515 87.475 79.478 ;
      RECT MASK 2 87.727 79.2515 87.807 79.478 ;
      RECT MASK 2 88.059 79.2515 88.139 79.478 ;
      RECT MASK 2 88.557 79.2515 88.637 79.478 ;
      RECT MASK 2 88.889 79.2515 88.969 79.478 ;
      RECT MASK 2 89.221 79.2515 89.301 79.478 ;
      RECT MASK 2 91.689 79.2515 91.769 79.478 ;
      RECT MASK 2 92.021 79.2515 92.101 79.478 ;
      RECT MASK 2 92.353 79.2515 92.433 79.478 ;
      RECT MASK 2 92.851 79.2515 92.931 79.478 ;
      RECT MASK 2 93.183 79.2515 93.263 79.478 ;
      RECT MASK 2 93.515 79.2515 93.595 79.478 ;
      RECT MASK 2 94.013 79.2515 94.093 79.478 ;
      RECT MASK 2 94.345 79.2515 94.425 79.478 ;
      RECT MASK 2 94.677 79.2515 94.757 79.478 ;
      RECT MASK 2 95.175 79.2515 95.255 79.478 ;
      RECT MASK 2 95.507 79.2515 95.587 79.478 ;
      RECT MASK 2 95.839 79.2515 95.919 79.478 ;
      RECT MASK 2 98.307 79.2515 98.387 79.478 ;
      RECT MASK 2 98.639 79.2515 98.719 79.478 ;
      RECT MASK 2 98.971 79.2515 99.051 79.478 ;
      RECT MASK 2 99.469 79.2515 99.549 79.478 ;
      RECT MASK 2 99.801 79.2515 99.881 79.478 ;
      RECT MASK 2 100.133 79.2515 100.213 79.478 ;
      RECT MASK 2 100.631 79.2515 100.711 79.478 ;
      RECT MASK 2 100.963 79.2515 101.043 79.478 ;
      RECT MASK 2 101.295 79.2515 101.375 79.478 ;
      RECT MASK 2 101.793 79.2515 101.873 79.478 ;
      RECT MASK 2 102.125 79.2515 102.205 79.478 ;
      RECT MASK 2 102.457 79.2515 102.537 79.478 ;
      RECT MASK 2 104.925 79.2515 105.005 79.478 ;
      RECT MASK 2 105.257 79.2515 105.337 79.478 ;
      RECT MASK 2 105.589 79.2515 105.669 79.478 ;
      RECT MASK 2 106.087 79.2515 106.167 79.478 ;
      RECT MASK 2 106.419 79.2515 106.499 79.478 ;
      RECT MASK 2 106.751 79.2515 106.831 79.478 ;
      RECT MASK 2 107.249 79.2515 107.329 79.478 ;
      RECT MASK 2 107.581 79.2515 107.661 79.478 ;
      RECT MASK 2 107.913 79.2515 107.993 79.478 ;
      RECT MASK 2 108.411 79.2515 108.491 79.478 ;
      RECT MASK 2 108.743 79.2515 108.823 79.478 ;
      RECT MASK 2 109.075 79.2515 109.155 79.478 ;
      RECT MASK 2 2.204 79.26 2.264 80.31 ;
      RECT MASK 2 2.478 79.26 2.538 80.31 ;
      RECT MASK 2 2.752 79.26 2.812 80.31 ;
      RECT MASK 2 3.026 79.26 3.086 80.31 ;
      RECT MASK 2 3.3 79.26 3.36 80.31 ;
      RECT MASK 2 3.574 79.26 3.634 80.31 ;
      RECT MASK 2 3.848 79.26 3.908 80.31 ;
      RECT MASK 2 4.122 79.26 4.182 80.31 ;
      RECT MASK 2 4.396 79.26 4.456 80.31 ;
      RECT MASK 2 111.122 79.331 113.352 79.371 ;
      RECT MASK 2 116.437 79.448 116.497 79.672 ;
      RECT MASK 2 116.769 79.448 116.829 79.672 ;
      RECT MASK 2 117.101 79.448 117.161 79.672 ;
      RECT MASK 2 117.433 79.448 117.493 79.672 ;
      RECT MASK 2 117.765 79.448 117.825 79.672 ;
      RECT MASK 2 118.097 79.448 118.157 79.672 ;
      RECT MASK 2 118.429 79.448 118.489 79.672 ;
      RECT MASK 2 118.761 79.448 118.821 79.672 ;
      RECT MASK 2 119.093 79.448 119.153 79.672 ;
      RECT MASK 2 119.425 79.448 119.485 79.672 ;
      RECT MASK 2 119.757 79.448 119.817 79.672 ;
      RECT MASK 2 120.089 79.448 120.149 79.672 ;
      RECT MASK 2 120.421 79.448 120.481 79.672 ;
      RECT MASK 2 120.753 79.448 120.813 79.672 ;
      RECT MASK 2 121.085 79.448 121.145 79.672 ;
      RECT MASK 2 121.417 79.448 121.477 79.672 ;
      RECT MASK 2 121.749 79.448 121.809 79.672 ;
      RECT MASK 2 122.081 79.448 122.141 79.672 ;
      RECT MASK 2 122.413 79.448 122.473 79.672 ;
      RECT MASK 2 122.745 79.448 122.805 79.672 ;
      RECT MASK 2 123.077 79.448 123.137 79.672 ;
      RECT MASK 2 123.409 79.448 123.469 79.672 ;
      RECT MASK 2 123.741 79.448 123.801 79.672 ;
      RECT MASK 2 124.073 79.448 124.133 79.672 ;
      RECT MASK 2 124.405 79.448 124.465 79.672 ;
      RECT MASK 2 124.737 79.448 124.797 79.672 ;
      RECT MASK 2 125.069 79.448 125.129 79.672 ;
      RECT MASK 2 125.401 79.448 125.461 79.672 ;
      RECT MASK 2 125.733 79.448 125.793 79.672 ;
      RECT MASK 2 126.065 79.448 126.125 79.672 ;
      RECT MASK 2 111.122 79.499 113.352 79.539 ;
      RECT MASK 2 111.767 79.683 111.95 79.723 ;
      RECT MASK 2 112.431 79.683 112.614 79.723 ;
      RECT MASK 2 116.079 79.8925 116.2725 79.9325 ;
      RECT MASK 2 126.2895 79.8925 126.483 79.9325 ;
      RECT MASK 2 111.151 79.905 111.331 79.945 ;
      RECT MASK 2 113.143 79.905 113.323 79.945 ;
      RECT MASK 2 6.2775 80 110.065 80.04 ;
      RECT MASK 2 115.539 80.18 126.947 80.22 ;
      RECT MASK 2 6.2775 80.19 110.065 80.23 ;
      RECT MASK 2 111.186 80.315 113.288 80.355 ;
      RECT MASK 2 115.539 80.37 126.947 80.41 ;
      RECT MASK 2 6.2775 80.45 109.836 80.49 ;
      RECT MASK 2 6.2775 80.64 109.836 80.68 ;
      RECT MASK 2 111.186 80.835 113.288 80.875 ;
      RECT MASK 2 2.204 80.97 2.264 82.02 ;
      RECT MASK 2 2.478 80.97 2.538 82.02 ;
      RECT MASK 2 2.752 80.97 2.812 82.02 ;
      RECT MASK 2 3.026 80.97 3.086 82.02 ;
      RECT MASK 2 3.3 80.97 3.36 82.02 ;
      RECT MASK 2 3.574 80.97 3.634 82.02 ;
      RECT MASK 2 3.848 80.97 3.908 82.02 ;
      RECT MASK 2 4.122 80.97 4.182 82.02 ;
      RECT MASK 2 4.396 80.97 4.456 82.02 ;
      RECT MASK 2 6.817 80.986 6.897 81.211 ;
      RECT MASK 2 7.149 80.986 7.229 81.211 ;
      RECT MASK 2 7.481 80.986 7.561 81.211 ;
      RECT MASK 2 7.979 80.986 8.059 81.211 ;
      RECT MASK 2 8.311 80.986 8.391 81.211 ;
      RECT MASK 2 8.643 80.986 8.723 81.211 ;
      RECT MASK 2 9.141 80.986 9.221 81.211 ;
      RECT MASK 2 9.473 80.986 9.553 81.211 ;
      RECT MASK 2 9.805 80.986 9.885 81.211 ;
      RECT MASK 2 12.273 80.986 12.353 81.211 ;
      RECT MASK 2 12.605 80.986 12.685 81.211 ;
      RECT MASK 2 12.937 80.986 13.017 81.211 ;
      RECT MASK 2 13.435 80.986 13.515 81.211 ;
      RECT MASK 2 13.767 80.986 13.847 81.211 ;
      RECT MASK 2 14.099 80.986 14.179 81.211 ;
      RECT MASK 2 14.597 80.986 14.677 81.211 ;
      RECT MASK 2 14.929 80.986 15.009 81.211 ;
      RECT MASK 2 15.261 80.986 15.341 81.211 ;
      RECT MASK 2 15.759 80.986 15.839 81.211 ;
      RECT MASK 2 16.091 80.986 16.171 81.211 ;
      RECT MASK 2 16.423 80.986 16.503 81.211 ;
      RECT MASK 2 18.891 80.986 18.971 81.211 ;
      RECT MASK 2 19.223 80.986 19.303 81.211 ;
      RECT MASK 2 19.555 80.986 19.635 81.211 ;
      RECT MASK 2 20.053 80.986 20.133 81.211 ;
      RECT MASK 2 20.385 80.986 20.465 81.211 ;
      RECT MASK 2 20.717 80.986 20.797 81.211 ;
      RECT MASK 2 21.215 80.986 21.295 81.211 ;
      RECT MASK 2 21.547 80.986 21.627 81.211 ;
      RECT MASK 2 21.879 80.986 21.959 81.211 ;
      RECT MASK 2 22.377 80.986 22.457 81.211 ;
      RECT MASK 2 22.709 80.986 22.789 81.211 ;
      RECT MASK 2 23.041 80.986 23.121 81.211 ;
      RECT MASK 2 25.509 80.986 25.589 81.211 ;
      RECT MASK 2 25.841 80.986 25.921 81.211 ;
      RECT MASK 2 26.173 80.986 26.253 81.211 ;
      RECT MASK 2 26.671 80.986 26.751 81.211 ;
      RECT MASK 2 27.003 80.986 27.083 81.211 ;
      RECT MASK 2 27.335 80.986 27.415 81.211 ;
      RECT MASK 2 27.833 80.986 27.913 81.211 ;
      RECT MASK 2 28.165 80.986 28.245 81.211 ;
      RECT MASK 2 28.497 80.986 28.577 81.211 ;
      RECT MASK 2 28.995 80.986 29.075 81.211 ;
      RECT MASK 2 29.327 80.986 29.407 81.211 ;
      RECT MASK 2 29.659 80.986 29.739 81.211 ;
      RECT MASK 2 32.127 80.986 32.207 81.211 ;
      RECT MASK 2 32.459 80.986 32.539 81.211 ;
      RECT MASK 2 32.791 80.986 32.871 81.211 ;
      RECT MASK 2 33.289 80.986 33.369 81.211 ;
      RECT MASK 2 33.621 80.986 33.701 81.211 ;
      RECT MASK 2 33.953 80.986 34.033 81.211 ;
      RECT MASK 2 34.451 80.986 34.531 81.211 ;
      RECT MASK 2 34.783 80.986 34.863 81.211 ;
      RECT MASK 2 35.115 80.986 35.195 81.211 ;
      RECT MASK 2 35.613 80.986 35.693 81.211 ;
      RECT MASK 2 35.945 80.986 36.025 81.211 ;
      RECT MASK 2 36.277 80.986 36.357 81.211 ;
      RECT MASK 2 38.745 80.986 38.825 81.211 ;
      RECT MASK 2 39.077 80.986 39.157 81.211 ;
      RECT MASK 2 39.409 80.986 39.489 81.211 ;
      RECT MASK 2 39.907 80.986 39.987 81.211 ;
      RECT MASK 2 40.239 80.986 40.319 81.211 ;
      RECT MASK 2 40.571 80.986 40.651 81.211 ;
      RECT MASK 2 41.069 80.986 41.149 81.211 ;
      RECT MASK 2 41.401 80.986 41.481 81.211 ;
      RECT MASK 2 41.733 80.986 41.813 81.211 ;
      RECT MASK 2 42.231 80.986 42.311 81.211 ;
      RECT MASK 2 42.563 80.986 42.643 81.211 ;
      RECT MASK 2 42.895 80.986 42.975 81.211 ;
      RECT MASK 2 45.363 80.986 45.443 81.211 ;
      RECT MASK 2 45.695 80.986 45.775 81.211 ;
      RECT MASK 2 46.027 80.986 46.107 81.211 ;
      RECT MASK 2 46.525 80.986 46.605 81.211 ;
      RECT MASK 2 46.857 80.986 46.937 81.211 ;
      RECT MASK 2 47.189 80.986 47.269 81.211 ;
      RECT MASK 2 47.687 80.986 47.767 81.211 ;
      RECT MASK 2 48.019 80.986 48.099 81.211 ;
      RECT MASK 2 48.351 80.986 48.431 81.211 ;
      RECT MASK 2 48.849 80.986 48.929 81.211 ;
      RECT MASK 2 49.181 80.986 49.261 81.211 ;
      RECT MASK 2 49.513 80.986 49.593 81.211 ;
      RECT MASK 2 51.981 80.986 52.061 81.211 ;
      RECT MASK 2 52.313 80.986 52.393 81.211 ;
      RECT MASK 2 52.645 80.986 52.725 81.211 ;
      RECT MASK 2 53.143 80.986 53.223 81.211 ;
      RECT MASK 2 53.475 80.986 53.555 81.211 ;
      RECT MASK 2 53.807 80.986 53.887 81.211 ;
      RECT MASK 2 54.305 80.986 54.385 81.211 ;
      RECT MASK 2 54.637 80.986 54.717 81.211 ;
      RECT MASK 2 54.969 80.986 55.049 81.211 ;
      RECT MASK 2 55.467 80.986 55.547 81.211 ;
      RECT MASK 2 55.799 80.986 55.879 81.211 ;
      RECT MASK 2 56.131 80.986 56.211 81.211 ;
      RECT MASK 2 58.599 80.986 58.679 81.211 ;
      RECT MASK 2 58.931 80.986 59.011 81.211 ;
      RECT MASK 2 59.263 80.986 59.343 81.211 ;
      RECT MASK 2 59.761 80.986 59.841 81.211 ;
      RECT MASK 2 60.093 80.986 60.173 81.211 ;
      RECT MASK 2 60.425 80.986 60.505 81.211 ;
      RECT MASK 2 60.923 80.986 61.003 81.211 ;
      RECT MASK 2 61.255 80.986 61.335 81.211 ;
      RECT MASK 2 61.587 80.986 61.667 81.211 ;
      RECT MASK 2 62.085 80.986 62.165 81.211 ;
      RECT MASK 2 62.417 80.986 62.497 81.211 ;
      RECT MASK 2 62.749 80.986 62.829 81.211 ;
      RECT MASK 2 65.217 80.986 65.297 81.211 ;
      RECT MASK 2 65.549 80.986 65.629 81.211 ;
      RECT MASK 2 65.881 80.986 65.961 81.211 ;
      RECT MASK 2 66.379 80.986 66.459 81.211 ;
      RECT MASK 2 66.711 80.986 66.791 81.211 ;
      RECT MASK 2 67.043 80.986 67.123 81.211 ;
      RECT MASK 2 67.541 80.986 67.621 81.211 ;
      RECT MASK 2 67.873 80.986 67.953 81.211 ;
      RECT MASK 2 68.205 80.986 68.285 81.211 ;
      RECT MASK 2 68.703 80.986 68.783 81.211 ;
      RECT MASK 2 69.035 80.986 69.115 81.211 ;
      RECT MASK 2 69.367 80.986 69.447 81.211 ;
      RECT MASK 2 71.835 80.986 71.915 81.211 ;
      RECT MASK 2 72.167 80.986 72.247 81.211 ;
      RECT MASK 2 72.499 80.986 72.579 81.211 ;
      RECT MASK 2 72.997 80.986 73.077 81.211 ;
      RECT MASK 2 73.329 80.986 73.409 81.211 ;
      RECT MASK 2 73.661 80.986 73.741 81.211 ;
      RECT MASK 2 74.159 80.986 74.239 81.211 ;
      RECT MASK 2 74.491 80.986 74.571 81.211 ;
      RECT MASK 2 74.823 80.986 74.903 81.211 ;
      RECT MASK 2 75.321 80.986 75.401 81.211 ;
      RECT MASK 2 75.653 80.986 75.733 81.211 ;
      RECT MASK 2 75.985 80.986 76.065 81.211 ;
      RECT MASK 2 78.453 80.986 78.533 81.211 ;
      RECT MASK 2 78.785 80.986 78.865 81.211 ;
      RECT MASK 2 79.117 80.986 79.197 81.211 ;
      RECT MASK 2 79.615 80.986 79.695 81.211 ;
      RECT MASK 2 79.947 80.986 80.027 81.211 ;
      RECT MASK 2 80.279 80.986 80.359 81.211 ;
      RECT MASK 2 80.777 80.986 80.857 81.211 ;
      RECT MASK 2 81.109 80.986 81.189 81.211 ;
      RECT MASK 2 81.441 80.986 81.521 81.211 ;
      RECT MASK 2 81.939 80.986 82.019 81.211 ;
      RECT MASK 2 82.271 80.986 82.351 81.211 ;
      RECT MASK 2 82.603 80.986 82.683 81.211 ;
      RECT MASK 2 85.071 80.986 85.151 81.211 ;
      RECT MASK 2 85.403 80.986 85.483 81.211 ;
      RECT MASK 2 85.735 80.986 85.815 81.211 ;
      RECT MASK 2 86.233 80.986 86.313 81.211 ;
      RECT MASK 2 86.565 80.986 86.645 81.211 ;
      RECT MASK 2 86.897 80.986 86.977 81.211 ;
      RECT MASK 2 87.395 80.986 87.475 81.211 ;
      RECT MASK 2 87.727 80.986 87.807 81.211 ;
      RECT MASK 2 88.059 80.986 88.139 81.211 ;
      RECT MASK 2 88.557 80.986 88.637 81.211 ;
      RECT MASK 2 88.889 80.986 88.969 81.211 ;
      RECT MASK 2 89.221 80.986 89.301 81.211 ;
      RECT MASK 2 91.689 80.986 91.769 81.211 ;
      RECT MASK 2 92.021 80.986 92.101 81.211 ;
      RECT MASK 2 92.353 80.986 92.433 81.211 ;
      RECT MASK 2 92.851 80.986 92.931 81.211 ;
      RECT MASK 2 93.183 80.986 93.263 81.211 ;
      RECT MASK 2 93.515 80.986 93.595 81.211 ;
      RECT MASK 2 94.013 80.986 94.093 81.211 ;
      RECT MASK 2 94.345 80.986 94.425 81.211 ;
      RECT MASK 2 94.677 80.986 94.757 81.211 ;
      RECT MASK 2 95.175 80.986 95.255 81.211 ;
      RECT MASK 2 95.507 80.986 95.587 81.211 ;
      RECT MASK 2 95.839 80.986 95.919 81.211 ;
      RECT MASK 2 98.307 80.986 98.387 81.211 ;
      RECT MASK 2 98.639 80.986 98.719 81.211 ;
      RECT MASK 2 98.971 80.986 99.051 81.211 ;
      RECT MASK 2 99.469 80.986 99.549 81.211 ;
      RECT MASK 2 99.801 80.986 99.881 81.211 ;
      RECT MASK 2 100.133 80.986 100.213 81.211 ;
      RECT MASK 2 100.631 80.986 100.711 81.211 ;
      RECT MASK 2 100.963 80.986 101.043 81.211 ;
      RECT MASK 2 101.295 80.986 101.375 81.211 ;
      RECT MASK 2 101.793 80.986 101.873 81.211 ;
      RECT MASK 2 102.125 80.986 102.205 81.211 ;
      RECT MASK 2 102.457 80.986 102.537 81.211 ;
      RECT MASK 2 104.925 80.986 105.005 81.211 ;
      RECT MASK 2 105.257 80.986 105.337 81.211 ;
      RECT MASK 2 105.589 80.986 105.669 81.211 ;
      RECT MASK 2 106.087 80.986 106.167 81.211 ;
      RECT MASK 2 106.419 80.986 106.499 81.211 ;
      RECT MASK 2 106.751 80.986 106.831 81.211 ;
      RECT MASK 2 107.249 80.986 107.329 81.211 ;
      RECT MASK 2 107.581 80.986 107.661 81.211 ;
      RECT MASK 2 107.913 80.986 107.993 81.211 ;
      RECT MASK 2 108.411 80.986 108.491 81.211 ;
      RECT MASK 2 108.743 80.986 108.823 81.211 ;
      RECT MASK 2 109.075 80.986 109.155 81.211 ;
      RECT MASK 2 111.151 81.281 111.331 81.321 ;
      RECT MASK 2 113.143 81.281 113.323 81.321 ;
      RECT MASK 2 115.613 81.35 128.525 81.39 ;
      RECT MASK 2 10.873 81.463 10.953 81.7345 ;
      RECT MASK 2 11.205 81.463 11.285 81.7345 ;
      RECT MASK 2 17.491 81.463 17.571 81.7345 ;
      RECT MASK 2 17.823 81.463 17.903 81.7345 ;
      RECT MASK 2 24.109 81.463 24.189 81.7345 ;
      RECT MASK 2 24.441 81.463 24.521 81.7345 ;
      RECT MASK 2 30.727 81.463 30.807 81.7345 ;
      RECT MASK 2 31.059 81.463 31.139 81.7345 ;
      RECT MASK 2 37.345 81.463 37.425 81.7345 ;
      RECT MASK 2 37.677 81.463 37.757 81.7345 ;
      RECT MASK 2 43.963 81.463 44.043 81.7345 ;
      RECT MASK 2 44.295 81.463 44.375 81.7345 ;
      RECT MASK 2 50.581 81.463 50.661 81.7345 ;
      RECT MASK 2 50.913 81.463 50.993 81.7345 ;
      RECT MASK 2 57.199 81.463 57.279 81.7345 ;
      RECT MASK 2 57.531 81.463 57.611 81.7345 ;
      RECT MASK 2 63.817 81.463 63.897 81.7345 ;
      RECT MASK 2 64.149 81.463 64.229 81.7345 ;
      RECT MASK 2 70.435 81.463 70.515 81.7345 ;
      RECT MASK 2 70.767 81.463 70.847 81.7345 ;
      RECT MASK 2 77.053 81.463 77.133 81.7345 ;
      RECT MASK 2 77.385 81.463 77.465 81.7345 ;
      RECT MASK 2 83.671 81.463 83.751 81.7345 ;
      RECT MASK 2 84.003 81.463 84.083 81.7345 ;
      RECT MASK 2 90.289 81.463 90.369 81.7345 ;
      RECT MASK 2 90.621 81.463 90.701 81.7345 ;
      RECT MASK 2 96.907 81.463 96.987 81.7345 ;
      RECT MASK 2 97.239 81.463 97.319 81.7345 ;
      RECT MASK 2 103.525 81.463 103.605 81.7345 ;
      RECT MASK 2 103.857 81.463 103.937 81.7345 ;
      RECT MASK 2 111.86 81.467 112.043 81.507 ;
      RECT MASK 2 112.524 81.467 112.707 81.507 ;
      RECT MASK 2 115.613 81.54 128.525 81.58 ;
      RECT MASK 2 111.151 81.651 113.323 81.691 ;
      RECT MASK 2 6.817 81.6515 6.897 81.882 ;
      RECT MASK 2 7.149 81.6515 7.229 81.882 ;
      RECT MASK 2 7.481 81.6515 7.561 81.882 ;
      RECT MASK 2 7.979 81.6515 8.059 81.882 ;
      RECT MASK 2 8.311 81.6515 8.391 81.882 ;
      RECT MASK 2 8.643 81.6515 8.723 81.882 ;
      RECT MASK 2 9.141 81.6515 9.221 81.882 ;
      RECT MASK 2 9.473 81.6515 9.553 81.882 ;
      RECT MASK 2 9.805 81.6515 9.885 81.882 ;
      RECT MASK 2 12.273 81.6515 12.353 81.882 ;
      RECT MASK 2 12.605 81.6515 12.685 81.882 ;
      RECT MASK 2 12.937 81.6515 13.017 81.882 ;
      RECT MASK 2 13.435 81.6515 13.515 81.882 ;
      RECT MASK 2 13.767 81.6515 13.847 81.882 ;
      RECT MASK 2 14.099 81.6515 14.179 81.882 ;
      RECT MASK 2 14.597 81.6515 14.677 81.882 ;
      RECT MASK 2 14.929 81.6515 15.009 81.882 ;
      RECT MASK 2 15.261 81.6515 15.341 81.882 ;
      RECT MASK 2 15.759 81.6515 15.839 81.882 ;
      RECT MASK 2 16.091 81.6515 16.171 81.882 ;
      RECT MASK 2 16.423 81.6515 16.503 81.882 ;
      RECT MASK 2 18.891 81.6515 18.971 81.882 ;
      RECT MASK 2 19.223 81.6515 19.303 81.882 ;
      RECT MASK 2 19.555 81.6515 19.635 81.882 ;
      RECT MASK 2 20.053 81.6515 20.133 81.882 ;
      RECT MASK 2 20.385 81.6515 20.465 81.882 ;
      RECT MASK 2 20.717 81.6515 20.797 81.882 ;
      RECT MASK 2 21.215 81.6515 21.295 81.882 ;
      RECT MASK 2 21.547 81.6515 21.627 81.882 ;
      RECT MASK 2 21.879 81.6515 21.959 81.882 ;
      RECT MASK 2 22.377 81.6515 22.457 81.882 ;
      RECT MASK 2 22.709 81.6515 22.789 81.882 ;
      RECT MASK 2 23.041 81.6515 23.121 81.882 ;
      RECT MASK 2 25.509 81.6515 25.589 81.882 ;
      RECT MASK 2 25.841 81.6515 25.921 81.882 ;
      RECT MASK 2 26.173 81.6515 26.253 81.882 ;
      RECT MASK 2 26.671 81.6515 26.751 81.882 ;
      RECT MASK 2 27.003 81.6515 27.083 81.882 ;
      RECT MASK 2 27.335 81.6515 27.415 81.882 ;
      RECT MASK 2 27.833 81.6515 27.913 81.882 ;
      RECT MASK 2 28.165 81.6515 28.245 81.882 ;
      RECT MASK 2 28.497 81.6515 28.577 81.882 ;
      RECT MASK 2 28.995 81.6515 29.075 81.882 ;
      RECT MASK 2 29.327 81.6515 29.407 81.882 ;
      RECT MASK 2 29.659 81.6515 29.739 81.882 ;
      RECT MASK 2 32.127 81.6515 32.207 81.882 ;
      RECT MASK 2 32.459 81.6515 32.539 81.882 ;
      RECT MASK 2 32.791 81.6515 32.871 81.882 ;
      RECT MASK 2 33.289 81.6515 33.369 81.882 ;
      RECT MASK 2 33.621 81.6515 33.701 81.882 ;
      RECT MASK 2 33.953 81.6515 34.033 81.882 ;
      RECT MASK 2 34.451 81.6515 34.531 81.882 ;
      RECT MASK 2 34.783 81.6515 34.863 81.882 ;
      RECT MASK 2 35.115 81.6515 35.195 81.882 ;
      RECT MASK 2 35.613 81.6515 35.693 81.882 ;
      RECT MASK 2 35.945 81.6515 36.025 81.882 ;
      RECT MASK 2 36.277 81.6515 36.357 81.882 ;
      RECT MASK 2 38.745 81.6515 38.825 81.882 ;
      RECT MASK 2 39.077 81.6515 39.157 81.882 ;
      RECT MASK 2 39.409 81.6515 39.489 81.882 ;
      RECT MASK 2 39.907 81.6515 39.987 81.882 ;
      RECT MASK 2 40.239 81.6515 40.319 81.882 ;
      RECT MASK 2 40.571 81.6515 40.651 81.882 ;
      RECT MASK 2 41.069 81.6515 41.149 81.882 ;
      RECT MASK 2 41.401 81.6515 41.481 81.882 ;
      RECT MASK 2 41.733 81.6515 41.813 81.882 ;
      RECT MASK 2 42.231 81.6515 42.311 81.882 ;
      RECT MASK 2 42.563 81.6515 42.643 81.882 ;
      RECT MASK 2 42.895 81.6515 42.975 81.882 ;
      RECT MASK 2 45.363 81.6515 45.443 81.882 ;
      RECT MASK 2 45.695 81.6515 45.775 81.882 ;
      RECT MASK 2 46.027 81.6515 46.107 81.882 ;
      RECT MASK 2 46.525 81.6515 46.605 81.882 ;
      RECT MASK 2 46.857 81.6515 46.937 81.882 ;
      RECT MASK 2 47.189 81.6515 47.269 81.882 ;
      RECT MASK 2 47.687 81.6515 47.767 81.882 ;
      RECT MASK 2 48.019 81.6515 48.099 81.882 ;
      RECT MASK 2 48.351 81.6515 48.431 81.882 ;
      RECT MASK 2 48.849 81.6515 48.929 81.882 ;
      RECT MASK 2 49.181 81.6515 49.261 81.882 ;
      RECT MASK 2 49.513 81.6515 49.593 81.882 ;
      RECT MASK 2 51.981 81.6515 52.061 81.882 ;
      RECT MASK 2 52.313 81.6515 52.393 81.882 ;
      RECT MASK 2 52.645 81.6515 52.725 81.882 ;
      RECT MASK 2 53.143 81.6515 53.223 81.882 ;
      RECT MASK 2 53.475 81.6515 53.555 81.882 ;
      RECT MASK 2 53.807 81.6515 53.887 81.882 ;
      RECT MASK 2 54.305 81.6515 54.385 81.882 ;
      RECT MASK 2 54.637 81.6515 54.717 81.882 ;
      RECT MASK 2 54.969 81.6515 55.049 81.882 ;
      RECT MASK 2 55.467 81.6515 55.547 81.882 ;
      RECT MASK 2 55.799 81.6515 55.879 81.882 ;
      RECT MASK 2 56.131 81.6515 56.211 81.882 ;
      RECT MASK 2 58.599 81.6515 58.679 81.882 ;
      RECT MASK 2 58.931 81.6515 59.011 81.882 ;
      RECT MASK 2 59.263 81.6515 59.343 81.882 ;
      RECT MASK 2 59.761 81.6515 59.841 81.882 ;
      RECT MASK 2 60.093 81.6515 60.173 81.882 ;
      RECT MASK 2 60.425 81.6515 60.505 81.882 ;
      RECT MASK 2 60.923 81.6515 61.003 81.882 ;
      RECT MASK 2 61.255 81.6515 61.335 81.882 ;
      RECT MASK 2 61.587 81.6515 61.667 81.882 ;
      RECT MASK 2 62.085 81.6515 62.165 81.882 ;
      RECT MASK 2 62.417 81.6515 62.497 81.882 ;
      RECT MASK 2 62.749 81.6515 62.829 81.882 ;
      RECT MASK 2 65.217 81.6515 65.297 81.882 ;
      RECT MASK 2 65.549 81.6515 65.629 81.882 ;
      RECT MASK 2 65.881 81.6515 65.961 81.882 ;
      RECT MASK 2 66.379 81.6515 66.459 81.882 ;
      RECT MASK 2 66.711 81.6515 66.791 81.882 ;
      RECT MASK 2 67.043 81.6515 67.123 81.882 ;
      RECT MASK 2 67.541 81.6515 67.621 81.882 ;
      RECT MASK 2 67.873 81.6515 67.953 81.882 ;
      RECT MASK 2 68.205 81.6515 68.285 81.882 ;
      RECT MASK 2 68.703 81.6515 68.783 81.882 ;
      RECT MASK 2 69.035 81.6515 69.115 81.882 ;
      RECT MASK 2 69.367 81.6515 69.447 81.882 ;
      RECT MASK 2 71.835 81.6515 71.915 81.882 ;
      RECT MASK 2 72.167 81.6515 72.247 81.882 ;
      RECT MASK 2 72.499 81.6515 72.579 81.882 ;
      RECT MASK 2 72.997 81.6515 73.077 81.882 ;
      RECT MASK 2 73.329 81.6515 73.409 81.882 ;
      RECT MASK 2 73.661 81.6515 73.741 81.882 ;
      RECT MASK 2 74.159 81.6515 74.239 81.882 ;
      RECT MASK 2 74.491 81.6515 74.571 81.882 ;
      RECT MASK 2 74.823 81.6515 74.903 81.882 ;
      RECT MASK 2 75.321 81.6515 75.401 81.882 ;
      RECT MASK 2 75.653 81.6515 75.733 81.882 ;
      RECT MASK 2 75.985 81.6515 76.065 81.882 ;
      RECT MASK 2 78.453 81.6515 78.533 81.882 ;
      RECT MASK 2 78.785 81.6515 78.865 81.882 ;
      RECT MASK 2 79.117 81.6515 79.197 81.882 ;
      RECT MASK 2 79.615 81.6515 79.695 81.882 ;
      RECT MASK 2 79.947 81.6515 80.027 81.882 ;
      RECT MASK 2 80.279 81.6515 80.359 81.882 ;
      RECT MASK 2 80.777 81.6515 80.857 81.882 ;
      RECT MASK 2 81.109 81.6515 81.189 81.882 ;
      RECT MASK 2 81.441 81.6515 81.521 81.882 ;
      RECT MASK 2 81.939 81.6515 82.019 81.882 ;
      RECT MASK 2 82.271 81.6515 82.351 81.882 ;
      RECT MASK 2 82.603 81.6515 82.683 81.882 ;
      RECT MASK 2 85.071 81.6515 85.151 81.882 ;
      RECT MASK 2 85.403 81.6515 85.483 81.882 ;
      RECT MASK 2 85.735 81.6515 85.815 81.882 ;
      RECT MASK 2 86.233 81.6515 86.313 81.882 ;
      RECT MASK 2 86.565 81.6515 86.645 81.882 ;
      RECT MASK 2 86.897 81.6515 86.977 81.882 ;
      RECT MASK 2 87.395 81.6515 87.475 81.882 ;
      RECT MASK 2 87.727 81.6515 87.807 81.882 ;
      RECT MASK 2 88.059 81.6515 88.139 81.882 ;
      RECT MASK 2 88.557 81.6515 88.637 81.882 ;
      RECT MASK 2 88.889 81.6515 88.969 81.882 ;
      RECT MASK 2 89.221 81.6515 89.301 81.882 ;
      RECT MASK 2 91.689 81.6515 91.769 81.882 ;
      RECT MASK 2 92.021 81.6515 92.101 81.882 ;
      RECT MASK 2 92.353 81.6515 92.433 81.882 ;
      RECT MASK 2 92.851 81.6515 92.931 81.882 ;
      RECT MASK 2 93.183 81.6515 93.263 81.882 ;
      RECT MASK 2 93.515 81.6515 93.595 81.882 ;
      RECT MASK 2 94.013 81.6515 94.093 81.882 ;
      RECT MASK 2 94.345 81.6515 94.425 81.882 ;
      RECT MASK 2 94.677 81.6515 94.757 81.882 ;
      RECT MASK 2 95.175 81.6515 95.255 81.882 ;
      RECT MASK 2 95.507 81.6515 95.587 81.882 ;
      RECT MASK 2 95.839 81.6515 95.919 81.882 ;
      RECT MASK 2 98.307 81.6515 98.387 81.882 ;
      RECT MASK 2 98.639 81.6515 98.719 81.882 ;
      RECT MASK 2 98.971 81.6515 99.051 81.882 ;
      RECT MASK 2 99.469 81.6515 99.549 81.882 ;
      RECT MASK 2 99.801 81.6515 99.881 81.882 ;
      RECT MASK 2 100.133 81.6515 100.213 81.882 ;
      RECT MASK 2 100.631 81.6515 100.711 81.882 ;
      RECT MASK 2 100.963 81.6515 101.043 81.882 ;
      RECT MASK 2 101.295 81.6515 101.375 81.882 ;
      RECT MASK 2 101.793 81.6515 101.873 81.882 ;
      RECT MASK 2 102.125 81.6515 102.205 81.882 ;
      RECT MASK 2 102.457 81.6515 102.537 81.882 ;
      RECT MASK 2 104.925 81.6515 105.005 81.882 ;
      RECT MASK 2 105.257 81.6515 105.337 81.882 ;
      RECT MASK 2 105.589 81.6515 105.669 81.882 ;
      RECT MASK 2 106.087 81.6515 106.167 81.882 ;
      RECT MASK 2 106.419 81.6515 106.499 81.882 ;
      RECT MASK 2 106.751 81.6515 106.831 81.882 ;
      RECT MASK 2 107.249 81.6515 107.329 81.882 ;
      RECT MASK 2 107.581 81.6515 107.661 81.882 ;
      RECT MASK 2 107.913 81.6515 107.993 81.882 ;
      RECT MASK 2 108.411 81.6515 108.491 81.882 ;
      RECT MASK 2 108.743 81.6515 108.823 81.882 ;
      RECT MASK 2 109.075 81.6515 109.155 81.882 ;
      RECT MASK 2 111.151 81.819 113.323 81.859 ;
      RECT MASK 2 116.599 82.05 116.659 83.1 ;
      RECT MASK 2 116.873 82.05 116.933 83.1 ;
      RECT MASK 2 117.147 82.05 117.207 83.1 ;
      RECT MASK 2 117.421 82.05 117.481 83.1 ;
      RECT MASK 2 117.695 82.05 117.755 83.1 ;
      RECT MASK 2 117.969 82.05 118.029 83.1 ;
      RECT MASK 2 118.243 82.05 118.303 83.1 ;
      RECT MASK 2 118.517 82.05 118.577 83.1 ;
      RECT MASK 2 118.791 82.05 118.851 83.1 ;
      RECT MASK 2 119.065 82.05 119.125 83.1 ;
      RECT MASK 2 119.339 82.05 119.399 83.1 ;
      RECT MASK 2 119.613 82.05 119.673 83.1 ;
      RECT MASK 2 119.887 82.05 119.947 83.1 ;
      RECT MASK 2 120.161 82.05 120.221 83.1 ;
      RECT MASK 2 120.435 82.05 120.495 83.1 ;
      RECT MASK 2 120.709 82.05 120.769 83.1 ;
      RECT MASK 2 120.983 82.05 121.043 83.1 ;
      RECT MASK 2 121.257 82.05 121.317 83.1 ;
      RECT MASK 2 121.531 82.05 121.591 83.1 ;
      RECT MASK 2 121.805 82.05 121.865 83.1 ;
      RECT MASK 2 122.079 82.05 122.139 83.1 ;
      RECT MASK 2 122.353 82.05 122.413 83.1 ;
      RECT MASK 2 122.627 82.05 122.687 83.1 ;
      RECT MASK 2 122.901 82.05 122.961 83.1 ;
      RECT MASK 2 123.175 82.05 123.235 83.1 ;
      RECT MASK 2 123.449 82.05 123.509 83.1 ;
      RECT MASK 2 123.723 82.05 123.783 83.1 ;
      RECT MASK 2 123.997 82.05 124.057 83.1 ;
      RECT MASK 2 124.271 82.05 124.331 83.1 ;
      RECT MASK 2 124.545 82.05 124.605 83.1 ;
      RECT MASK 2 124.819 82.05 124.879 83.1 ;
      RECT MASK 2 125.093 82.05 125.153 83.1 ;
      RECT MASK 2 125.367 82.05 125.427 83.1 ;
      RECT MASK 2 125.641 82.05 125.701 83.1 ;
      RECT MASK 2 125.915 82.05 125.975 83.1 ;
      RECT MASK 2 126.189 82.05 126.249 83.1 ;
      RECT MASK 2 126.463 82.05 126.523 83.1 ;
      RECT MASK 2 126.737 82.05 126.797 83.1 ;
      RECT MASK 2 127.011 82.05 127.071 83.1 ;
      RECT MASK 2 127.285 82.05 127.345 83.1 ;
      RECT MASK 2 127.559 82.05 127.619 83.1 ;
      RECT MASK 2 111.186 82.16 113.288 82.2 ;
      RECT MASK 2 111.186 82.35 113.288 82.39 ;
      RECT MASK 2 6.2775 82.4 109.836 82.44 ;
      RECT MASK 2 6.2775 82.59 109.836 82.63 ;
      RECT MASK 2 2.204 82.68 2.264 83.73 ;
      RECT MASK 2 2.478 82.68 2.538 83.73 ;
      RECT MASK 2 2.752 82.68 2.812 83.73 ;
      RECT MASK 2 3.026 82.68 3.086 83.73 ;
      RECT MASK 2 3.3 82.68 3.36 83.73 ;
      RECT MASK 2 3.574 82.68 3.634 83.73 ;
      RECT MASK 2 3.848 82.68 3.908 83.73 ;
      RECT MASK 2 4.122 82.68 4.182 83.73 ;
      RECT MASK 2 4.396 82.68 4.456 83.73 ;
      RECT MASK 2 6.269 82.961 109.869 83.001 ;
      RECT MASK 2 6.269 83.129 109.869 83.169 ;
      RECT MASK 2 6.978 83.313 7.161 83.353 ;
      RECT MASK 2 7.383 83.313 7.566 83.353 ;
      RECT MASK 2 8.14 83.313 8.323 83.353 ;
      RECT MASK 2 8.545 83.313 8.728 83.353 ;
      RECT MASK 2 9.302 83.313 9.485 83.353 ;
      RECT MASK 2 9.707 83.313 9.89 83.353 ;
      RECT MASK 2 12.434 83.313 12.617 83.353 ;
      RECT MASK 2 12.839 83.313 13.022 83.353 ;
      RECT MASK 2 13.596 83.313 13.779 83.353 ;
      RECT MASK 2 14.001 83.313 14.184 83.353 ;
      RECT MASK 2 14.758 83.313 14.941 83.353 ;
      RECT MASK 2 15.163 83.313 15.346 83.353 ;
      RECT MASK 2 15.92 83.313 16.103 83.353 ;
      RECT MASK 2 16.325 83.313 16.508 83.353 ;
      RECT MASK 2 19.052 83.313 19.235 83.353 ;
      RECT MASK 2 19.457 83.313 19.64 83.353 ;
      RECT MASK 2 20.214 83.313 20.397 83.353 ;
      RECT MASK 2 20.619 83.313 20.802 83.353 ;
      RECT MASK 2 21.376 83.313 21.559 83.353 ;
      RECT MASK 2 21.781 83.313 21.964 83.353 ;
      RECT MASK 2 22.538 83.313 22.721 83.353 ;
      RECT MASK 2 22.943 83.313 23.126 83.353 ;
      RECT MASK 2 25.67 83.313 25.853 83.353 ;
      RECT MASK 2 26.075 83.313 26.258 83.353 ;
      RECT MASK 2 26.832 83.313 27.015 83.353 ;
      RECT MASK 2 27.237 83.313 27.42 83.353 ;
      RECT MASK 2 27.994 83.313 28.177 83.353 ;
      RECT MASK 2 28.399 83.313 28.582 83.353 ;
      RECT MASK 2 29.156 83.313 29.339 83.353 ;
      RECT MASK 2 29.561 83.313 29.744 83.353 ;
      RECT MASK 2 32.288 83.313 32.471 83.353 ;
      RECT MASK 2 32.693 83.313 32.876 83.353 ;
      RECT MASK 2 33.45 83.313 33.633 83.353 ;
      RECT MASK 2 33.855 83.313 34.038 83.353 ;
      RECT MASK 2 34.612 83.313 34.795 83.353 ;
      RECT MASK 2 35.017 83.313 35.2 83.353 ;
      RECT MASK 2 35.774 83.313 35.957 83.353 ;
      RECT MASK 2 36.179 83.313 36.362 83.353 ;
      RECT MASK 2 38.906 83.313 39.089 83.353 ;
      RECT MASK 2 39.311 83.313 39.494 83.353 ;
      RECT MASK 2 40.068 83.313 40.251 83.353 ;
      RECT MASK 2 40.473 83.313 40.656 83.353 ;
      RECT MASK 2 41.23 83.313 41.413 83.353 ;
      RECT MASK 2 41.635 83.313 41.818 83.353 ;
      RECT MASK 2 42.392 83.313 42.575 83.353 ;
      RECT MASK 2 42.797 83.313 42.98 83.353 ;
      RECT MASK 2 45.524 83.313 45.707 83.353 ;
      RECT MASK 2 45.929 83.313 46.112 83.353 ;
      RECT MASK 2 46.686 83.313 46.869 83.353 ;
      RECT MASK 2 47.091 83.313 47.274 83.353 ;
      RECT MASK 2 47.848 83.313 48.031 83.353 ;
      RECT MASK 2 48.253 83.313 48.436 83.353 ;
      RECT MASK 2 49.01 83.313 49.193 83.353 ;
      RECT MASK 2 49.415 83.313 49.598 83.353 ;
      RECT MASK 2 52.142 83.313 52.325 83.353 ;
      RECT MASK 2 52.547 83.313 52.73 83.353 ;
      RECT MASK 2 53.304 83.313 53.487 83.353 ;
      RECT MASK 2 53.709 83.313 53.892 83.353 ;
      RECT MASK 2 54.466 83.313 54.649 83.353 ;
      RECT MASK 2 54.871 83.313 55.054 83.353 ;
      RECT MASK 2 55.628 83.313 55.811 83.353 ;
      RECT MASK 2 56.033 83.313 56.216 83.353 ;
      RECT MASK 2 58.76 83.313 58.943 83.353 ;
      RECT MASK 2 59.165 83.313 59.348 83.353 ;
      RECT MASK 2 59.922 83.313 60.105 83.353 ;
      RECT MASK 2 60.327 83.313 60.51 83.353 ;
      RECT MASK 2 61.084 83.313 61.267 83.353 ;
      RECT MASK 2 61.489 83.313 61.672 83.353 ;
      RECT MASK 2 62.246 83.313 62.429 83.353 ;
      RECT MASK 2 62.651 83.313 62.834 83.353 ;
      RECT MASK 2 65.378 83.313 65.561 83.353 ;
      RECT MASK 2 65.783 83.313 65.966 83.353 ;
      RECT MASK 2 66.54 83.313 66.723 83.353 ;
      RECT MASK 2 66.945 83.313 67.128 83.353 ;
      RECT MASK 2 67.702 83.313 67.885 83.353 ;
      RECT MASK 2 68.107 83.313 68.29 83.353 ;
      RECT MASK 2 68.864 83.313 69.047 83.353 ;
      RECT MASK 2 69.269 83.313 69.452 83.353 ;
      RECT MASK 2 71.996 83.313 72.179 83.353 ;
      RECT MASK 2 72.401 83.313 72.584 83.353 ;
      RECT MASK 2 73.158 83.313 73.341 83.353 ;
      RECT MASK 2 73.563 83.313 73.746 83.353 ;
      RECT MASK 2 74.32 83.313 74.503 83.353 ;
      RECT MASK 2 74.725 83.313 74.908 83.353 ;
      RECT MASK 2 75.482 83.313 75.665 83.353 ;
      RECT MASK 2 75.887 83.313 76.07 83.353 ;
      RECT MASK 2 78.614 83.313 78.797 83.353 ;
      RECT MASK 2 79.019 83.313 79.202 83.353 ;
      RECT MASK 2 79.776 83.313 79.959 83.353 ;
      RECT MASK 2 80.181 83.313 80.364 83.353 ;
      RECT MASK 2 80.938 83.313 81.121 83.353 ;
      RECT MASK 2 81.343 83.313 81.526 83.353 ;
      RECT MASK 2 82.1 83.313 82.283 83.353 ;
      RECT MASK 2 82.505 83.313 82.688 83.353 ;
      RECT MASK 2 85.232 83.313 85.415 83.353 ;
      RECT MASK 2 85.637 83.313 85.82 83.353 ;
      RECT MASK 2 86.394 83.313 86.577 83.353 ;
      RECT MASK 2 86.799 83.313 86.982 83.353 ;
      RECT MASK 2 87.556 83.313 87.739 83.353 ;
      RECT MASK 2 87.961 83.313 88.144 83.353 ;
      RECT MASK 2 88.718 83.313 88.901 83.353 ;
      RECT MASK 2 89.123 83.313 89.306 83.353 ;
      RECT MASK 2 91.85 83.313 92.033 83.353 ;
      RECT MASK 2 92.255 83.313 92.438 83.353 ;
      RECT MASK 2 93.012 83.313 93.195 83.353 ;
      RECT MASK 2 93.417 83.313 93.6 83.353 ;
      RECT MASK 2 94.174 83.313 94.357 83.353 ;
      RECT MASK 2 94.579 83.313 94.762 83.353 ;
      RECT MASK 2 95.336 83.313 95.519 83.353 ;
      RECT MASK 2 95.741 83.313 95.924 83.353 ;
      RECT MASK 2 98.468 83.313 98.651 83.353 ;
      RECT MASK 2 98.873 83.313 99.056 83.353 ;
      RECT MASK 2 99.63 83.313 99.813 83.353 ;
      RECT MASK 2 100.035 83.313 100.218 83.353 ;
      RECT MASK 2 100.792 83.313 100.975 83.353 ;
      RECT MASK 2 101.197 83.313 101.38 83.353 ;
      RECT MASK 2 101.954 83.313 102.137 83.353 ;
      RECT MASK 2 102.359 83.313 102.542 83.353 ;
      RECT MASK 2 105.086 83.313 105.269 83.353 ;
      RECT MASK 2 105.491 83.313 105.674 83.353 ;
      RECT MASK 2 106.248 83.313 106.431 83.353 ;
      RECT MASK 2 106.653 83.313 106.836 83.353 ;
      RECT MASK 2 107.41 83.313 107.593 83.353 ;
      RECT MASK 2 107.815 83.313 107.998 83.353 ;
      RECT MASK 2 108.572 83.313 108.755 83.353 ;
      RECT MASK 2 108.977 83.313 109.16 83.353 ;
      RECT MASK 2 6.269 83.499 6.449 83.539 ;
      RECT MASK 2 10.419 83.499 10.599 83.539 ;
      RECT MASK 2 11.725 83.499 11.905 83.539 ;
      RECT MASK 2 17.037 83.499 17.217 83.539 ;
      RECT MASK 2 18.343 83.499 18.523 83.539 ;
      RECT MASK 2 23.655 83.499 23.835 83.539 ;
      RECT MASK 2 24.961 83.499 25.141 83.539 ;
      RECT MASK 2 30.273 83.499 30.453 83.539 ;
      RECT MASK 2 31.579 83.499 31.759 83.539 ;
      RECT MASK 2 36.891 83.499 37.071 83.539 ;
      RECT MASK 2 38.197 83.499 38.377 83.539 ;
      RECT MASK 2 43.509 83.499 43.689 83.539 ;
      RECT MASK 2 44.815 83.499 44.995 83.539 ;
      RECT MASK 2 50.127 83.499 50.307 83.539 ;
      RECT MASK 2 51.433 83.499 51.613 83.539 ;
      RECT MASK 2 56.745 83.499 56.925 83.539 ;
      RECT MASK 2 58.051 83.499 58.231 83.539 ;
      RECT MASK 2 63.363 83.499 63.543 83.539 ;
      RECT MASK 2 64.669 83.499 64.849 83.539 ;
      RECT MASK 2 69.981 83.499 70.161 83.539 ;
      RECT MASK 2 71.287 83.499 71.467 83.539 ;
      RECT MASK 2 76.599 83.499 76.779 83.539 ;
      RECT MASK 2 77.905 83.499 78.085 83.539 ;
      RECT MASK 2 83.217 83.499 83.397 83.539 ;
      RECT MASK 2 84.523 83.499 84.703 83.539 ;
      RECT MASK 2 89.835 83.499 90.015 83.539 ;
      RECT MASK 2 91.141 83.499 91.321 83.539 ;
      RECT MASK 2 96.453 83.499 96.633 83.539 ;
      RECT MASK 2 97.759 83.499 97.939 83.539 ;
      RECT MASK 2 103.071 83.499 103.251 83.539 ;
      RECT MASK 2 104.377 83.499 104.557 83.539 ;
      RECT MASK 2 109.689 83.499 109.869 83.539 ;
      RECT MASK 2 116.599 83.76 116.659 84.81 ;
      RECT MASK 2 116.873 83.76 116.933 84.81 ;
      RECT MASK 2 117.147 83.76 117.207 84.81 ;
      RECT MASK 2 117.421 83.76 117.481 84.81 ;
      RECT MASK 2 117.695 83.76 117.755 84.81 ;
      RECT MASK 2 117.969 83.76 118.029 84.81 ;
      RECT MASK 2 118.243 83.76 118.303 84.81 ;
      RECT MASK 2 118.517 83.76 118.577 84.81 ;
      RECT MASK 2 118.791 83.76 118.851 84.81 ;
      RECT MASK 2 119.065 83.76 119.125 84.81 ;
      RECT MASK 2 119.339 83.76 119.399 84.81 ;
      RECT MASK 2 119.613 83.76 119.673 84.81 ;
      RECT MASK 2 119.887 83.76 119.947 84.81 ;
      RECT MASK 2 120.161 83.76 120.221 84.81 ;
      RECT MASK 2 120.435 83.76 120.495 84.81 ;
      RECT MASK 2 120.709 83.76 120.769 84.81 ;
      RECT MASK 2 120.983 83.76 121.043 84.81 ;
      RECT MASK 2 121.257 83.76 121.317 84.81 ;
      RECT MASK 2 121.531 83.76 121.591 84.81 ;
      RECT MASK 2 121.805 83.76 121.865 84.81 ;
      RECT MASK 2 122.079 83.76 122.139 84.81 ;
      RECT MASK 2 122.353 83.76 122.413 84.81 ;
      RECT MASK 2 122.627 83.76 122.687 84.81 ;
      RECT MASK 2 122.901 83.76 122.961 84.81 ;
      RECT MASK 2 123.175 83.76 123.235 84.81 ;
      RECT MASK 2 123.449 83.76 123.509 84.81 ;
      RECT MASK 2 123.723 83.76 123.783 84.81 ;
      RECT MASK 2 123.997 83.76 124.057 84.81 ;
      RECT MASK 2 124.271 83.76 124.331 84.81 ;
      RECT MASK 2 124.545 83.76 124.605 84.81 ;
      RECT MASK 2 124.819 83.76 124.879 84.81 ;
      RECT MASK 2 125.093 83.76 125.153 84.81 ;
      RECT MASK 2 125.367 83.76 125.427 84.81 ;
      RECT MASK 2 125.641 83.76 125.701 84.81 ;
      RECT MASK 2 125.915 83.76 125.975 84.81 ;
      RECT MASK 2 126.189 83.76 126.249 84.81 ;
      RECT MASK 2 126.463 83.76 126.523 84.81 ;
      RECT MASK 2 126.737 83.76 126.797 84.81 ;
      RECT MASK 2 127.011 83.76 127.071 84.81 ;
      RECT MASK 2 127.285 83.76 127.345 84.81 ;
      RECT MASK 2 127.559 83.76 127.619 84.81 ;
      RECT MASK 2 6.224 83.945 109.834 83.985 ;
      RECT MASK 2 2.204 84.39 2.264 85.44 ;
      RECT MASK 2 2.478 84.39 2.538 85.44 ;
      RECT MASK 2 2.752 84.39 2.812 85.44 ;
      RECT MASK 2 3.026 84.39 3.086 85.44 ;
      RECT MASK 2 3.3 84.39 3.36 85.44 ;
      RECT MASK 2 3.574 84.39 3.634 85.44 ;
      RECT MASK 2 3.848 84.39 3.908 85.44 ;
      RECT MASK 2 4.122 84.39 4.182 85.44 ;
      RECT MASK 2 4.396 84.39 4.456 85.44 ;
      RECT MASK 2 6.224 84.465 109.834 84.505 ;
      RECT MASK 2 6.269 84.875 6.449 84.915 ;
      RECT MASK 2 10.419 84.875 10.599 84.915 ;
      RECT MASK 2 11.725 84.875 11.905 84.915 ;
      RECT MASK 2 17.037 84.875 17.217 84.915 ;
      RECT MASK 2 18.343 84.875 18.523 84.915 ;
      RECT MASK 2 23.655 84.875 23.835 84.915 ;
      RECT MASK 2 24.961 84.875 25.141 84.915 ;
      RECT MASK 2 30.273 84.875 30.453 84.915 ;
      RECT MASK 2 31.579 84.875 31.759 84.915 ;
      RECT MASK 2 36.891 84.875 37.071 84.915 ;
      RECT MASK 2 38.197 84.875 38.377 84.915 ;
      RECT MASK 2 43.509 84.875 43.689 84.915 ;
      RECT MASK 2 44.815 84.875 44.995 84.915 ;
      RECT MASK 2 50.127 84.875 50.307 84.915 ;
      RECT MASK 2 51.433 84.875 51.613 84.915 ;
      RECT MASK 2 56.745 84.875 56.925 84.915 ;
      RECT MASK 2 58.051 84.875 58.231 84.915 ;
      RECT MASK 2 63.363 84.875 63.543 84.915 ;
      RECT MASK 2 64.669 84.875 64.849 84.915 ;
      RECT MASK 2 69.981 84.875 70.161 84.915 ;
      RECT MASK 2 71.287 84.875 71.467 84.915 ;
      RECT MASK 2 76.599 84.875 76.779 84.915 ;
      RECT MASK 2 77.905 84.875 78.085 84.915 ;
      RECT MASK 2 83.217 84.875 83.397 84.915 ;
      RECT MASK 2 84.523 84.875 84.703 84.915 ;
      RECT MASK 2 89.835 84.875 90.015 84.915 ;
      RECT MASK 2 91.141 84.875 91.321 84.915 ;
      RECT MASK 2 96.453 84.875 96.633 84.915 ;
      RECT MASK 2 97.759 84.875 97.939 84.915 ;
      RECT MASK 2 103.071 84.875 103.251 84.915 ;
      RECT MASK 2 104.377 84.875 104.557 84.915 ;
      RECT MASK 2 109.689 84.875 109.869 84.915 ;
      RECT MASK 2 10.873 84.9185 10.953 85.141 ;
      RECT MASK 2 11.205 84.9185 11.285 85.141 ;
      RECT MASK 2 17.491 84.9185 17.571 85.141 ;
      RECT MASK 2 17.823 84.9185 17.903 85.141 ;
      RECT MASK 2 24.109 84.9185 24.189 85.141 ;
      RECT MASK 2 24.441 84.9185 24.521 85.141 ;
      RECT MASK 2 30.727 84.9185 30.807 85.141 ;
      RECT MASK 2 31.059 84.9185 31.139 85.141 ;
      RECT MASK 2 37.345 84.9185 37.425 85.141 ;
      RECT MASK 2 37.677 84.9185 37.757 85.141 ;
      RECT MASK 2 43.963 84.9185 44.043 85.141 ;
      RECT MASK 2 44.295 84.9185 44.375 85.141 ;
      RECT MASK 2 50.581 84.9185 50.661 85.141 ;
      RECT MASK 2 50.913 84.9185 50.993 85.141 ;
      RECT MASK 2 57.199 84.9185 57.279 85.141 ;
      RECT MASK 2 57.531 84.9185 57.611 85.141 ;
      RECT MASK 2 63.817 84.9185 63.897 85.141 ;
      RECT MASK 2 64.149 84.9185 64.229 85.141 ;
      RECT MASK 2 70.435 84.9185 70.515 85.141 ;
      RECT MASK 2 70.767 84.9185 70.847 85.141 ;
      RECT MASK 2 77.053 84.9185 77.133 85.141 ;
      RECT MASK 2 77.385 84.9185 77.465 85.141 ;
      RECT MASK 2 83.671 84.9185 83.751 85.141 ;
      RECT MASK 2 84.003 84.9185 84.083 85.141 ;
      RECT MASK 2 90.289 84.9185 90.369 85.141 ;
      RECT MASK 2 90.621 84.9185 90.701 85.141 ;
      RECT MASK 2 96.907 84.9185 96.987 85.141 ;
      RECT MASK 2 97.239 84.9185 97.319 85.141 ;
      RECT MASK 2 103.525 84.9185 103.605 85.141 ;
      RECT MASK 2 103.857 84.9185 103.937 85.141 ;
      RECT MASK 2 6.978 85.097 7.161 85.137 ;
      RECT MASK 2 7.383 85.097 7.566 85.137 ;
      RECT MASK 2 8.14 85.097 8.323 85.137 ;
      RECT MASK 2 8.545 85.097 8.728 85.137 ;
      RECT MASK 2 9.302 85.097 9.485 85.137 ;
      RECT MASK 2 9.707 85.097 9.89 85.137 ;
      RECT MASK 2 12.434 85.097 12.617 85.137 ;
      RECT MASK 2 12.839 85.097 13.022 85.137 ;
      RECT MASK 2 13.596 85.097 13.779 85.137 ;
      RECT MASK 2 14.001 85.097 14.184 85.137 ;
      RECT MASK 2 14.758 85.097 14.941 85.137 ;
      RECT MASK 2 15.163 85.097 15.346 85.137 ;
      RECT MASK 2 15.92 85.097 16.103 85.137 ;
      RECT MASK 2 16.325 85.097 16.508 85.137 ;
      RECT MASK 2 19.052 85.097 19.235 85.137 ;
      RECT MASK 2 19.457 85.097 19.64 85.137 ;
      RECT MASK 2 20.214 85.097 20.397 85.137 ;
      RECT MASK 2 20.619 85.097 20.802 85.137 ;
      RECT MASK 2 21.376 85.097 21.559 85.137 ;
      RECT MASK 2 21.781 85.097 21.964 85.137 ;
      RECT MASK 2 22.538 85.097 22.721 85.137 ;
      RECT MASK 2 22.943 85.097 23.126 85.137 ;
      RECT MASK 2 25.67 85.097 25.853 85.137 ;
      RECT MASK 2 26.075 85.097 26.258 85.137 ;
      RECT MASK 2 26.832 85.097 27.015 85.137 ;
      RECT MASK 2 27.237 85.097 27.42 85.137 ;
      RECT MASK 2 27.994 85.097 28.177 85.137 ;
      RECT MASK 2 28.399 85.097 28.582 85.137 ;
      RECT MASK 2 29.156 85.097 29.339 85.137 ;
      RECT MASK 2 29.561 85.097 29.744 85.137 ;
      RECT MASK 2 32.288 85.097 32.471 85.137 ;
      RECT MASK 2 32.693 85.097 32.876 85.137 ;
      RECT MASK 2 33.45 85.097 33.633 85.137 ;
      RECT MASK 2 33.855 85.097 34.038 85.137 ;
      RECT MASK 2 34.612 85.097 34.795 85.137 ;
      RECT MASK 2 35.017 85.097 35.2 85.137 ;
      RECT MASK 2 35.774 85.097 35.957 85.137 ;
      RECT MASK 2 36.179 85.097 36.362 85.137 ;
      RECT MASK 2 38.906 85.097 39.089 85.137 ;
      RECT MASK 2 39.311 85.097 39.494 85.137 ;
      RECT MASK 2 40.068 85.097 40.251 85.137 ;
      RECT MASK 2 40.473 85.097 40.656 85.137 ;
      RECT MASK 2 41.23 85.097 41.413 85.137 ;
      RECT MASK 2 41.635 85.097 41.818 85.137 ;
      RECT MASK 2 42.392 85.097 42.575 85.137 ;
      RECT MASK 2 42.797 85.097 42.98 85.137 ;
      RECT MASK 2 45.524 85.097 45.707 85.137 ;
      RECT MASK 2 45.929 85.097 46.112 85.137 ;
      RECT MASK 2 46.686 85.097 46.869 85.137 ;
      RECT MASK 2 47.091 85.097 47.274 85.137 ;
      RECT MASK 2 47.848 85.097 48.031 85.137 ;
      RECT MASK 2 48.253 85.097 48.436 85.137 ;
      RECT MASK 2 49.01 85.097 49.193 85.137 ;
      RECT MASK 2 49.415 85.097 49.598 85.137 ;
      RECT MASK 2 52.142 85.097 52.325 85.137 ;
      RECT MASK 2 52.547 85.097 52.73 85.137 ;
      RECT MASK 2 53.304 85.097 53.487 85.137 ;
      RECT MASK 2 53.709 85.097 53.892 85.137 ;
      RECT MASK 2 54.466 85.097 54.649 85.137 ;
      RECT MASK 2 54.871 85.097 55.054 85.137 ;
      RECT MASK 2 55.628 85.097 55.811 85.137 ;
      RECT MASK 2 56.033 85.097 56.216 85.137 ;
      RECT MASK 2 58.76 85.097 58.943 85.137 ;
      RECT MASK 2 59.165 85.097 59.348 85.137 ;
      RECT MASK 2 59.922 85.097 60.105 85.137 ;
      RECT MASK 2 60.327 85.097 60.51 85.137 ;
      RECT MASK 2 61.084 85.097 61.267 85.137 ;
      RECT MASK 2 61.489 85.097 61.672 85.137 ;
      RECT MASK 2 62.246 85.097 62.429 85.137 ;
      RECT MASK 2 62.651 85.097 62.834 85.137 ;
      RECT MASK 2 65.378 85.097 65.561 85.137 ;
      RECT MASK 2 65.783 85.097 65.966 85.137 ;
      RECT MASK 2 66.54 85.097 66.723 85.137 ;
      RECT MASK 2 66.945 85.097 67.128 85.137 ;
      RECT MASK 2 67.702 85.097 67.885 85.137 ;
      RECT MASK 2 68.107 85.097 68.29 85.137 ;
      RECT MASK 2 68.864 85.097 69.047 85.137 ;
      RECT MASK 2 69.269 85.097 69.452 85.137 ;
      RECT MASK 2 71.996 85.097 72.179 85.137 ;
      RECT MASK 2 72.401 85.097 72.584 85.137 ;
      RECT MASK 2 73.158 85.097 73.341 85.137 ;
      RECT MASK 2 73.563 85.097 73.746 85.137 ;
      RECT MASK 2 74.32 85.097 74.503 85.137 ;
      RECT MASK 2 74.725 85.097 74.908 85.137 ;
      RECT MASK 2 75.482 85.097 75.665 85.137 ;
      RECT MASK 2 75.887 85.097 76.07 85.137 ;
      RECT MASK 2 78.614 85.097 78.797 85.137 ;
      RECT MASK 2 79.019 85.097 79.202 85.137 ;
      RECT MASK 2 79.776 85.097 79.959 85.137 ;
      RECT MASK 2 80.181 85.097 80.364 85.137 ;
      RECT MASK 2 80.938 85.097 81.121 85.137 ;
      RECT MASK 2 81.343 85.097 81.526 85.137 ;
      RECT MASK 2 82.1 85.097 82.283 85.137 ;
      RECT MASK 2 82.505 85.097 82.688 85.137 ;
      RECT MASK 2 85.232 85.097 85.415 85.137 ;
      RECT MASK 2 85.637 85.097 85.82 85.137 ;
      RECT MASK 2 86.394 85.097 86.577 85.137 ;
      RECT MASK 2 86.799 85.097 86.982 85.137 ;
      RECT MASK 2 87.556 85.097 87.739 85.137 ;
      RECT MASK 2 87.961 85.097 88.144 85.137 ;
      RECT MASK 2 88.718 85.097 88.901 85.137 ;
      RECT MASK 2 89.123 85.097 89.306 85.137 ;
      RECT MASK 2 91.85 85.097 92.033 85.137 ;
      RECT MASK 2 92.255 85.097 92.438 85.137 ;
      RECT MASK 2 93.012 85.097 93.195 85.137 ;
      RECT MASK 2 93.417 85.097 93.6 85.137 ;
      RECT MASK 2 94.174 85.097 94.357 85.137 ;
      RECT MASK 2 94.579 85.097 94.762 85.137 ;
      RECT MASK 2 95.336 85.097 95.519 85.137 ;
      RECT MASK 2 95.741 85.097 95.924 85.137 ;
      RECT MASK 2 98.468 85.097 98.651 85.137 ;
      RECT MASK 2 98.873 85.097 99.056 85.137 ;
      RECT MASK 2 99.63 85.097 99.813 85.137 ;
      RECT MASK 2 100.035 85.097 100.218 85.137 ;
      RECT MASK 2 100.792 85.097 100.975 85.137 ;
      RECT MASK 2 101.197 85.097 101.38 85.137 ;
      RECT MASK 2 101.954 85.097 102.137 85.137 ;
      RECT MASK 2 102.359 85.097 102.542 85.137 ;
      RECT MASK 2 105.086 85.097 105.269 85.137 ;
      RECT MASK 2 105.491 85.097 105.674 85.137 ;
      RECT MASK 2 106.248 85.097 106.431 85.137 ;
      RECT MASK 2 106.653 85.097 106.836 85.137 ;
      RECT MASK 2 107.41 85.097 107.593 85.137 ;
      RECT MASK 2 107.815 85.097 107.998 85.137 ;
      RECT MASK 2 108.572 85.097 108.755 85.137 ;
      RECT MASK 2 108.977 85.097 109.16 85.137 ;
      RECT MASK 2 6.224 85.281 109.898 85.321 ;
      RECT MASK 2 6.224 85.449 109.898 85.489 ;
      RECT MASK 2 116.599 85.47 116.659 86.52 ;
      RECT MASK 2 116.873 85.47 116.933 86.52 ;
      RECT MASK 2 117.147 85.47 117.207 86.52 ;
      RECT MASK 2 117.421 85.47 117.481 86.52 ;
      RECT MASK 2 117.695 85.47 117.755 86.52 ;
      RECT MASK 2 117.969 85.47 118.029 86.52 ;
      RECT MASK 2 118.243 85.47 118.303 86.52 ;
      RECT MASK 2 118.517 85.47 118.577 86.52 ;
      RECT MASK 2 118.791 85.47 118.851 86.52 ;
      RECT MASK 2 119.065 85.47 119.125 86.52 ;
      RECT MASK 2 119.339 85.47 119.399 86.52 ;
      RECT MASK 2 119.613 85.47 119.673 86.52 ;
      RECT MASK 2 119.887 85.47 119.947 86.52 ;
      RECT MASK 2 120.161 85.47 120.221 86.52 ;
      RECT MASK 2 120.435 85.47 120.495 86.52 ;
      RECT MASK 2 120.709 85.47 120.769 86.52 ;
      RECT MASK 2 120.983 85.47 121.043 86.52 ;
      RECT MASK 2 121.257 85.47 121.317 86.52 ;
      RECT MASK 2 121.531 85.47 121.591 86.52 ;
      RECT MASK 2 121.805 85.47 121.865 86.52 ;
      RECT MASK 2 122.079 85.47 122.139 86.52 ;
      RECT MASK 2 122.353 85.47 122.413 86.52 ;
      RECT MASK 2 122.627 85.47 122.687 86.52 ;
      RECT MASK 2 122.901 85.47 122.961 86.52 ;
      RECT MASK 2 123.175 85.47 123.235 86.52 ;
      RECT MASK 2 123.449 85.47 123.509 86.52 ;
      RECT MASK 2 123.723 85.47 123.783 86.52 ;
      RECT MASK 2 123.997 85.47 124.057 86.52 ;
      RECT MASK 2 124.271 85.47 124.331 86.52 ;
      RECT MASK 2 124.545 85.47 124.605 86.52 ;
      RECT MASK 2 124.819 85.47 124.879 86.52 ;
      RECT MASK 2 125.093 85.47 125.153 86.52 ;
      RECT MASK 2 125.367 85.47 125.427 86.52 ;
      RECT MASK 2 125.641 85.47 125.701 86.52 ;
      RECT MASK 2 125.915 85.47 125.975 86.52 ;
      RECT MASK 2 126.189 85.47 126.249 86.52 ;
      RECT MASK 2 126.463 85.47 126.523 86.52 ;
      RECT MASK 2 126.737 85.47 126.797 86.52 ;
      RECT MASK 2 127.011 85.47 127.071 86.52 ;
      RECT MASK 2 127.285 85.47 127.345 86.52 ;
      RECT MASK 2 127.559 85.47 127.619 86.52 ;
      RECT MASK 2 6.224 85.79 109.826 85.83 ;
      RECT MASK 2 6.224 85.98 109.826 86.02 ;
      RECT MASK 2 2.204 86.1 2.264 87.15 ;
      RECT MASK 2 2.478 86.1 2.538 87.15 ;
      RECT MASK 2 2.752 86.1 2.812 87.15 ;
      RECT MASK 2 3.026 86.1 3.086 87.15 ;
      RECT MASK 2 3.3 86.1 3.36 87.15 ;
      RECT MASK 2 3.574 86.1 3.634 87.15 ;
      RECT MASK 2 3.848 86.1 3.908 87.15 ;
      RECT MASK 2 4.122 86.1 4.182 87.15 ;
      RECT MASK 2 4.396 86.1 4.456 87.15 ;
      RECT MASK 2 71.997 86.259 103.585 86.319 ;
      RECT MASK 2 69.797 86.27 71.728 86.31 ;
      RECT MASK 2 103.854 86.27 105.785 86.31 ;
      RECT MASK 2 33.407 86.36 35.338 86.4 ;
      RECT MASK 2 67.472 86.36 69.229 86.4 ;
      RECT MASK 2 69.797 86.46 71.728 86.5 ;
      RECT MASK 2 103.854 86.46 105.785 86.5 ;
      RECT MASK 2 33.407 86.55 35.338 86.59 ;
      RECT MASK 2 67.472 86.55 69.229 86.59 ;
      RECT MASK 2 70.129 86.72 71.728 86.76 ;
      RECT MASK 2 103.854 86.72 105.453 86.76 ;
      RECT MASK 2 33.739 86.81 35.338 86.85 ;
      RECT MASK 2 67.472 86.81 68.897 86.85 ;
      RECT MASK 2 115.613 86.81 128.525 86.85 ;
      RECT MASK 2 70.129 86.91 71.728 86.95 ;
      RECT MASK 2 103.854 86.91 105.453 86.95 ;
      RECT MASK 2 33.739 87 35.338 87.04 ;
      RECT MASK 2 67.472 87 68.897 87.04 ;
      RECT MASK 2 115.613 87 128.525 87.04 ;
      RECT MASK 2 36.326 87.021 66.476 87.081 ;
      RECT MASK 2 72.716 87.021 102.866 87.081 ;
      RECT MASK 2 25.67 87.101 30.62 87.161 ;
      RECT MASK 2 5.984 87.23 12.811 87.27 ;
      RECT MASK 2 13.208 87.23 17.19 87.27 ;
      RECT MASK 2 17.592 87.23 22.239 87.27 ;
      RECT MASK 2 107.479 87.26 128.525 87.3 ;
      RECT MASK 2 36.326 87.273 66.476 87.333 ;
      RECT MASK 2 72.716 87.273 102.866 87.333 ;
      RECT MASK 2 25.67 87.363 30.62 87.423 ;
      RECT MASK 2 34.36 87.38 35.134 87.42 ;
      RECT MASK 2 67.676 87.38 68.276 87.42 ;
      RECT MASK 2 70.75 87.38 71.524 87.42 ;
      RECT MASK 2 104.058 87.38 104.832 87.42 ;
      RECT MASK 2 22.444 87.41 24.198 87.45 ;
      RECT MASK 2 5.984 87.42 12.811 87.46 ;
      RECT MASK 2 13.208 87.42 17.19 87.46 ;
      RECT MASK 2 17.592 87.42 22.239 87.46 ;
      RECT MASK 2 107.479 87.45 128.525 87.49 ;
      RECT MASK 2 36.326 87.499 66.476 87.559 ;
      RECT MASK 2 72.716 87.499 102.866 87.559 ;
      RECT MASK 2 34.36 87.54 35.134 87.58 ;
      RECT MASK 2 67.676 87.54 68.276 87.58 ;
      RECT MASK 2 70.75 87.54 71.524 87.58 ;
      RECT MASK 2 104.058 87.54 104.832 87.58 ;
      RECT MASK 2 71.997 87.56 72.269 87.62 ;
      RECT MASK 2 103.313 87.56 103.585 87.62 ;
      RECT MASK 2 22.444 87.57 24.198 87.61 ;
      RECT MASK 2 8.7735 87.68 12.2035 87.72 ;
      RECT MASK 2 13.8215 87.68 16.5875 87.72 ;
      RECT MASK 2 18.2055 87.68 21.6355 87.72 ;
      RECT MASK 2 5.92 87.761 7.154 87.801 ;
      RECT MASK 2 2.204 87.81 2.264 88.86 ;
      RECT MASK 2 2.478 87.81 2.538 88.86 ;
      RECT MASK 2 2.752 87.81 2.812 88.86 ;
      RECT MASK 2 3.026 87.81 3.086 88.86 ;
      RECT MASK 2 3.3 87.81 3.36 88.86 ;
      RECT MASK 2 3.574 87.81 3.634 88.86 ;
      RECT MASK 2 3.848 87.81 3.908 88.86 ;
      RECT MASK 2 4.122 87.81 4.182 88.86 ;
      RECT MASK 2 4.396 87.81 4.456 88.86 ;
      RECT MASK 2 22.444 87.83 24.198 87.87 ;
      RECT MASK 2 8.7735 87.87 12.2035 87.91 ;
      RECT MASK 2 13.8215 87.87 16.5875 87.91 ;
      RECT MASK 2 18.2055 87.87 21.6355 87.91 ;
      RECT MASK 2 34.36 87.914 35.134 87.994 ;
      RECT MASK 2 67.676 87.914 68.276 87.994 ;
      RECT MASK 2 70.75 87.914 71.524 87.994 ;
      RECT MASK 2 104.058 87.914 104.832 87.994 ;
      RECT MASK 2 36.326 87.921 36.778 87.981 ;
      RECT MASK 2 37.048 87.921 65.754 87.981 ;
      RECT MASK 2 66.024 87.921 66.476 87.981 ;
      RECT MASK 2 72.716 87.921 73.168 87.981 ;
      RECT MASK 2 73.438 87.921 102.144 87.981 ;
      RECT MASK 2 102.414 87.921 102.866 87.981 ;
      RECT MASK 2 5.92 87.929 7.154 87.969 ;
      RECT MASK 2 108.379 87.93 108.439 88.98 ;
      RECT MASK 2 108.653 87.93 108.713 88.98 ;
      RECT MASK 2 108.927 87.93 108.987 88.98 ;
      RECT MASK 2 109.201 87.93 109.261 88.98 ;
      RECT MASK 2 109.475 87.93 109.535 88.98 ;
      RECT MASK 2 109.749 87.93 109.809 88.98 ;
      RECT MASK 2 110.023 87.93 110.083 88.98 ;
      RECT MASK 2 110.297 87.93 110.357 88.98 ;
      RECT MASK 2 110.571 87.93 110.631 88.98 ;
      RECT MASK 2 110.845 87.93 110.905 88.98 ;
      RECT MASK 2 111.119 87.93 111.179 88.98 ;
      RECT MASK 2 111.393 87.93 111.453 88.98 ;
      RECT MASK 2 111.667 87.93 111.727 88.98 ;
      RECT MASK 2 111.941 87.93 112.001 88.98 ;
      RECT MASK 2 112.215 87.93 112.275 88.98 ;
      RECT MASK 2 112.489 87.93 112.549 88.98 ;
      RECT MASK 2 112.763 87.93 112.823 88.98 ;
      RECT MASK 2 113.037 87.93 113.097 88.98 ;
      RECT MASK 2 113.311 87.93 113.371 88.98 ;
      RECT MASK 2 113.585 87.93 113.645 88.98 ;
      RECT MASK 2 113.859 87.93 113.919 88.98 ;
      RECT MASK 2 114.133 87.93 114.193 88.98 ;
      RECT MASK 2 114.407 87.93 114.467 88.98 ;
      RECT MASK 2 114.681 87.93 114.741 88.98 ;
      RECT MASK 2 114.955 87.93 115.015 88.98 ;
      RECT MASK 2 115.229 87.93 115.289 88.98 ;
      RECT MASK 2 115.503 87.93 115.563 88.98 ;
      RECT MASK 2 115.777 87.93 115.837 88.98 ;
      RECT MASK 2 116.051 87.93 116.111 88.98 ;
      RECT MASK 2 116.325 87.93 116.385 88.98 ;
      RECT MASK 2 116.599 87.93 116.659 88.98 ;
      RECT MASK 2 116.873 87.93 116.933 88.98 ;
      RECT MASK 2 117.147 87.93 117.207 88.98 ;
      RECT MASK 2 117.421 87.93 117.481 88.98 ;
      RECT MASK 2 117.695 87.93 117.755 88.98 ;
      RECT MASK 2 117.969 87.93 118.029 88.98 ;
      RECT MASK 2 118.243 87.93 118.303 88.98 ;
      RECT MASK 2 118.517 87.93 118.577 88.98 ;
      RECT MASK 2 118.791 87.93 118.851 88.98 ;
      RECT MASK 2 119.065 87.93 119.125 88.98 ;
      RECT MASK 2 119.339 87.93 119.399 88.98 ;
      RECT MASK 2 119.613 87.93 119.673 88.98 ;
      RECT MASK 2 119.887 87.93 119.947 88.98 ;
      RECT MASK 2 120.161 87.93 120.221 88.98 ;
      RECT MASK 2 120.435 87.93 120.495 88.98 ;
      RECT MASK 2 120.709 87.93 120.769 88.98 ;
      RECT MASK 2 120.983 87.93 121.043 88.98 ;
      RECT MASK 2 121.257 87.93 121.317 88.98 ;
      RECT MASK 2 121.531 87.93 121.591 88.98 ;
      RECT MASK 2 121.805 87.93 121.865 88.98 ;
      RECT MASK 2 122.079 87.93 122.139 88.98 ;
      RECT MASK 2 122.353 87.93 122.413 88.98 ;
      RECT MASK 2 122.627 87.93 122.687 88.98 ;
      RECT MASK 2 122.901 87.93 122.961 88.98 ;
      RECT MASK 2 123.175 87.93 123.235 88.98 ;
      RECT MASK 2 123.449 87.93 123.509 88.98 ;
      RECT MASK 2 123.723 87.93 123.783 88.98 ;
      RECT MASK 2 123.997 87.93 124.057 88.98 ;
      RECT MASK 2 124.271 87.93 124.331 88.98 ;
      RECT MASK 2 124.545 87.93 124.605 88.98 ;
      RECT MASK 2 124.819 87.93 124.879 88.98 ;
      RECT MASK 2 125.093 87.93 125.153 88.98 ;
      RECT MASK 2 125.367 87.93 125.427 88.98 ;
      RECT MASK 2 125.641 87.93 125.701 88.98 ;
      RECT MASK 2 125.915 87.93 125.975 88.98 ;
      RECT MASK 2 126.189 87.93 126.249 88.98 ;
      RECT MASK 2 126.463 87.93 126.523 88.98 ;
      RECT MASK 2 126.737 87.93 126.797 88.98 ;
      RECT MASK 2 127.011 87.93 127.071 88.98 ;
      RECT MASK 2 127.285 87.93 127.345 88.98 ;
      RECT MASK 2 127.559 87.93 127.619 88.98 ;
      RECT MASK 2 25.67 87.957 25.938 88.017 ;
      RECT MASK 2 26.212 87.957 30.078 88.017 ;
      RECT MASK 2 30.352 87.957 30.62 88.017 ;
      RECT MASK 2 22.444 87.99 24.198 88.03 ;
      RECT MASK 2 6.492 88.113 6.675 88.153 ;
      RECT MASK 2 9.1055 88.13 11.8715 88.17 ;
      RECT MASK 2 14.1405 88.13 16.2815 88.17 ;
      RECT MASK 2 18.5375 88.13 21.3035 88.17 ;
      RECT MASK 2 36.326 88.173 36.778 88.233 ;
      RECT MASK 2 37.048 88.173 65.754 88.233 ;
      RECT MASK 2 66.024 88.173 66.476 88.233 ;
      RECT MASK 2 72.716 88.173 73.168 88.233 ;
      RECT MASK 2 73.438 88.173 102.144 88.233 ;
      RECT MASK 2 102.414 88.173 102.866 88.233 ;
      RECT MASK 2 34.36 88.226 35.134 88.306 ;
      RECT MASK 2 67.676 88.226 68.276 88.306 ;
      RECT MASK 2 70.75 88.226 71.524 88.306 ;
      RECT MASK 2 104.058 88.226 104.832 88.306 ;
      RECT MASK 2 22.444 88.25 24.198 88.29 ;
      RECT MASK 2 9.1055 88.32 11.8715 88.36 ;
      RECT MASK 2 14.1405 88.32 16.2815 88.36 ;
      RECT MASK 2 18.5375 88.32 21.3035 88.36 ;
      RECT MASK 2 5.949 88.335 6.129 88.375 ;
      RECT MASK 2 6.945 88.335 7.125 88.375 ;
      RECT MASK 2 36.323 88.399 36.787 88.459 ;
      RECT MASK 2 37.047 88.399 65.755 88.459 ;
      RECT MASK 2 66.015 88.399 66.479 88.459 ;
      RECT MASK 2 72.713 88.399 73.177 88.459 ;
      RECT MASK 2 73.437 88.399 102.145 88.459 ;
      RECT MASK 2 102.405 88.399 102.869 88.459 ;
      RECT MASK 2 22.444 88.41 24.198 88.45 ;
      RECT MASK 2 25.67 88.541 30.62 88.601 ;
      RECT MASK 2 22.444 88.67 24.198 88.71 ;
      RECT MASK 2 9.2965 88.688 9.3565 88.912 ;
      RECT MASK 2 9.6285 88.688 9.6885 88.912 ;
      RECT MASK 2 9.9605 88.688 10.0205 88.912 ;
      RECT MASK 2 10.2925 88.688 10.3525 88.912 ;
      RECT MASK 2 10.6245 88.688 10.6845 88.912 ;
      RECT MASK 2 10.9565 88.688 11.0165 88.912 ;
      RECT MASK 2 11.2885 88.688 11.3485 88.912 ;
      RECT MASK 2 11.6205 88.688 11.6805 88.912 ;
      RECT MASK 2 14.3445 88.688 14.4045 88.912 ;
      RECT MASK 2 14.6765 88.688 14.7365 88.912 ;
      RECT MASK 2 15.0085 88.688 15.0685 88.912 ;
      RECT MASK 2 15.3405 88.688 15.4005 88.912 ;
      RECT MASK 2 15.6725 88.688 15.7325 88.912 ;
      RECT MASK 2 16.0045 88.688 16.0645 88.912 ;
      RECT MASK 2 18.5625 88.688 18.6225 88.912 ;
      RECT MASK 2 18.8945 88.688 18.9545 88.912 ;
      RECT MASK 2 19.2265 88.688 19.2865 88.912 ;
      RECT MASK 2 19.5585 88.688 19.6185 88.912 ;
      RECT MASK 2 19.8905 88.688 19.9505 88.912 ;
      RECT MASK 2 20.2225 88.688 20.2825 88.912 ;
      RECT MASK 2 20.5545 88.688 20.6145 88.912 ;
      RECT MASK 2 20.8865 88.688 20.9465 88.912 ;
      RECT MASK 2 21.2185 88.688 21.2785 88.912 ;
      RECT MASK 2 5.984 88.745 7.09 88.785 ;
      RECT MASK 2 34.36 88.754 35.134 88.834 ;
      RECT MASK 2 67.676 88.754 68.276 88.834 ;
      RECT MASK 2 70.75 88.754 71.524 88.834 ;
      RECT MASK 2 104.058 88.754 104.832 88.834 ;
      RECT MASK 2 25.67 88.803 30.62 88.863 ;
      RECT MASK 2 36.326 88.821 66.476 88.881 ;
      RECT MASK 2 72.716 88.821 102.866 88.881 ;
      RECT MASK 2 22.444 88.83 24.198 88.87 ;
      RECT MASK 2 34.36 89.066 35.134 89.146 ;
      RECT MASK 2 67.676 89.066 68.276 89.146 ;
      RECT MASK 2 70.75 89.066 71.524 89.146 ;
      RECT MASK 2 104.058 89.066 104.832 89.146 ;
      RECT MASK 2 8.9875 89.07 9.4995 89.11 ;
      RECT MASK 2 11.4775 89.07 11.9545 89.11 ;
      RECT MASK 2 14.0355 89.07 14.5475 89.11 ;
      RECT MASK 2 15.8615 89.07 16.3385 89.11 ;
      RECT MASK 2 18.4195 89.07 18.9315 89.11 ;
      RECT MASK 2 20.9095 89.07 21.3865 89.11 ;
      RECT MASK 2 36.326 89.073 66.476 89.133 ;
      RECT MASK 2 72.716 89.073 102.866 89.133 ;
      RECT MASK 2 22.444 89.09 24.198 89.13 ;
      RECT MASK 2 22.444 89.25 24.198 89.29 ;
      RECT MASK 2 5.984 89.265 7.09 89.305 ;
      RECT MASK 2 8.9875 89.27 9.4995 89.31 ;
      RECT MASK 2 11.4775 89.27 11.9545 89.31 ;
      RECT MASK 2 14.0355 89.27 14.5475 89.31 ;
      RECT MASK 2 15.8615 89.27 16.3385 89.31 ;
      RECT MASK 2 18.4195 89.27 18.9315 89.31 ;
      RECT MASK 2 20.9095 89.27 21.3865 89.31 ;
      RECT MASK 2 36.326 89.299 66.476 89.359 ;
      RECT MASK 2 72.716 89.299 102.866 89.359 ;
      RECT MASK 2 71.997 89.36 72.269 89.42 ;
      RECT MASK 2 103.313 89.36 103.585 89.42 ;
      RECT MASK 2 108.379 89.43 108.439 90.48 ;
      RECT MASK 2 108.653 89.43 108.713 90.48 ;
      RECT MASK 2 108.927 89.43 108.987 90.48 ;
      RECT MASK 2 109.201 89.43 109.261 90.48 ;
      RECT MASK 2 109.475 89.43 109.535 90.48 ;
      RECT MASK 2 109.749 89.43 109.809 90.48 ;
      RECT MASK 2 110.023 89.43 110.083 90.48 ;
      RECT MASK 2 110.297 89.43 110.357 90.48 ;
      RECT MASK 2 110.571 89.43 110.631 90.48 ;
      RECT MASK 2 110.845 89.43 110.905 90.48 ;
      RECT MASK 2 111.119 89.43 111.179 90.48 ;
      RECT MASK 2 111.393 89.43 111.453 90.48 ;
      RECT MASK 2 111.667 89.43 111.727 90.48 ;
      RECT MASK 2 111.941 89.43 112.001 90.48 ;
      RECT MASK 2 112.215 89.43 112.275 90.48 ;
      RECT MASK 2 112.489 89.43 112.549 90.48 ;
      RECT MASK 2 112.763 89.43 112.823 90.48 ;
      RECT MASK 2 113.037 89.43 113.097 90.48 ;
      RECT MASK 2 113.311 89.43 113.371 90.48 ;
      RECT MASK 2 113.585 89.43 113.645 90.48 ;
      RECT MASK 2 113.859 89.43 113.919 90.48 ;
      RECT MASK 2 114.133 89.43 114.193 90.48 ;
      RECT MASK 2 114.407 89.43 114.467 90.48 ;
      RECT MASK 2 114.681 89.43 114.741 90.48 ;
      RECT MASK 2 114.955 89.43 115.015 90.48 ;
      RECT MASK 2 115.229 89.43 115.289 90.48 ;
      RECT MASK 2 115.503 89.43 115.563 90.48 ;
      RECT MASK 2 115.777 89.43 115.837 90.48 ;
      RECT MASK 2 116.051 89.43 116.111 90.48 ;
      RECT MASK 2 116.325 89.43 116.385 90.48 ;
      RECT MASK 2 116.599 89.43 116.659 90.48 ;
      RECT MASK 2 116.873 89.43 116.933 90.48 ;
      RECT MASK 2 117.147 89.43 117.207 90.48 ;
      RECT MASK 2 117.421 89.43 117.481 90.48 ;
      RECT MASK 2 117.695 89.43 117.755 90.48 ;
      RECT MASK 2 117.969 89.43 118.029 90.48 ;
      RECT MASK 2 118.243 89.43 118.303 90.48 ;
      RECT MASK 2 118.517 89.43 118.577 90.48 ;
      RECT MASK 2 118.791 89.43 118.851 90.48 ;
      RECT MASK 2 119.065 89.43 119.125 90.48 ;
      RECT MASK 2 119.339 89.43 119.399 90.48 ;
      RECT MASK 2 119.613 89.43 119.673 90.48 ;
      RECT MASK 2 119.887 89.43 119.947 90.48 ;
      RECT MASK 2 120.161 89.43 120.221 90.48 ;
      RECT MASK 2 120.435 89.43 120.495 90.48 ;
      RECT MASK 2 120.709 89.43 120.769 90.48 ;
      RECT MASK 2 120.983 89.43 121.043 90.48 ;
      RECT MASK 2 121.257 89.43 121.317 90.48 ;
      RECT MASK 2 121.531 89.43 121.591 90.48 ;
      RECT MASK 2 121.805 89.43 121.865 90.48 ;
      RECT MASK 2 122.079 89.43 122.139 90.48 ;
      RECT MASK 2 122.353 89.43 122.413 90.48 ;
      RECT MASK 2 122.627 89.43 122.687 90.48 ;
      RECT MASK 2 122.901 89.43 122.961 90.48 ;
      RECT MASK 2 123.175 89.43 123.235 90.48 ;
      RECT MASK 2 123.449 89.43 123.509 90.48 ;
      RECT MASK 2 123.723 89.43 123.783 90.48 ;
      RECT MASK 2 123.997 89.43 124.057 90.48 ;
      RECT MASK 2 124.271 89.43 124.331 90.48 ;
      RECT MASK 2 124.545 89.43 124.605 90.48 ;
      RECT MASK 2 124.819 89.43 124.879 90.48 ;
      RECT MASK 2 125.093 89.43 125.153 90.48 ;
      RECT MASK 2 125.367 89.43 125.427 90.48 ;
      RECT MASK 2 125.641 89.43 125.701 90.48 ;
      RECT MASK 2 125.915 89.43 125.975 90.48 ;
      RECT MASK 2 126.189 89.43 126.249 90.48 ;
      RECT MASK 2 126.463 89.43 126.523 90.48 ;
      RECT MASK 2 126.737 89.43 126.797 90.48 ;
      RECT MASK 2 127.011 89.43 127.071 90.48 ;
      RECT MASK 2 127.285 89.43 127.345 90.48 ;
      RECT MASK 2 127.559 89.43 127.619 90.48 ;
      RECT MASK 2 25.67 89.441 30.62 89.501 ;
      RECT MASK 2 9.2965 89.468 9.3565 89.692 ;
      RECT MASK 2 9.6285 89.468 9.6885 89.692 ;
      RECT MASK 2 9.9605 89.468 10.0205 89.692 ;
      RECT MASK 2 10.2925 89.468 10.3525 89.692 ;
      RECT MASK 2 10.6245 89.468 10.6845 89.692 ;
      RECT MASK 2 10.9565 89.468 11.0165 89.692 ;
      RECT MASK 2 11.2885 89.468 11.3485 89.692 ;
      RECT MASK 2 11.6205 89.468 11.6805 89.692 ;
      RECT MASK 2 14.3445 89.468 14.4045 89.692 ;
      RECT MASK 2 14.6765 89.468 14.7365 89.692 ;
      RECT MASK 2 15.0085 89.468 15.0685 89.692 ;
      RECT MASK 2 15.3405 89.468 15.4005 89.692 ;
      RECT MASK 2 15.6725 89.468 15.7325 89.692 ;
      RECT MASK 2 16.0045 89.468 16.0645 89.692 ;
      RECT MASK 2 18.5625 89.468 18.6225 89.692 ;
      RECT MASK 2 18.8945 89.468 18.9545 89.692 ;
      RECT MASK 2 19.2265 89.468 19.2865 89.692 ;
      RECT MASK 2 19.5585 89.468 19.6185 89.692 ;
      RECT MASK 2 19.8905 89.468 19.9505 89.692 ;
      RECT MASK 2 20.2225 89.468 20.2825 89.692 ;
      RECT MASK 2 20.5545 89.468 20.6145 89.692 ;
      RECT MASK 2 20.8865 89.468 20.9465 89.692 ;
      RECT MASK 2 21.2185 89.468 21.2785 89.692 ;
      RECT MASK 2 22.444 89.51 24.198 89.55 ;
      RECT MASK 2 2.204 89.52 2.264 90.57 ;
      RECT MASK 2 2.478 89.52 2.538 90.57 ;
      RECT MASK 2 2.752 89.52 2.812 90.57 ;
      RECT MASK 2 3.026 89.52 3.086 90.57 ;
      RECT MASK 2 3.3 89.52 3.36 90.57 ;
      RECT MASK 2 3.574 89.52 3.634 90.57 ;
      RECT MASK 2 3.848 89.52 3.908 90.57 ;
      RECT MASK 2 4.122 89.52 4.182 90.57 ;
      RECT MASK 2 4.396 89.52 4.456 90.57 ;
      RECT MASK 2 34.36 89.594 35.134 89.674 ;
      RECT MASK 2 67.676 89.594 68.276 89.674 ;
      RECT MASK 2 70.75 89.594 71.524 89.674 ;
      RECT MASK 2 104.058 89.594 104.832 89.674 ;
      RECT MASK 2 22.444 89.67 24.198 89.71 ;
      RECT MASK 2 25.67 89.703 30.62 89.763 ;
      RECT MASK 2 5.949 89.711 6.129 89.751 ;
      RECT MASK 2 6.945 89.711 7.125 89.751 ;
      RECT MASK 2 36.326 89.721 36.778 89.781 ;
      RECT MASK 2 37.048 89.721 65.754 89.781 ;
      RECT MASK 2 66.024 89.721 66.476 89.781 ;
      RECT MASK 2 72.716 89.721 73.168 89.781 ;
      RECT MASK 2 73.438 89.721 102.144 89.781 ;
      RECT MASK 2 102.414 89.721 102.866 89.781 ;
      RECT MASK 2 6.399 89.897 6.582 89.937 ;
      RECT MASK 2 34.36 89.906 35.134 89.986 ;
      RECT MASK 2 67.676 89.906 68.276 89.986 ;
      RECT MASK 2 70.75 89.906 71.524 89.986 ;
      RECT MASK 2 104.058 89.906 104.832 89.986 ;
      RECT MASK 2 22.444 89.93 24.198 89.97 ;
      RECT MASK 2 36.326 89.973 36.778 90.033 ;
      RECT MASK 2 37.048 89.973 65.754 90.033 ;
      RECT MASK 2 66.024 89.973 66.476 90.033 ;
      RECT MASK 2 72.716 89.973 73.168 90.033 ;
      RECT MASK 2 73.438 89.973 102.144 90.033 ;
      RECT MASK 2 102.414 89.973 102.866 90.033 ;
      RECT MASK 2 8.7735 89.99 12.2035 90.03 ;
      RECT MASK 2 13.8215 89.99 16.5875 90.03 ;
      RECT MASK 2 18.2055 89.99 21.6355 90.03 ;
      RECT MASK 2 5.949 90.081 7.125 90.121 ;
      RECT MASK 2 22.444 90.09 24.198 90.13 ;
      RECT MASK 2 8.7735 90.18 12.2035 90.22 ;
      RECT MASK 2 13.8215 90.18 16.5875 90.22 ;
      RECT MASK 2 18.2055 90.18 21.6355 90.22 ;
      RECT MASK 2 36.323 90.199 36.787 90.259 ;
      RECT MASK 2 37.047 90.199 65.755 90.259 ;
      RECT MASK 2 66.015 90.199 66.479 90.259 ;
      RECT MASK 2 72.713 90.199 73.177 90.259 ;
      RECT MASK 2 73.437 90.199 102.145 90.259 ;
      RECT MASK 2 102.405 90.199 102.869 90.259 ;
      RECT MASK 2 5.949 90.249 7.125 90.289 ;
      RECT MASK 2 25.67 90.297 25.938 90.357 ;
      RECT MASK 2 26.212 90.297 30.078 90.357 ;
      RECT MASK 2 30.352 90.297 30.62 90.357 ;
      RECT MASK 2 22.444 90.35 24.198 90.39 ;
      RECT MASK 2 34.36 90.434 35.134 90.514 ;
      RECT MASK 2 67.676 90.434 68.276 90.514 ;
      RECT MASK 2 70.75 90.434 71.524 90.514 ;
      RECT MASK 2 104.058 90.434 104.832 90.514 ;
      RECT MASK 2 8.16 90.44 12.807 90.48 ;
      RECT MASK 2 13.208 90.44 17.19 90.48 ;
      RECT MASK 2 17.592 90.44 22.239 90.48 ;
      RECT MASK 2 22.444 90.51 24.198 90.55 ;
      RECT MASK 2 36.326 90.621 66.476 90.681 ;
      RECT MASK 2 72.716 90.621 102.866 90.681 ;
      RECT MASK 2 8.16 90.63 12.807 90.67 ;
      RECT MASK 2 13.208 90.63 17.19 90.67 ;
      RECT MASK 2 17.592 90.63 22.239 90.67 ;
      RECT MASK 2 5.984 90.65 7.09 90.69 ;
      RECT MASK 2 34.36 90.746 35.134 90.826 ;
      RECT MASK 2 67.676 90.746 68.276 90.826 ;
      RECT MASK 2 70.75 90.746 71.524 90.826 ;
      RECT MASK 2 104.058 90.746 104.832 90.826 ;
      RECT MASK 2 22.444 90.77 24.198 90.81 ;
      RECT MASK 2 5.984 90.84 7.09 90.88 ;
      RECT MASK 2 36.326 90.873 66.476 90.933 ;
      RECT MASK 2 72.716 90.873 102.866 90.933 ;
      RECT MASK 2 25.67 90.881 30.62 90.941 ;
      RECT MASK 2 7.8125 90.89 12.807 90.93 ;
      RECT MASK 2 13.208 90.89 17.19 90.93 ;
      RECT MASK 2 17.592 90.89 22.239 90.93 ;
      RECT MASK 2 22.444 90.93 24.198 90.97 ;
      RECT MASK 2 108.379 90.93 108.439 91.98 ;
      RECT MASK 2 108.653 90.93 108.713 91.98 ;
      RECT MASK 2 108.927 90.93 108.987 91.98 ;
      RECT MASK 2 109.201 90.93 109.261 91.98 ;
      RECT MASK 2 109.475 90.93 109.535 91.98 ;
      RECT MASK 2 109.749 90.93 109.809 91.98 ;
      RECT MASK 2 110.023 90.93 110.083 91.98 ;
      RECT MASK 2 110.297 90.93 110.357 91.98 ;
      RECT MASK 2 110.571 90.93 110.631 91.98 ;
      RECT MASK 2 110.845 90.93 110.905 91.98 ;
      RECT MASK 2 111.119 90.93 111.179 91.98 ;
      RECT MASK 2 111.393 90.93 111.453 91.98 ;
      RECT MASK 2 111.667 90.93 111.727 91.98 ;
      RECT MASK 2 111.941 90.93 112.001 91.98 ;
      RECT MASK 2 112.215 90.93 112.275 91.98 ;
      RECT MASK 2 112.489 90.93 112.549 91.98 ;
      RECT MASK 2 112.763 90.93 112.823 91.98 ;
      RECT MASK 2 113.037 90.93 113.097 91.98 ;
      RECT MASK 2 113.311 90.93 113.371 91.98 ;
      RECT MASK 2 113.585 90.93 113.645 91.98 ;
      RECT MASK 2 113.859 90.93 113.919 91.98 ;
      RECT MASK 2 114.133 90.93 114.193 91.98 ;
      RECT MASK 2 114.407 90.93 114.467 91.98 ;
      RECT MASK 2 114.681 90.93 114.741 91.98 ;
      RECT MASK 2 114.955 90.93 115.015 91.98 ;
      RECT MASK 2 115.229 90.93 115.289 91.98 ;
      RECT MASK 2 115.503 90.93 115.563 91.98 ;
      RECT MASK 2 115.777 90.93 115.837 91.98 ;
      RECT MASK 2 116.051 90.93 116.111 91.98 ;
      RECT MASK 2 116.325 90.93 116.385 91.98 ;
      RECT MASK 2 116.599 90.93 116.659 91.98 ;
      RECT MASK 2 116.873 90.93 116.933 91.98 ;
      RECT MASK 2 117.147 90.93 117.207 91.98 ;
      RECT MASK 2 117.421 90.93 117.481 91.98 ;
      RECT MASK 2 117.695 90.93 117.755 91.98 ;
      RECT MASK 2 117.969 90.93 118.029 91.98 ;
      RECT MASK 2 118.243 90.93 118.303 91.98 ;
      RECT MASK 2 118.517 90.93 118.577 91.98 ;
      RECT MASK 2 118.791 90.93 118.851 91.98 ;
      RECT MASK 2 119.065 90.93 119.125 91.98 ;
      RECT MASK 2 119.339 90.93 119.399 91.98 ;
      RECT MASK 2 119.613 90.93 119.673 91.98 ;
      RECT MASK 2 119.887 90.93 119.947 91.98 ;
      RECT MASK 2 120.161 90.93 120.221 91.98 ;
      RECT MASK 2 120.435 90.93 120.495 91.98 ;
      RECT MASK 2 120.709 90.93 120.769 91.98 ;
      RECT MASK 2 120.983 90.93 121.043 91.98 ;
      RECT MASK 2 121.257 90.93 121.317 91.98 ;
      RECT MASK 2 121.531 90.93 121.591 91.98 ;
      RECT MASK 2 121.805 90.93 121.865 91.98 ;
      RECT MASK 2 122.079 90.93 122.139 91.98 ;
      RECT MASK 2 122.353 90.93 122.413 91.98 ;
      RECT MASK 2 122.627 90.93 122.687 91.98 ;
      RECT MASK 2 122.901 90.93 122.961 91.98 ;
      RECT MASK 2 123.175 90.93 123.235 91.98 ;
      RECT MASK 2 123.449 90.93 123.509 91.98 ;
      RECT MASK 2 123.723 90.93 123.783 91.98 ;
      RECT MASK 2 123.997 90.93 124.057 91.98 ;
      RECT MASK 2 124.271 90.93 124.331 91.98 ;
      RECT MASK 2 124.545 90.93 124.605 91.98 ;
      RECT MASK 2 124.819 90.93 124.879 91.98 ;
      RECT MASK 2 125.093 90.93 125.153 91.98 ;
      RECT MASK 2 125.367 90.93 125.427 91.98 ;
      RECT MASK 2 125.641 90.93 125.701 91.98 ;
      RECT MASK 2 125.915 90.93 125.975 91.98 ;
      RECT MASK 2 126.189 90.93 126.249 91.98 ;
      RECT MASK 2 126.463 90.93 126.523 91.98 ;
      RECT MASK 2 126.737 90.93 126.797 91.98 ;
      RECT MASK 2 127.011 90.93 127.071 91.98 ;
      RECT MASK 2 127.285 90.93 127.345 91.98 ;
      RECT MASK 2 127.559 90.93 127.619 91.98 ;
      RECT MASK 2 7.8125 91.08 12.807 91.12 ;
      RECT MASK 2 13.208 91.08 17.19 91.12 ;
      RECT MASK 2 17.592 91.08 22.239 91.12 ;
      RECT MASK 2 36.326 91.099 66.476 91.159 ;
      RECT MASK 2 72.716 91.099 102.866 91.159 ;
      RECT MASK 2 25.67 91.143 30.62 91.203 ;
      RECT MASK 2 71.997 91.16 72.269 91.22 ;
      RECT MASK 2 103.313 91.16 103.585 91.22 ;
      RECT MASK 2 22.444 91.19 24.198 91.23 ;
      RECT MASK 2 2.204 91.23 2.264 92.28 ;
      RECT MASK 2 2.478 91.23 2.538 92.28 ;
      RECT MASK 2 2.752 91.23 2.812 92.28 ;
      RECT MASK 2 3.026 91.23 3.086 92.28 ;
      RECT MASK 2 3.3 91.23 3.36 92.28 ;
      RECT MASK 2 3.574 91.23 3.634 92.28 ;
      RECT MASK 2 3.848 91.23 3.908 92.28 ;
      RECT MASK 2 4.122 91.23 4.182 92.28 ;
      RECT MASK 2 4.396 91.23 4.456 92.28 ;
      RECT MASK 2 5.949 91.271 7.125 91.311 ;
      RECT MASK 2 34.36 91.274 35.134 91.354 ;
      RECT MASK 2 67.676 91.274 68.276 91.354 ;
      RECT MASK 2 70.75 91.274 71.524 91.354 ;
      RECT MASK 2 104.058 91.274 104.832 91.354 ;
      RECT MASK 2 8.446 91.34 11.876 91.38 ;
      RECT MASK 2 13.8215 91.34 16.5875 91.38 ;
      RECT MASK 2 18.2055 91.34 21.6355 91.38 ;
      RECT MASK 2 22.444 91.35 24.198 91.39 ;
      RECT MASK 2 5.949 91.439 7.125 91.479 ;
      RECT MASK 2 36.326 91.521 36.778 91.581 ;
      RECT MASK 2 37.048 91.521 65.754 91.581 ;
      RECT MASK 2 66.024 91.521 66.476 91.581 ;
      RECT MASK 2 72.716 91.521 73.168 91.581 ;
      RECT MASK 2 73.438 91.521 102.144 91.581 ;
      RECT MASK 2 102.414 91.521 102.866 91.581 ;
      RECT MASK 2 8.446 91.53 11.876 91.57 ;
      RECT MASK 2 13.8215 91.53 16.5875 91.57 ;
      RECT MASK 2 18.2055 91.53 21.6355 91.57 ;
      RECT MASK 2 25.188 91.55 31.092 91.59 ;
      RECT MASK 2 34.36 91.586 35.134 91.666 ;
      RECT MASK 2 67.676 91.586 68.276 91.666 ;
      RECT MASK 2 70.75 91.586 71.524 91.666 ;
      RECT MASK 2 104.058 91.586 104.832 91.666 ;
      RECT MASK 2 22.444 91.61 24.198 91.65 ;
      RECT MASK 2 6.492 91.623 6.675 91.663 ;
      RECT MASK 2 25.188 91.71 31.092 91.75 ;
      RECT MASK 2 22.444 91.77 24.198 91.81 ;
      RECT MASK 2 36.326 91.773 36.778 91.833 ;
      RECT MASK 2 37.048 91.773 65.754 91.833 ;
      RECT MASK 2 66.024 91.773 66.476 91.833 ;
      RECT MASK 2 72.716 91.773 73.168 91.833 ;
      RECT MASK 2 73.438 91.773 102.144 91.833 ;
      RECT MASK 2 102.414 91.773 102.866 91.833 ;
      RECT MASK 2 5.949 91.809 6.129 91.849 ;
      RECT MASK 2 6.945 91.809 7.125 91.849 ;
      RECT MASK 2 8.969 91.868 9.029 92.092 ;
      RECT MASK 2 9.301 91.868 9.361 92.092 ;
      RECT MASK 2 9.633 91.868 9.693 92.092 ;
      RECT MASK 2 9.965 91.868 10.025 92.092 ;
      RECT MASK 2 10.297 91.868 10.357 92.092 ;
      RECT MASK 2 10.629 91.868 10.689 92.092 ;
      RECT MASK 2 10.961 91.868 11.021 92.092 ;
      RECT MASK 2 11.293 91.868 11.353 92.092 ;
      RECT MASK 2 14.3445 91.868 14.4045 92.092 ;
      RECT MASK 2 14.6765 91.868 14.7365 92.092 ;
      RECT MASK 2 15.0085 91.868 15.0685 92.092 ;
      RECT MASK 2 15.3405 91.868 15.4005 92.092 ;
      RECT MASK 2 15.6725 91.868 15.7325 92.092 ;
      RECT MASK 2 16.0045 91.868 16.0645 92.092 ;
      RECT MASK 2 18.5625 91.868 18.6225 92.092 ;
      RECT MASK 2 18.8945 91.868 18.9545 92.092 ;
      RECT MASK 2 19.2265 91.868 19.2865 92.092 ;
      RECT MASK 2 19.5585 91.868 19.6185 92.092 ;
      RECT MASK 2 19.8905 91.868 19.9505 92.092 ;
      RECT MASK 2 20.2225 91.868 20.2825 92.092 ;
      RECT MASK 2 20.5545 91.868 20.6145 92.092 ;
      RECT MASK 2 20.8865 91.868 20.9465 92.092 ;
      RECT MASK 2 21.2185 91.868 21.2785 92.092 ;
      RECT MASK 2 36.323 91.999 36.787 92.059 ;
      RECT MASK 2 37.047 91.999 65.755 92.059 ;
      RECT MASK 2 66.015 91.999 66.479 92.059 ;
      RECT MASK 2 72.713 91.999 73.177 92.059 ;
      RECT MASK 2 73.437 91.999 102.145 92.059 ;
      RECT MASK 2 102.405 91.999 102.869 92.059 ;
      RECT MASK 2 22.444 92.03 24.198 92.07 ;
      RECT MASK 2 34.36 92.114 35.134 92.194 ;
      RECT MASK 2 67.676 92.114 68.276 92.194 ;
      RECT MASK 2 70.75 92.114 71.524 92.194 ;
      RECT MASK 2 104.058 92.114 104.832 92.194 ;
      RECT MASK 2 25.237 92.149 31.053 92.289 ;
      RECT MASK 2 22.444 92.19 24.198 92.23 ;
      RECT MASK 2 8.66 92.25 9.172 92.29 ;
      RECT MASK 2 11.15 92.25 11.627 92.29 ;
      RECT MASK 2 14.0355 92.25 14.5475 92.29 ;
      RECT MASK 2 15.8615 92.25 16.3385 92.29 ;
      RECT MASK 2 18.4195 92.25 18.9315 92.29 ;
      RECT MASK 2 20.9095 92.25 21.3865 92.29 ;
      RECT MASK 2 5.984 92.255 7.09 92.295 ;
      RECT MASK 2 36.326 92.421 66.476 92.481 ;
      RECT MASK 2 72.716 92.421 102.866 92.481 ;
      RECT MASK 2 34.36 92.426 35.134 92.506 ;
      RECT MASK 2 67.676 92.426 68.276 92.506 ;
      RECT MASK 2 70.75 92.426 71.524 92.506 ;
      RECT MASK 2 104.058 92.426 104.832 92.506 ;
      RECT MASK 2 108.379 92.43 108.439 93.48 ;
      RECT MASK 2 108.653 92.43 108.713 93.48 ;
      RECT MASK 2 108.927 92.43 108.987 93.48 ;
      RECT MASK 2 109.201 92.43 109.261 93.48 ;
      RECT MASK 2 109.475 92.43 109.535 93.48 ;
      RECT MASK 2 109.749 92.43 109.809 93.48 ;
      RECT MASK 2 110.023 92.43 110.083 93.48 ;
      RECT MASK 2 110.297 92.43 110.357 93.48 ;
      RECT MASK 2 110.571 92.43 110.631 93.48 ;
      RECT MASK 2 110.845 92.43 110.905 93.48 ;
      RECT MASK 2 111.119 92.43 111.179 93.48 ;
      RECT MASK 2 111.393 92.43 111.453 93.48 ;
      RECT MASK 2 111.667 92.43 111.727 93.48 ;
      RECT MASK 2 111.941 92.43 112.001 93.48 ;
      RECT MASK 2 112.215 92.43 112.275 93.48 ;
      RECT MASK 2 112.489 92.43 112.549 93.48 ;
      RECT MASK 2 112.763 92.43 112.823 93.48 ;
      RECT MASK 2 113.037 92.43 113.097 93.48 ;
      RECT MASK 2 113.311 92.43 113.371 93.48 ;
      RECT MASK 2 113.585 92.43 113.645 93.48 ;
      RECT MASK 2 113.859 92.43 113.919 93.48 ;
      RECT MASK 2 114.133 92.43 114.193 93.48 ;
      RECT MASK 2 114.407 92.43 114.467 93.48 ;
      RECT MASK 2 114.681 92.43 114.741 93.48 ;
      RECT MASK 2 114.955 92.43 115.015 93.48 ;
      RECT MASK 2 115.229 92.43 115.289 93.48 ;
      RECT MASK 2 115.503 92.43 115.563 93.48 ;
      RECT MASK 2 115.777 92.43 115.837 93.48 ;
      RECT MASK 2 116.051 92.43 116.111 93.48 ;
      RECT MASK 2 116.325 92.43 116.385 93.48 ;
      RECT MASK 2 116.599 92.43 116.659 93.48 ;
      RECT MASK 2 116.873 92.43 116.933 93.48 ;
      RECT MASK 2 117.147 92.43 117.207 93.48 ;
      RECT MASK 2 117.421 92.43 117.481 93.48 ;
      RECT MASK 2 117.695 92.43 117.755 93.48 ;
      RECT MASK 2 117.969 92.43 118.029 93.48 ;
      RECT MASK 2 118.243 92.43 118.303 93.48 ;
      RECT MASK 2 118.517 92.43 118.577 93.48 ;
      RECT MASK 2 118.791 92.43 118.851 93.48 ;
      RECT MASK 2 119.065 92.43 119.125 93.48 ;
      RECT MASK 2 119.339 92.43 119.399 93.48 ;
      RECT MASK 2 119.613 92.43 119.673 93.48 ;
      RECT MASK 2 119.887 92.43 119.947 93.48 ;
      RECT MASK 2 120.161 92.43 120.221 93.48 ;
      RECT MASK 2 120.435 92.43 120.495 93.48 ;
      RECT MASK 2 120.709 92.43 120.769 93.48 ;
      RECT MASK 2 120.983 92.43 121.043 93.48 ;
      RECT MASK 2 121.257 92.43 121.317 93.48 ;
      RECT MASK 2 121.531 92.43 121.591 93.48 ;
      RECT MASK 2 121.805 92.43 121.865 93.48 ;
      RECT MASK 2 122.079 92.43 122.139 93.48 ;
      RECT MASK 2 122.353 92.43 122.413 93.48 ;
      RECT MASK 2 122.627 92.43 122.687 93.48 ;
      RECT MASK 2 122.901 92.43 122.961 93.48 ;
      RECT MASK 2 123.175 92.43 123.235 93.48 ;
      RECT MASK 2 123.449 92.43 123.509 93.48 ;
      RECT MASK 2 123.723 92.43 123.783 93.48 ;
      RECT MASK 2 123.997 92.43 124.057 93.48 ;
      RECT MASK 2 124.271 92.43 124.331 93.48 ;
      RECT MASK 2 124.545 92.43 124.605 93.48 ;
      RECT MASK 2 124.819 92.43 124.879 93.48 ;
      RECT MASK 2 125.093 92.43 125.153 93.48 ;
      RECT MASK 2 125.367 92.43 125.427 93.48 ;
      RECT MASK 2 125.641 92.43 125.701 93.48 ;
      RECT MASK 2 125.915 92.43 125.975 93.48 ;
      RECT MASK 2 126.189 92.43 126.249 93.48 ;
      RECT MASK 2 126.463 92.43 126.523 93.48 ;
      RECT MASK 2 126.737 92.43 126.797 93.48 ;
      RECT MASK 2 127.011 92.43 127.071 93.48 ;
      RECT MASK 2 127.285 92.43 127.345 93.48 ;
      RECT MASK 2 127.559 92.43 127.619 93.48 ;
      RECT MASK 2 8.66 92.45 9.172 92.49 ;
      RECT MASK 2 11.15 92.45 11.627 92.49 ;
      RECT MASK 2 14.0355 92.45 14.5475 92.49 ;
      RECT MASK 2 15.8615 92.45 16.3385 92.49 ;
      RECT MASK 2 18.4195 92.45 18.9315 92.49 ;
      RECT MASK 2 20.9095 92.45 21.3865 92.49 ;
      RECT MASK 2 22.444 92.45 24.198 92.49 ;
      RECT MASK 2 22.444 92.61 24.198 92.65 ;
      RECT MASK 2 8.969 92.648 9.029 92.872 ;
      RECT MASK 2 9.301 92.648 9.361 92.872 ;
      RECT MASK 2 9.633 92.648 9.693 92.872 ;
      RECT MASK 2 9.965 92.648 10.025 92.872 ;
      RECT MASK 2 10.297 92.648 10.357 92.872 ;
      RECT MASK 2 10.629 92.648 10.689 92.872 ;
      RECT MASK 2 10.961 92.648 11.021 92.872 ;
      RECT MASK 2 11.293 92.648 11.353 92.872 ;
      RECT MASK 2 14.3445 92.648 14.4045 92.872 ;
      RECT MASK 2 14.6765 92.648 14.7365 92.872 ;
      RECT MASK 2 15.0085 92.648 15.0685 92.872 ;
      RECT MASK 2 15.3405 92.648 15.4005 92.872 ;
      RECT MASK 2 15.6725 92.648 15.7325 92.872 ;
      RECT MASK 2 16.0045 92.648 16.0645 92.872 ;
      RECT MASK 2 18.5625 92.648 18.6225 92.872 ;
      RECT MASK 2 18.8945 92.648 18.9545 92.872 ;
      RECT MASK 2 19.2265 92.648 19.2865 92.872 ;
      RECT MASK 2 19.5585 92.648 19.6185 92.872 ;
      RECT MASK 2 19.8905 92.648 19.9505 92.872 ;
      RECT MASK 2 20.2225 92.648 20.2825 92.872 ;
      RECT MASK 2 20.5545 92.648 20.6145 92.872 ;
      RECT MASK 2 20.8865 92.648 20.9465 92.872 ;
      RECT MASK 2 21.2185 92.648 21.2785 92.872 ;
      RECT MASK 2 36.326 92.673 66.476 92.733 ;
      RECT MASK 2 72.716 92.673 102.866 92.733 ;
      RECT MASK 2 5.984 92.775 7.09 92.815 ;
      RECT MASK 2 22.444 92.87 24.198 92.91 ;
      RECT MASK 2 36.326 92.899 66.476 92.959 ;
      RECT MASK 2 72.716 92.899 102.866 92.959 ;
      RECT MASK 2 2.204 92.94 2.264 93.99 ;
      RECT MASK 2 2.478 92.94 2.538 93.99 ;
      RECT MASK 2 2.752 92.94 2.812 93.99 ;
      RECT MASK 2 3.026 92.94 3.086 93.99 ;
      RECT MASK 2 3.3 92.94 3.36 93.99 ;
      RECT MASK 2 3.574 92.94 3.634 93.99 ;
      RECT MASK 2 3.848 92.94 3.908 93.99 ;
      RECT MASK 2 4.122 92.94 4.182 93.99 ;
      RECT MASK 2 4.396 92.94 4.456 93.99 ;
      RECT MASK 2 34.36 92.954 35.134 93.034 ;
      RECT MASK 2 67.676 92.954 68.276 93.034 ;
      RECT MASK 2 70.75 92.954 71.524 93.034 ;
      RECT MASK 2 104.058 92.954 104.832 93.034 ;
      RECT MASK 2 71.997 92.96 72.269 93.02 ;
      RECT MASK 2 103.313 92.96 103.585 93.02 ;
      RECT MASK 2 22.444 93.03 24.198 93.07 ;
      RECT MASK 2 5.949 93.185 6.129 93.225 ;
      RECT MASK 2 6.945 93.185 7.125 93.225 ;
      RECT MASK 2 8.778 93.2 11.544 93.24 ;
      RECT MASK 2 14.1405 93.2 16.2815 93.24 ;
      RECT MASK 2 18.5375 93.2 21.3035 93.24 ;
      RECT MASK 2 34.36 93.266 35.134 93.346 ;
      RECT MASK 2 67.676 93.266 68.276 93.346 ;
      RECT MASK 2 70.75 93.266 71.524 93.346 ;
      RECT MASK 2 104.058 93.266 104.832 93.346 ;
      RECT MASK 2 22.444 93.29 24.198 93.33 ;
      RECT MASK 2 36.326 93.321 36.778 93.381 ;
      RECT MASK 2 37.048 93.321 65.754 93.381 ;
      RECT MASK 2 66.024 93.321 66.476 93.381 ;
      RECT MASK 2 72.716 93.321 73.168 93.381 ;
      RECT MASK 2 73.438 93.321 102.144 93.381 ;
      RECT MASK 2 102.414 93.321 102.866 93.381 ;
      RECT MASK 2 8.778 93.39 11.544 93.43 ;
      RECT MASK 2 14.1405 93.39 16.2815 93.43 ;
      RECT MASK 2 18.5375 93.39 21.3035 93.43 ;
      RECT MASK 2 6.399 93.407 6.582 93.447 ;
      RECT MASK 2 22.444 93.45 24.198 93.49 ;
      RECT MASK 2 36.326 93.573 36.778 93.633 ;
      RECT MASK 2 37.048 93.573 65.754 93.633 ;
      RECT MASK 2 66.024 93.573 66.476 93.633 ;
      RECT MASK 2 72.716 93.573 73.168 93.633 ;
      RECT MASK 2 73.438 93.573 102.144 93.633 ;
      RECT MASK 2 102.414 93.573 102.866 93.633 ;
      RECT MASK 2 5.92 93.591 7.154 93.631 ;
      RECT MASK 2 8.446 93.65 11.876 93.69 ;
      RECT MASK 2 13.8215 93.65 16.5875 93.69 ;
      RECT MASK 2 18.2055 93.65 21.6355 93.69 ;
      RECT MASK 2 22.444 93.71 24.198 93.75 ;
      RECT MASK 2 5.92 93.759 7.154 93.799 ;
      RECT MASK 2 34.36 93.794 35.134 93.874 ;
      RECT MASK 2 67.676 93.794 68.276 93.874 ;
      RECT MASK 2 70.75 93.794 71.524 93.874 ;
      RECT MASK 2 104.058 93.794 104.832 93.874 ;
      RECT MASK 2 36.323 93.799 36.787 93.859 ;
      RECT MASK 2 37.047 93.799 65.755 93.859 ;
      RECT MASK 2 66.015 93.799 66.479 93.859 ;
      RECT MASK 2 72.713 93.799 73.177 93.859 ;
      RECT MASK 2 73.437 93.799 102.145 93.859 ;
      RECT MASK 2 102.405 93.799 102.869 93.859 ;
      RECT MASK 2 8.446 93.84 11.876 93.88 ;
      RECT MASK 2 13.8215 93.84 16.5875 93.88 ;
      RECT MASK 2 18.2055 93.84 21.6355 93.88 ;
      RECT MASK 2 22.444 93.87 24.198 93.91 ;
      RECT MASK 2 25.237 93.871 31.053 94.011 ;
      RECT MASK 2 108.379 93.93 108.439 94.98 ;
      RECT MASK 2 108.653 93.93 108.713 94.98 ;
      RECT MASK 2 108.927 93.93 108.987 94.98 ;
      RECT MASK 2 109.201 93.93 109.261 94.98 ;
      RECT MASK 2 109.475 93.93 109.535 94.98 ;
      RECT MASK 2 109.749 93.93 109.809 94.98 ;
      RECT MASK 2 110.023 93.93 110.083 94.98 ;
      RECT MASK 2 110.297 93.93 110.357 94.98 ;
      RECT MASK 2 110.571 93.93 110.631 94.98 ;
      RECT MASK 2 110.845 93.93 110.905 94.98 ;
      RECT MASK 2 111.119 93.93 111.179 94.98 ;
      RECT MASK 2 111.393 93.93 111.453 94.98 ;
      RECT MASK 2 111.667 93.93 111.727 94.98 ;
      RECT MASK 2 111.941 93.93 112.001 94.98 ;
      RECT MASK 2 112.215 93.93 112.275 94.98 ;
      RECT MASK 2 112.489 93.93 112.549 94.98 ;
      RECT MASK 2 112.763 93.93 112.823 94.98 ;
      RECT MASK 2 113.037 93.93 113.097 94.98 ;
      RECT MASK 2 113.311 93.93 113.371 94.98 ;
      RECT MASK 2 113.585 93.93 113.645 94.98 ;
      RECT MASK 2 113.859 93.93 113.919 94.98 ;
      RECT MASK 2 114.133 93.93 114.193 94.98 ;
      RECT MASK 2 114.407 93.93 114.467 94.98 ;
      RECT MASK 2 114.681 93.93 114.741 94.98 ;
      RECT MASK 2 114.955 93.93 115.015 94.98 ;
      RECT MASK 2 115.229 93.93 115.289 94.98 ;
      RECT MASK 2 115.503 93.93 115.563 94.98 ;
      RECT MASK 2 115.777 93.93 115.837 94.98 ;
      RECT MASK 2 116.051 93.93 116.111 94.98 ;
      RECT MASK 2 116.325 93.93 116.385 94.98 ;
      RECT MASK 2 116.599 93.93 116.659 94.98 ;
      RECT MASK 2 116.873 93.93 116.933 94.98 ;
      RECT MASK 2 117.147 93.93 117.207 94.98 ;
      RECT MASK 2 117.421 93.93 117.481 94.98 ;
      RECT MASK 2 117.695 93.93 117.755 94.98 ;
      RECT MASK 2 117.969 93.93 118.029 94.98 ;
      RECT MASK 2 118.243 93.93 118.303 94.98 ;
      RECT MASK 2 118.517 93.93 118.577 94.98 ;
      RECT MASK 2 118.791 93.93 118.851 94.98 ;
      RECT MASK 2 119.065 93.93 119.125 94.98 ;
      RECT MASK 2 119.339 93.93 119.399 94.98 ;
      RECT MASK 2 119.613 93.93 119.673 94.98 ;
      RECT MASK 2 119.887 93.93 119.947 94.98 ;
      RECT MASK 2 120.161 93.93 120.221 94.98 ;
      RECT MASK 2 120.435 93.93 120.495 94.98 ;
      RECT MASK 2 120.709 93.93 120.769 94.98 ;
      RECT MASK 2 120.983 93.93 121.043 94.98 ;
      RECT MASK 2 121.257 93.93 121.317 94.98 ;
      RECT MASK 2 121.531 93.93 121.591 94.98 ;
      RECT MASK 2 121.805 93.93 121.865 94.98 ;
      RECT MASK 2 122.079 93.93 122.139 94.98 ;
      RECT MASK 2 122.353 93.93 122.413 94.98 ;
      RECT MASK 2 122.627 93.93 122.687 94.98 ;
      RECT MASK 2 122.901 93.93 122.961 94.98 ;
      RECT MASK 2 123.175 93.93 123.235 94.98 ;
      RECT MASK 2 123.449 93.93 123.509 94.98 ;
      RECT MASK 2 123.723 93.93 123.783 94.98 ;
      RECT MASK 2 123.997 93.93 124.057 94.98 ;
      RECT MASK 2 124.271 93.93 124.331 94.98 ;
      RECT MASK 2 124.545 93.93 124.605 94.98 ;
      RECT MASK 2 124.819 93.93 124.879 94.98 ;
      RECT MASK 2 125.093 93.93 125.153 94.98 ;
      RECT MASK 2 125.367 93.93 125.427 94.98 ;
      RECT MASK 2 125.641 93.93 125.701 94.98 ;
      RECT MASK 2 125.915 93.93 125.975 94.98 ;
      RECT MASK 2 126.189 93.93 126.249 94.98 ;
      RECT MASK 2 126.463 93.93 126.523 94.98 ;
      RECT MASK 2 126.737 93.93 126.797 94.98 ;
      RECT MASK 2 127.011 93.93 127.071 94.98 ;
      RECT MASK 2 127.285 93.93 127.345 94.98 ;
      RECT MASK 2 127.559 93.93 127.619 94.98 ;
      RECT MASK 2 5.984 94.1 12.811 94.14 ;
      RECT MASK 2 13.208 94.1 17.19 94.14 ;
      RECT MASK 2 17.592 94.1 22.239 94.14 ;
      RECT MASK 2 34.36 94.106 35.134 94.186 ;
      RECT MASK 2 67.676 94.106 68.276 94.186 ;
      RECT MASK 2 70.75 94.106 71.524 94.186 ;
      RECT MASK 2 104.058 94.106 104.832 94.186 ;
      RECT MASK 2 22.444 94.13 24.198 94.17 ;
      RECT MASK 2 36.326 94.221 66.476 94.281 ;
      RECT MASK 2 72.716 94.221 102.866 94.281 ;
      RECT MASK 2 5.984 94.29 12.811 94.33 ;
      RECT MASK 2 13.208 94.29 17.19 94.33 ;
      RECT MASK 2 17.592 94.29 22.239 94.33 ;
      RECT MASK 2 22.444 94.29 24.198 94.33 ;
      RECT MASK 2 36.326 94.473 66.476 94.533 ;
      RECT MASK 2 72.716 94.473 102.866 94.533 ;
      RECT MASK 2 22.444 94.55 31.502 94.59 ;
      RECT MASK 2 33.739 94.64 35.338 94.68 ;
      RECT MASK 2 67.467 94.64 68.897 94.68 ;
      RECT MASK 2 2.204 94.65 2.264 95.7 ;
      RECT MASK 2 2.478 94.65 2.538 95.7 ;
      RECT MASK 2 2.752 94.65 2.812 95.7 ;
      RECT MASK 2 3.026 94.65 3.086 95.7 ;
      RECT MASK 2 3.3 94.65 3.36 95.7 ;
      RECT MASK 2 3.574 94.65 3.634 95.7 ;
      RECT MASK 2 3.848 94.65 3.908 95.7 ;
      RECT MASK 2 4.122 94.65 4.182 95.7 ;
      RECT MASK 2 4.396 94.65 4.456 95.7 ;
      RECT MASK 2 36.326 94.699 66.476 94.759 ;
      RECT MASK 2 72.716 94.699 102.866 94.759 ;
      RECT MASK 2 22.444 94.71 31.502 94.75 ;
      RECT MASK 2 70.129 94.73 71.728 94.77 ;
      RECT MASK 2 103.854 94.73 105.453 94.77 ;
      RECT MASK 2 71.997 94.76 72.269 94.82 ;
      RECT MASK 2 103.313 94.76 103.585 94.82 ;
      RECT MASK 2 33.739 94.83 35.338 94.87 ;
      RECT MASK 2 67.467 94.83 68.897 94.87 ;
      RECT MASK 2 70.129 94.92 71.728 94.96 ;
      RECT MASK 2 103.854 94.92 105.453 94.96 ;
      RECT MASK 2 22.444 94.97 31.502 95.01 ;
      RECT MASK 2 33.407 95.09 35.338 95.13 ;
      RECT MASK 2 67.467 95.09 69.229 95.13 ;
      RECT MASK 2 22.444 95.13 31.502 95.17 ;
      RECT MASK 2 69.797 95.18 71.728 95.22 ;
      RECT MASK 2 103.854 95.18 105.785 95.22 ;
      RECT MASK 2 33.407 95.28 35.338 95.32 ;
      RECT MASK 2 67.467 95.28 69.229 95.32 ;
      RECT MASK 2 71.997 95.361 103.585 95.421 ;
      RECT MASK 2 69.797 95.37 71.728 95.41 ;
      RECT MASK 2 103.854 95.37 105.785 95.41 ;
      RECT MASK 2 22.444 95.39 31.502 95.43 ;
      RECT MASK 2 108.379 95.43 108.439 96.48 ;
      RECT MASK 2 108.653 95.43 108.713 96.48 ;
      RECT MASK 2 108.927 95.43 108.987 96.48 ;
      RECT MASK 2 109.201 95.43 109.261 96.48 ;
      RECT MASK 2 109.475 95.43 109.535 96.48 ;
      RECT MASK 2 109.749 95.43 109.809 96.48 ;
      RECT MASK 2 110.023 95.43 110.083 96.48 ;
      RECT MASK 2 110.297 95.43 110.357 96.48 ;
      RECT MASK 2 110.571 95.43 110.631 96.48 ;
      RECT MASK 2 110.845 95.43 110.905 96.48 ;
      RECT MASK 2 111.119 95.43 111.179 96.48 ;
      RECT MASK 2 111.393 95.43 111.453 96.48 ;
      RECT MASK 2 111.667 95.43 111.727 96.48 ;
      RECT MASK 2 111.941 95.43 112.001 96.48 ;
      RECT MASK 2 112.215 95.43 112.275 96.48 ;
      RECT MASK 2 112.489 95.43 112.549 96.48 ;
      RECT MASK 2 112.763 95.43 112.823 96.48 ;
      RECT MASK 2 113.037 95.43 113.097 96.48 ;
      RECT MASK 2 113.311 95.43 113.371 96.48 ;
      RECT MASK 2 113.585 95.43 113.645 96.48 ;
      RECT MASK 2 113.859 95.43 113.919 96.48 ;
      RECT MASK 2 114.133 95.43 114.193 96.48 ;
      RECT MASK 2 114.407 95.43 114.467 96.48 ;
      RECT MASK 2 114.681 95.43 114.741 96.48 ;
      RECT MASK 2 114.955 95.43 115.015 96.48 ;
      RECT MASK 2 115.229 95.43 115.289 96.48 ;
      RECT MASK 2 115.503 95.43 115.563 96.48 ;
      RECT MASK 2 115.777 95.43 115.837 96.48 ;
      RECT MASK 2 116.051 95.43 116.111 96.48 ;
      RECT MASK 2 116.325 95.43 116.385 96.48 ;
      RECT MASK 2 116.599 95.43 116.659 96.48 ;
      RECT MASK 2 116.873 95.43 116.933 96.48 ;
      RECT MASK 2 117.147 95.43 117.207 96.48 ;
      RECT MASK 2 117.421 95.43 117.481 96.48 ;
      RECT MASK 2 117.695 95.43 117.755 96.48 ;
      RECT MASK 2 117.969 95.43 118.029 96.48 ;
      RECT MASK 2 118.243 95.43 118.303 96.48 ;
      RECT MASK 2 118.517 95.43 118.577 96.48 ;
      RECT MASK 2 118.791 95.43 118.851 96.48 ;
      RECT MASK 2 119.065 95.43 119.125 96.48 ;
      RECT MASK 2 119.339 95.43 119.399 96.48 ;
      RECT MASK 2 119.613 95.43 119.673 96.48 ;
      RECT MASK 2 119.887 95.43 119.947 96.48 ;
      RECT MASK 2 120.161 95.43 120.221 96.48 ;
      RECT MASK 2 120.435 95.43 120.495 96.48 ;
      RECT MASK 2 120.709 95.43 120.769 96.48 ;
      RECT MASK 2 120.983 95.43 121.043 96.48 ;
      RECT MASK 2 121.257 95.43 121.317 96.48 ;
      RECT MASK 2 121.531 95.43 121.591 96.48 ;
      RECT MASK 2 121.805 95.43 121.865 96.48 ;
      RECT MASK 2 122.079 95.43 122.139 96.48 ;
      RECT MASK 2 122.353 95.43 122.413 96.48 ;
      RECT MASK 2 122.627 95.43 122.687 96.48 ;
      RECT MASK 2 122.901 95.43 122.961 96.48 ;
      RECT MASK 2 123.175 95.43 123.235 96.48 ;
      RECT MASK 2 123.449 95.43 123.509 96.48 ;
      RECT MASK 2 123.723 95.43 123.783 96.48 ;
      RECT MASK 2 123.997 95.43 124.057 96.48 ;
      RECT MASK 2 124.271 95.43 124.331 96.48 ;
      RECT MASK 2 124.545 95.43 124.605 96.48 ;
      RECT MASK 2 124.819 95.43 124.879 96.48 ;
      RECT MASK 2 125.093 95.43 125.153 96.48 ;
      RECT MASK 2 125.367 95.43 125.427 96.48 ;
      RECT MASK 2 125.641 95.43 125.701 96.48 ;
      RECT MASK 2 125.915 95.43 125.975 96.48 ;
      RECT MASK 2 126.189 95.43 126.249 96.48 ;
      RECT MASK 2 126.463 95.43 126.523 96.48 ;
      RECT MASK 2 126.737 95.43 126.797 96.48 ;
      RECT MASK 2 127.011 95.43 127.071 96.48 ;
      RECT MASK 2 127.285 95.43 127.345 96.48 ;
      RECT MASK 2 127.559 95.43 127.619 96.48 ;
      RECT MASK 2 22.444 95.55 31.502 95.59 ;
      RECT MASK 2 22.444 95.81 36.656 95.85 ;
      RECT MASK 2 22.444 95.97 36.656 96.01 ;
      RECT MASK 2 1.248 96.14 5.362 96.18 ;
      RECT MASK 2 22.444 96.23 36.656 96.27 ;
      RECT MASK 2 1.248 96.33 5.362 96.37 ;
      RECT MASK 2 22.444 96.39 36.656 96.43 ;
      RECT MASK 2 107.479 96.83 128.525 96.87 ;
      RECT MASK 2 107.479 97.02 128.525 97.06 ;
      RECT MASK 2 1.439 97.28 44.397 97.32 ;
      RECT MASK 2 44.831 97.28 87.789 97.32 ;
      RECT MASK 2 88.223 97.28 128.525 97.32 ;
      RECT MASK 2 1.439 97.47 44.397 97.51 ;
      RECT MASK 2 44.831 97.47 87.789 97.51 ;
      RECT MASK 2 88.223 97.47 128.525 97.51 ;
      RECT MASK 2 2.338 97.83 2.398 98.88 ;
      RECT MASK 2 2.612 97.83 2.672 98.88 ;
      RECT MASK 2 2.886 97.83 2.946 98.88 ;
      RECT MASK 2 3.16 97.83 3.22 98.88 ;
      RECT MASK 2 3.434 97.83 3.494 98.88 ;
      RECT MASK 2 3.708 97.83 3.768 98.88 ;
      RECT MASK 2 3.982 97.83 4.042 98.88 ;
      RECT MASK 2 4.256 97.83 4.316 98.88 ;
      RECT MASK 2 4.53 97.83 4.59 98.88 ;
      RECT MASK 2 4.804 97.83 4.864 98.88 ;
      RECT MASK 2 5.078 97.83 5.138 98.88 ;
      RECT MASK 2 5.352 97.83 5.412 98.88 ;
      RECT MASK 2 5.626 97.83 5.686 98.88 ;
      RECT MASK 2 5.9 97.83 5.96 98.88 ;
      RECT MASK 2 6.174 97.83 6.234 98.88 ;
      RECT MASK 2 6.448 97.83 6.508 98.88 ;
      RECT MASK 2 6.722 97.83 6.782 98.88 ;
      RECT MASK 2 6.996 97.83 7.056 98.88 ;
      RECT MASK 2 7.27 97.83 7.33 98.88 ;
      RECT MASK 2 7.544 97.83 7.604 98.88 ;
      RECT MASK 2 7.818 97.83 7.878 98.88 ;
      RECT MASK 2 8.092 97.83 8.152 98.88 ;
      RECT MASK 2 8.366 97.83 8.426 98.88 ;
      RECT MASK 2 8.64 97.83 8.7 98.88 ;
      RECT MASK 2 8.914 97.83 8.974 98.88 ;
      RECT MASK 2 9.188 97.83 9.248 98.88 ;
      RECT MASK 2 9.462 97.83 9.522 98.88 ;
      RECT MASK 2 9.736 97.83 9.796 98.88 ;
      RECT MASK 2 10.01 97.83 10.07 98.88 ;
      RECT MASK 2 10.284 97.83 10.344 98.88 ;
      RECT MASK 2 10.558 97.83 10.618 98.88 ;
      RECT MASK 2 10.832 97.83 10.892 98.88 ;
      RECT MASK 2 11.106 97.83 11.166 98.88 ;
      RECT MASK 2 11.38 97.83 11.44 98.88 ;
      RECT MASK 2 11.654 97.83 11.714 98.88 ;
      RECT MASK 2 11.928 97.83 11.988 98.88 ;
      RECT MASK 2 12.202 97.83 12.262 98.88 ;
      RECT MASK 2 12.476 97.83 12.536 98.88 ;
      RECT MASK 2 12.75 97.83 12.81 98.88 ;
      RECT MASK 2 13.024 97.83 13.084 98.88 ;
      RECT MASK 2 13.298 97.83 13.358 98.88 ;
      RECT MASK 2 13.572 97.83 13.632 98.88 ;
      RECT MASK 2 13.846 97.83 13.906 98.88 ;
      RECT MASK 2 14.12 97.83 14.18 98.88 ;
      RECT MASK 2 14.394 97.83 14.454 98.88 ;
      RECT MASK 2 14.668 97.83 14.728 98.88 ;
      RECT MASK 2 14.942 97.83 15.002 98.88 ;
      RECT MASK 2 15.216 97.83 15.276 98.88 ;
      RECT MASK 2 15.49 97.83 15.55 98.88 ;
      RECT MASK 2 15.764 97.83 15.824 98.88 ;
      RECT MASK 2 16.038 97.83 16.098 98.88 ;
      RECT MASK 2 16.312 97.83 16.372 98.88 ;
      RECT MASK 2 16.586 97.83 16.646 98.88 ;
      RECT MASK 2 16.86 97.83 16.92 98.88 ;
      RECT MASK 2 17.134 97.83 17.194 98.88 ;
      RECT MASK 2 17.408 97.83 17.468 98.88 ;
      RECT MASK 2 17.682 97.83 17.742 98.88 ;
      RECT MASK 2 17.956 97.83 18.016 98.88 ;
      RECT MASK 2 18.23 97.83 18.29 98.88 ;
      RECT MASK 2 18.504 97.83 18.564 98.88 ;
      RECT MASK 2 18.778 97.83 18.838 98.88 ;
      RECT MASK 2 19.052 97.83 19.112 98.88 ;
      RECT MASK 2 19.326 97.83 19.386 98.88 ;
      RECT MASK 2 19.6 97.83 19.66 98.88 ;
      RECT MASK 2 19.874 97.83 19.934 98.88 ;
      RECT MASK 2 20.148 97.83 20.208 98.88 ;
      RECT MASK 2 20.422 97.83 20.482 98.88 ;
      RECT MASK 2 20.696 97.83 20.756 98.88 ;
      RECT MASK 2 20.97 97.83 21.03 98.88 ;
      RECT MASK 2 21.244 97.83 21.304 98.88 ;
      RECT MASK 2 21.518 97.83 21.578 98.88 ;
      RECT MASK 2 21.792 97.83 21.852 98.88 ;
      RECT MASK 2 22.066 97.83 22.126 98.88 ;
      RECT MASK 2 22.34 97.83 22.4 98.88 ;
      RECT MASK 2 22.614 97.83 22.674 98.88 ;
      RECT MASK 2 22.888 97.83 22.948 98.88 ;
      RECT MASK 2 23.162 97.83 23.222 98.88 ;
      RECT MASK 2 23.436 97.83 23.496 98.88 ;
      RECT MASK 2 23.71 97.83 23.77 98.88 ;
      RECT MASK 2 23.984 97.83 24.044 98.88 ;
      RECT MASK 2 24.258 97.83 24.318 98.88 ;
      RECT MASK 2 24.532 97.83 24.592 98.88 ;
      RECT MASK 2 24.806 97.83 24.866 98.88 ;
      RECT MASK 2 25.08 97.83 25.14 98.88 ;
      RECT MASK 2 25.354 97.83 25.414 98.88 ;
      RECT MASK 2 25.628 97.83 25.688 98.88 ;
      RECT MASK 2 25.902 97.83 25.962 98.88 ;
      RECT MASK 2 26.176 97.83 26.236 98.88 ;
      RECT MASK 2 26.45 97.83 26.51 98.88 ;
      RECT MASK 2 26.724 97.83 26.784 98.88 ;
      RECT MASK 2 26.998 97.83 27.058 98.88 ;
      RECT MASK 2 27.272 97.83 27.332 98.88 ;
      RECT MASK 2 27.546 97.83 27.606 98.88 ;
      RECT MASK 2 27.82 97.83 27.88 98.88 ;
      RECT MASK 2 28.094 97.83 28.154 98.88 ;
      RECT MASK 2 28.368 97.83 28.428 98.88 ;
      RECT MASK 2 28.642 97.83 28.702 98.88 ;
      RECT MASK 2 28.916 97.83 28.976 98.88 ;
      RECT MASK 2 29.19 97.83 29.25 98.88 ;
      RECT MASK 2 29.464 97.83 29.524 98.88 ;
      RECT MASK 2 29.738 97.83 29.798 98.88 ;
      RECT MASK 2 30.012 97.83 30.072 98.88 ;
      RECT MASK 2 30.286 97.83 30.346 98.88 ;
      RECT MASK 2 30.56 97.83 30.62 98.88 ;
      RECT MASK 2 30.834 97.83 30.894 98.88 ;
      RECT MASK 2 31.108 97.83 31.168 98.88 ;
      RECT MASK 2 31.382 97.83 31.442 98.88 ;
      RECT MASK 2 31.656 97.83 31.716 98.88 ;
      RECT MASK 2 31.93 97.83 31.99 98.88 ;
      RECT MASK 2 32.204 97.83 32.264 98.88 ;
      RECT MASK 2 32.478 97.83 32.538 98.88 ;
      RECT MASK 2 32.752 97.83 32.812 98.88 ;
      RECT MASK 2 33.026 97.83 33.086 98.88 ;
      RECT MASK 2 33.3 97.83 33.36 98.88 ;
      RECT MASK 2 33.574 97.83 33.634 98.88 ;
      RECT MASK 2 33.848 97.83 33.908 98.88 ;
      RECT MASK 2 34.122 97.83 34.182 98.88 ;
      RECT MASK 2 34.396 97.83 34.456 98.88 ;
      RECT MASK 2 34.67 97.83 34.73 98.88 ;
      RECT MASK 2 34.944 97.83 35.004 98.88 ;
      RECT MASK 2 35.218 97.83 35.278 98.88 ;
      RECT MASK 2 35.492 97.83 35.552 98.88 ;
      RECT MASK 2 35.766 97.83 35.826 98.88 ;
      RECT MASK 2 36.04 97.83 36.1 98.88 ;
      RECT MASK 2 36.314 97.83 36.374 98.88 ;
      RECT MASK 2 36.588 97.83 36.648 98.88 ;
      RECT MASK 2 36.862 97.83 36.922 98.88 ;
      RECT MASK 2 37.136 97.83 37.196 98.88 ;
      RECT MASK 2 37.41 97.83 37.47 98.88 ;
      RECT MASK 2 37.684 97.83 37.744 98.88 ;
      RECT MASK 2 37.958 97.83 38.018 98.88 ;
      RECT MASK 2 38.232 97.83 38.292 98.88 ;
      RECT MASK 2 38.506 97.83 38.566 98.88 ;
      RECT MASK 2 38.78 97.83 38.84 98.88 ;
      RECT MASK 2 39.054 97.83 39.114 98.88 ;
      RECT MASK 2 39.328 97.83 39.388 98.88 ;
      RECT MASK 2 39.602 97.83 39.662 98.88 ;
      RECT MASK 2 39.876 97.83 39.936 98.88 ;
      RECT MASK 2 40.15 97.83 40.21 98.88 ;
      RECT MASK 2 40.424 97.83 40.484 98.88 ;
      RECT MASK 2 40.698 97.83 40.758 98.88 ;
      RECT MASK 2 40.972 97.83 41.032 98.88 ;
      RECT MASK 2 41.246 97.83 41.306 98.88 ;
      RECT MASK 2 41.52 97.83 41.58 98.88 ;
      RECT MASK 2 41.794 97.83 41.854 98.88 ;
      RECT MASK 2 42.068 97.83 42.128 98.88 ;
      RECT MASK 2 42.342 97.83 42.402 98.88 ;
      RECT MASK 2 42.616 97.83 42.676 98.88 ;
      RECT MASK 2 42.89 97.83 42.95 98.88 ;
      RECT MASK 2 43.164 97.83 43.224 98.88 ;
      RECT MASK 2 43.438 97.83 43.498 98.88 ;
      RECT MASK 2 45.73 97.83 45.79 98.88 ;
      RECT MASK 2 46.004 97.83 46.064 98.88 ;
      RECT MASK 2 46.278 97.83 46.338 98.88 ;
      RECT MASK 2 46.552 97.83 46.612 98.88 ;
      RECT MASK 2 46.826 97.83 46.886 98.88 ;
      RECT MASK 2 47.1 97.83 47.16 98.88 ;
      RECT MASK 2 47.374 97.83 47.434 98.88 ;
      RECT MASK 2 47.648 97.83 47.708 98.88 ;
      RECT MASK 2 47.922 97.83 47.982 98.88 ;
      RECT MASK 2 48.196 97.83 48.256 98.88 ;
      RECT MASK 2 48.47 97.83 48.53 98.88 ;
      RECT MASK 2 48.744 97.83 48.804 98.88 ;
      RECT MASK 2 49.018 97.83 49.078 98.88 ;
      RECT MASK 2 49.292 97.83 49.352 98.88 ;
      RECT MASK 2 49.566 97.83 49.626 98.88 ;
      RECT MASK 2 49.84 97.83 49.9 98.88 ;
      RECT MASK 2 50.114 97.83 50.174 98.88 ;
      RECT MASK 2 50.388 97.83 50.448 98.88 ;
      RECT MASK 2 50.662 97.83 50.722 98.88 ;
      RECT MASK 2 50.936 97.83 50.996 98.88 ;
      RECT MASK 2 51.21 97.83 51.27 98.88 ;
      RECT MASK 2 51.484 97.83 51.544 98.88 ;
      RECT MASK 2 51.758 97.83 51.818 98.88 ;
      RECT MASK 2 52.032 97.83 52.092 98.88 ;
      RECT MASK 2 52.306 97.83 52.366 98.88 ;
      RECT MASK 2 52.58 97.83 52.64 98.88 ;
      RECT MASK 2 52.854 97.83 52.914 98.88 ;
      RECT MASK 2 53.128 97.83 53.188 98.88 ;
      RECT MASK 2 53.402 97.83 53.462 98.88 ;
      RECT MASK 2 53.676 97.83 53.736 98.88 ;
      RECT MASK 2 53.95 97.83 54.01 98.88 ;
      RECT MASK 2 54.224 97.83 54.284 98.88 ;
      RECT MASK 2 54.498 97.83 54.558 98.88 ;
      RECT MASK 2 54.772 97.83 54.832 98.88 ;
      RECT MASK 2 55.046 97.83 55.106 98.88 ;
      RECT MASK 2 55.32 97.83 55.38 98.88 ;
      RECT MASK 2 55.594 97.83 55.654 98.88 ;
      RECT MASK 2 55.868 97.83 55.928 98.88 ;
      RECT MASK 2 56.142 97.83 56.202 98.88 ;
      RECT MASK 2 56.416 97.83 56.476 98.88 ;
      RECT MASK 2 56.69 97.83 56.75 98.88 ;
      RECT MASK 2 56.964 97.83 57.024 98.88 ;
      RECT MASK 2 57.238 97.83 57.298 98.88 ;
      RECT MASK 2 57.512 97.83 57.572 98.88 ;
      RECT MASK 2 57.786 97.83 57.846 98.88 ;
      RECT MASK 2 58.06 97.83 58.12 98.88 ;
      RECT MASK 2 58.334 97.83 58.394 98.88 ;
      RECT MASK 2 58.608 97.83 58.668 98.88 ;
      RECT MASK 2 58.882 97.83 58.942 98.88 ;
      RECT MASK 2 59.156 97.83 59.216 98.88 ;
      RECT MASK 2 59.43 97.83 59.49 98.88 ;
      RECT MASK 2 59.704 97.83 59.764 98.88 ;
      RECT MASK 2 59.978 97.83 60.038 98.88 ;
      RECT MASK 2 60.252 97.83 60.312 98.88 ;
      RECT MASK 2 60.526 97.83 60.586 98.88 ;
      RECT MASK 2 60.8 97.83 60.86 98.88 ;
      RECT MASK 2 61.074 97.83 61.134 98.88 ;
      RECT MASK 2 61.348 97.83 61.408 98.88 ;
      RECT MASK 2 61.622 97.83 61.682 98.88 ;
      RECT MASK 2 61.896 97.83 61.956 98.88 ;
      RECT MASK 2 62.17 97.83 62.23 98.88 ;
      RECT MASK 2 62.444 97.83 62.504 98.88 ;
      RECT MASK 2 62.718 97.83 62.778 98.88 ;
      RECT MASK 2 62.992 97.83 63.052 98.88 ;
      RECT MASK 2 63.266 97.83 63.326 98.88 ;
      RECT MASK 2 63.54 97.83 63.6 98.88 ;
      RECT MASK 2 63.814 97.83 63.874 98.88 ;
      RECT MASK 2 64.088 97.83 64.148 98.88 ;
      RECT MASK 2 64.362 97.83 64.422 98.88 ;
      RECT MASK 2 64.636 97.83 64.696 98.88 ;
      RECT MASK 2 64.91 97.83 64.97 98.88 ;
      RECT MASK 2 65.184 97.83 65.244 98.88 ;
      RECT MASK 2 65.458 97.83 65.518 98.88 ;
      RECT MASK 2 65.732 97.83 65.792 98.88 ;
      RECT MASK 2 66.006 97.83 66.066 98.88 ;
      RECT MASK 2 66.28 97.83 66.34 98.88 ;
      RECT MASK 2 66.554 97.83 66.614 98.88 ;
      RECT MASK 2 66.828 97.83 66.888 98.88 ;
      RECT MASK 2 67.102 97.83 67.162 98.88 ;
      RECT MASK 2 67.376 97.83 67.436 98.88 ;
      RECT MASK 2 67.65 97.83 67.71 98.88 ;
      RECT MASK 2 67.924 97.83 67.984 98.88 ;
      RECT MASK 2 68.198 97.83 68.258 98.88 ;
      RECT MASK 2 68.472 97.83 68.532 98.88 ;
      RECT MASK 2 68.746 97.83 68.806 98.88 ;
      RECT MASK 2 69.02 97.83 69.08 98.88 ;
      RECT MASK 2 69.294 97.83 69.354 98.88 ;
      RECT MASK 2 69.568 97.83 69.628 98.88 ;
      RECT MASK 2 69.842 97.83 69.902 98.88 ;
      RECT MASK 2 70.116 97.83 70.176 98.88 ;
      RECT MASK 2 70.39 97.83 70.45 98.88 ;
      RECT MASK 2 70.664 97.83 70.724 98.88 ;
      RECT MASK 2 70.938 97.83 70.998 98.88 ;
      RECT MASK 2 71.212 97.83 71.272 98.88 ;
      RECT MASK 2 71.486 97.83 71.546 98.88 ;
      RECT MASK 2 71.76 97.83 71.82 98.88 ;
      RECT MASK 2 72.034 97.83 72.094 98.88 ;
      RECT MASK 2 72.308 97.83 72.368 98.88 ;
      RECT MASK 2 72.582 97.83 72.642 98.88 ;
      RECT MASK 2 72.856 97.83 72.916 98.88 ;
      RECT MASK 2 73.13 97.83 73.19 98.88 ;
      RECT MASK 2 73.404 97.83 73.464 98.88 ;
      RECT MASK 2 73.678 97.83 73.738 98.88 ;
      RECT MASK 2 73.952 97.83 74.012 98.88 ;
      RECT MASK 2 74.226 97.83 74.286 98.88 ;
      RECT MASK 2 74.5 97.83 74.56 98.88 ;
      RECT MASK 2 74.774 97.83 74.834 98.88 ;
      RECT MASK 2 75.048 97.83 75.108 98.88 ;
      RECT MASK 2 75.322 97.83 75.382 98.88 ;
      RECT MASK 2 75.596 97.83 75.656 98.88 ;
      RECT MASK 2 75.87 97.83 75.93 98.88 ;
      RECT MASK 2 76.144 97.83 76.204 98.88 ;
      RECT MASK 2 76.418 97.83 76.478 98.88 ;
      RECT MASK 2 76.692 97.83 76.752 98.88 ;
      RECT MASK 2 76.966 97.83 77.026 98.88 ;
      RECT MASK 2 77.24 97.83 77.3 98.88 ;
      RECT MASK 2 77.514 97.83 77.574 98.88 ;
      RECT MASK 2 77.788 97.83 77.848 98.88 ;
      RECT MASK 2 78.062 97.83 78.122 98.88 ;
      RECT MASK 2 78.336 97.83 78.396 98.88 ;
      RECT MASK 2 78.61 97.83 78.67 98.88 ;
      RECT MASK 2 78.884 97.83 78.944 98.88 ;
      RECT MASK 2 79.158 97.83 79.218 98.88 ;
      RECT MASK 2 79.432 97.83 79.492 98.88 ;
      RECT MASK 2 79.706 97.83 79.766 98.88 ;
      RECT MASK 2 79.98 97.83 80.04 98.88 ;
      RECT MASK 2 80.254 97.83 80.314 98.88 ;
      RECT MASK 2 80.528 97.83 80.588 98.88 ;
      RECT MASK 2 80.802 97.83 80.862 98.88 ;
      RECT MASK 2 81.076 97.83 81.136 98.88 ;
      RECT MASK 2 81.35 97.83 81.41 98.88 ;
      RECT MASK 2 81.624 97.83 81.684 98.88 ;
      RECT MASK 2 81.898 97.83 81.958 98.88 ;
      RECT MASK 2 82.172 97.83 82.232 98.88 ;
      RECT MASK 2 82.446 97.83 82.506 98.88 ;
      RECT MASK 2 82.72 97.83 82.78 98.88 ;
      RECT MASK 2 82.994 97.83 83.054 98.88 ;
      RECT MASK 2 83.268 97.83 83.328 98.88 ;
      RECT MASK 2 83.542 97.83 83.602 98.88 ;
      RECT MASK 2 83.816 97.83 83.876 98.88 ;
      RECT MASK 2 84.09 97.83 84.15 98.88 ;
      RECT MASK 2 84.364 97.83 84.424 98.88 ;
      RECT MASK 2 84.638 97.83 84.698 98.88 ;
      RECT MASK 2 84.912 97.83 84.972 98.88 ;
      RECT MASK 2 85.186 97.83 85.246 98.88 ;
      RECT MASK 2 85.46 97.83 85.52 98.88 ;
      RECT MASK 2 85.734 97.83 85.794 98.88 ;
      RECT MASK 2 86.008 97.83 86.068 98.88 ;
      RECT MASK 2 86.282 97.83 86.342 98.88 ;
      RECT MASK 2 86.556 97.83 86.616 98.88 ;
      RECT MASK 2 86.83 97.83 86.89 98.88 ;
      RECT MASK 2 89.089 97.83 89.149 98.88 ;
      RECT MASK 2 89.363 97.83 89.423 98.88 ;
      RECT MASK 2 89.637 97.83 89.697 98.88 ;
      RECT MASK 2 89.911 97.83 89.971 98.88 ;
      RECT MASK 2 90.185 97.83 90.245 98.88 ;
      RECT MASK 2 90.459 97.83 90.519 98.88 ;
      RECT MASK 2 90.733 97.83 90.793 98.88 ;
      RECT MASK 2 91.007 97.83 91.067 98.88 ;
      RECT MASK 2 91.281 97.83 91.341 98.88 ;
      RECT MASK 2 91.555 97.83 91.615 98.88 ;
      RECT MASK 2 91.829 97.83 91.889 98.88 ;
      RECT MASK 2 92.103 97.83 92.163 98.88 ;
      RECT MASK 2 92.377 97.83 92.437 98.88 ;
      RECT MASK 2 92.651 97.83 92.711 98.88 ;
      RECT MASK 2 92.925 97.83 92.985 98.88 ;
      RECT MASK 2 93.199 97.83 93.259 98.88 ;
      RECT MASK 2 93.473 97.83 93.533 98.88 ;
      RECT MASK 2 93.747 97.83 93.807 98.88 ;
      RECT MASK 2 94.021 97.83 94.081 98.88 ;
      RECT MASK 2 94.295 97.83 94.355 98.88 ;
      RECT MASK 2 94.569 97.83 94.629 98.88 ;
      RECT MASK 2 94.843 97.83 94.903 98.88 ;
      RECT MASK 2 95.117 97.83 95.177 98.88 ;
      RECT MASK 2 95.391 97.83 95.451 98.88 ;
      RECT MASK 2 95.665 97.83 95.725 98.88 ;
      RECT MASK 2 95.939 97.83 95.999 98.88 ;
      RECT MASK 2 96.213 97.83 96.273 98.88 ;
      RECT MASK 2 96.487 97.83 96.547 98.88 ;
      RECT MASK 2 96.761 97.83 96.821 98.88 ;
      RECT MASK 2 97.035 97.83 97.095 98.88 ;
      RECT MASK 2 97.309 97.83 97.369 98.88 ;
      RECT MASK 2 97.583 97.83 97.643 98.88 ;
      RECT MASK 2 97.857 97.83 97.917 98.88 ;
      RECT MASK 2 98.131 97.83 98.191 98.88 ;
      RECT MASK 2 98.405 97.83 98.465 98.88 ;
      RECT MASK 2 98.679 97.83 98.739 98.88 ;
      RECT MASK 2 98.953 97.83 99.013 98.88 ;
      RECT MASK 2 99.227 97.83 99.287 98.88 ;
      RECT MASK 2 99.501 97.83 99.561 98.88 ;
      RECT MASK 2 99.775 97.83 99.835 98.88 ;
      RECT MASK 2 100.049 97.83 100.109 98.88 ;
      RECT MASK 2 100.323 97.83 100.383 98.88 ;
      RECT MASK 2 100.597 97.83 100.657 98.88 ;
      RECT MASK 2 100.871 97.83 100.931 98.88 ;
      RECT MASK 2 101.145 97.83 101.205 98.88 ;
      RECT MASK 2 101.419 97.83 101.479 98.88 ;
      RECT MASK 2 101.693 97.83 101.753 98.88 ;
      RECT MASK 2 101.967 97.83 102.027 98.88 ;
      RECT MASK 2 102.241 97.83 102.301 98.88 ;
      RECT MASK 2 102.515 97.83 102.575 98.88 ;
      RECT MASK 2 102.789 97.83 102.849 98.88 ;
      RECT MASK 2 103.063 97.83 103.123 98.88 ;
      RECT MASK 2 103.337 97.83 103.397 98.88 ;
      RECT MASK 2 103.611 97.83 103.671 98.88 ;
      RECT MASK 2 103.885 97.83 103.945 98.88 ;
      RECT MASK 2 104.159 97.83 104.219 98.88 ;
      RECT MASK 2 104.433 97.83 104.493 98.88 ;
      RECT MASK 2 104.707 97.83 104.767 98.88 ;
      RECT MASK 2 104.981 97.83 105.041 98.88 ;
      RECT MASK 2 105.255 97.83 105.315 98.88 ;
      RECT MASK 2 105.529 97.83 105.589 98.88 ;
      RECT MASK 2 105.803 97.83 105.863 98.88 ;
      RECT MASK 2 106.077 97.83 106.137 98.88 ;
      RECT MASK 2 106.351 97.83 106.411 98.88 ;
      RECT MASK 2 106.625 97.83 106.685 98.88 ;
      RECT MASK 2 106.899 97.83 106.959 98.88 ;
      RECT MASK 2 107.173 97.83 107.233 98.88 ;
      RECT MASK 2 107.447 97.83 107.507 98.88 ;
      RECT MASK 2 107.721 97.83 107.781 98.88 ;
      RECT MASK 2 107.995 97.83 108.055 98.88 ;
      RECT MASK 2 108.269 97.83 108.329 98.88 ;
      RECT MASK 2 108.543 97.83 108.603 98.88 ;
      RECT MASK 2 108.817 97.83 108.877 98.88 ;
      RECT MASK 2 109.091 97.83 109.151 98.88 ;
      RECT MASK 2 109.365 97.83 109.425 98.88 ;
      RECT MASK 2 109.639 97.83 109.699 98.88 ;
      RECT MASK 2 109.913 97.83 109.973 98.88 ;
      RECT MASK 2 110.187 97.83 110.247 98.88 ;
      RECT MASK 2 110.461 97.83 110.521 98.88 ;
      RECT MASK 2 110.735 97.83 110.795 98.88 ;
      RECT MASK 2 111.009 97.83 111.069 98.88 ;
      RECT MASK 2 111.283 97.83 111.343 98.88 ;
      RECT MASK 2 111.557 97.83 111.617 98.88 ;
      RECT MASK 2 111.831 97.83 111.891 98.88 ;
      RECT MASK 2 112.105 97.83 112.165 98.88 ;
      RECT MASK 2 112.379 97.83 112.439 98.88 ;
      RECT MASK 2 112.653 97.83 112.713 98.88 ;
      RECT MASK 2 112.927 97.83 112.987 98.88 ;
      RECT MASK 2 113.201 97.83 113.261 98.88 ;
      RECT MASK 2 113.475 97.83 113.535 98.88 ;
      RECT MASK 2 113.749 97.83 113.809 98.88 ;
      RECT MASK 2 114.023 97.83 114.083 98.88 ;
      RECT MASK 2 114.297 97.83 114.357 98.88 ;
      RECT MASK 2 114.571 97.83 114.631 98.88 ;
      RECT MASK 2 114.845 97.83 114.905 98.88 ;
      RECT MASK 2 115.119 97.83 115.179 98.88 ;
      RECT MASK 2 115.393 97.83 115.453 98.88 ;
      RECT MASK 2 115.667 97.83 115.727 98.88 ;
      RECT MASK 2 115.941 97.83 116.001 98.88 ;
      RECT MASK 2 116.215 97.83 116.275 98.88 ;
      RECT MASK 2 116.489 97.83 116.549 98.88 ;
      RECT MASK 2 116.763 97.83 116.823 98.88 ;
      RECT MASK 2 117.037 97.83 117.097 98.88 ;
      RECT MASK 2 117.311 97.83 117.371 98.88 ;
      RECT MASK 2 117.585 97.83 117.645 98.88 ;
      RECT MASK 2 117.859 97.83 117.919 98.88 ;
      RECT MASK 2 118.133 97.83 118.193 98.88 ;
      RECT MASK 2 118.407 97.83 118.467 98.88 ;
      RECT MASK 2 118.681 97.83 118.741 98.88 ;
      RECT MASK 2 118.955 97.83 119.015 98.88 ;
      RECT MASK 2 119.229 97.83 119.289 98.88 ;
      RECT MASK 2 119.503 97.83 119.563 98.88 ;
      RECT MASK 2 119.777 97.83 119.837 98.88 ;
      RECT MASK 2 120.051 97.83 120.111 98.88 ;
      RECT MASK 2 120.325 97.83 120.385 98.88 ;
      RECT MASK 2 120.599 97.83 120.659 98.88 ;
      RECT MASK 2 120.873 97.83 120.933 98.88 ;
      RECT MASK 2 121.147 97.83 121.207 98.88 ;
      RECT MASK 2 121.421 97.83 121.481 98.88 ;
      RECT MASK 2 121.695 97.83 121.755 98.88 ;
      RECT MASK 2 121.969 97.83 122.029 98.88 ;
      RECT MASK 2 122.243 97.83 122.303 98.88 ;
      RECT MASK 2 122.517 97.83 122.577 98.88 ;
      RECT MASK 2 122.791 97.83 122.851 98.88 ;
      RECT MASK 2 123.065 97.83 123.125 98.88 ;
      RECT MASK 2 123.339 97.83 123.399 98.88 ;
      RECT MASK 2 123.613 97.83 123.673 98.88 ;
      RECT MASK 2 123.887 97.83 123.947 98.88 ;
      RECT MASK 2 124.161 97.83 124.221 98.88 ;
      RECT MASK 2 124.435 97.83 124.495 98.88 ;
      RECT MASK 2 124.709 97.83 124.769 98.88 ;
      RECT MASK 2 124.983 97.83 125.043 98.88 ;
      RECT MASK 2 125.257 97.83 125.317 98.88 ;
      RECT MASK 2 125.531 97.83 125.591 98.88 ;
      RECT MASK 2 125.805 97.83 125.865 98.88 ;
      RECT MASK 2 126.079 97.83 126.139 98.88 ;
      RECT MASK 2 126.353 97.83 126.413 98.88 ;
      RECT MASK 2 126.627 97.83 126.687 98.88 ;
      RECT MASK 2 126.901 97.83 126.961 98.88 ;
      RECT MASK 2 127.175 97.83 127.235 98.88 ;
      RECT MASK 2 127.449 97.83 127.509 98.88 ;
      RECT MASK 2 2.338 99.54 2.398 100.59 ;
      RECT MASK 2 2.612 99.54 2.672 100.59 ;
      RECT MASK 2 2.886 99.54 2.946 100.59 ;
      RECT MASK 2 3.16 99.54 3.22 100.59 ;
      RECT MASK 2 3.434 99.54 3.494 100.59 ;
      RECT MASK 2 3.708 99.54 3.768 100.59 ;
      RECT MASK 2 3.982 99.54 4.042 100.59 ;
      RECT MASK 2 4.256 99.54 4.316 100.59 ;
      RECT MASK 2 4.53 99.54 4.59 100.59 ;
      RECT MASK 2 4.804 99.54 4.864 100.59 ;
      RECT MASK 2 5.078 99.54 5.138 100.59 ;
      RECT MASK 2 5.352 99.54 5.412 100.59 ;
      RECT MASK 2 5.626 99.54 5.686 100.59 ;
      RECT MASK 2 5.9 99.54 5.96 100.59 ;
      RECT MASK 2 6.174 99.54 6.234 100.59 ;
      RECT MASK 2 6.448 99.54 6.508 100.59 ;
      RECT MASK 2 6.722 99.54 6.782 100.59 ;
      RECT MASK 2 6.996 99.54 7.056 100.59 ;
      RECT MASK 2 7.27 99.54 7.33 100.59 ;
      RECT MASK 2 7.544 99.54 7.604 100.59 ;
      RECT MASK 2 7.818 99.54 7.878 100.59 ;
      RECT MASK 2 8.092 99.54 8.152 100.59 ;
      RECT MASK 2 8.366 99.54 8.426 100.59 ;
      RECT MASK 2 8.64 99.54 8.7 100.59 ;
      RECT MASK 2 8.914 99.54 8.974 100.59 ;
      RECT MASK 2 9.188 99.54 9.248 100.59 ;
      RECT MASK 2 9.462 99.54 9.522 100.59 ;
      RECT MASK 2 9.736 99.54 9.796 100.59 ;
      RECT MASK 2 10.01 99.54 10.07 100.59 ;
      RECT MASK 2 10.284 99.54 10.344 100.59 ;
      RECT MASK 2 10.558 99.54 10.618 100.59 ;
      RECT MASK 2 10.832 99.54 10.892 100.59 ;
      RECT MASK 2 11.106 99.54 11.166 100.59 ;
      RECT MASK 2 11.38 99.54 11.44 100.59 ;
      RECT MASK 2 11.654 99.54 11.714 100.59 ;
      RECT MASK 2 11.928 99.54 11.988 100.59 ;
      RECT MASK 2 12.202 99.54 12.262 100.59 ;
      RECT MASK 2 12.476 99.54 12.536 100.59 ;
      RECT MASK 2 12.75 99.54 12.81 100.59 ;
      RECT MASK 2 13.024 99.54 13.084 100.59 ;
      RECT MASK 2 13.298 99.54 13.358 100.59 ;
      RECT MASK 2 13.572 99.54 13.632 100.59 ;
      RECT MASK 2 13.846 99.54 13.906 100.59 ;
      RECT MASK 2 14.12 99.54 14.18 100.59 ;
      RECT MASK 2 14.394 99.54 14.454 100.59 ;
      RECT MASK 2 14.668 99.54 14.728 100.59 ;
      RECT MASK 2 14.942 99.54 15.002 100.59 ;
      RECT MASK 2 15.216 99.54 15.276 100.59 ;
      RECT MASK 2 15.49 99.54 15.55 100.59 ;
      RECT MASK 2 15.764 99.54 15.824 100.59 ;
      RECT MASK 2 16.038 99.54 16.098 100.59 ;
      RECT MASK 2 16.312 99.54 16.372 100.59 ;
      RECT MASK 2 16.586 99.54 16.646 100.59 ;
      RECT MASK 2 16.86 99.54 16.92 100.59 ;
      RECT MASK 2 17.134 99.54 17.194 100.59 ;
      RECT MASK 2 17.408 99.54 17.468 100.59 ;
      RECT MASK 2 17.682 99.54 17.742 100.59 ;
      RECT MASK 2 17.956 99.54 18.016 100.59 ;
      RECT MASK 2 18.23 99.54 18.29 100.59 ;
      RECT MASK 2 18.504 99.54 18.564 100.59 ;
      RECT MASK 2 18.778 99.54 18.838 100.59 ;
      RECT MASK 2 19.052 99.54 19.112 100.59 ;
      RECT MASK 2 19.326 99.54 19.386 100.59 ;
      RECT MASK 2 19.6 99.54 19.66 100.59 ;
      RECT MASK 2 19.874 99.54 19.934 100.59 ;
      RECT MASK 2 20.148 99.54 20.208 100.59 ;
      RECT MASK 2 20.422 99.54 20.482 100.59 ;
      RECT MASK 2 20.696 99.54 20.756 100.59 ;
      RECT MASK 2 20.97 99.54 21.03 100.59 ;
      RECT MASK 2 21.244 99.54 21.304 100.59 ;
      RECT MASK 2 21.518 99.54 21.578 100.59 ;
      RECT MASK 2 21.792 99.54 21.852 100.59 ;
      RECT MASK 2 22.066 99.54 22.126 100.59 ;
      RECT MASK 2 22.34 99.54 22.4 100.59 ;
      RECT MASK 2 22.614 99.54 22.674 100.59 ;
      RECT MASK 2 22.888 99.54 22.948 100.59 ;
      RECT MASK 2 23.162 99.54 23.222 100.59 ;
      RECT MASK 2 23.436 99.54 23.496 100.59 ;
      RECT MASK 2 23.71 99.54 23.77 100.59 ;
      RECT MASK 2 23.984 99.54 24.044 100.59 ;
      RECT MASK 2 24.258 99.54 24.318 100.59 ;
      RECT MASK 2 24.532 99.54 24.592 100.59 ;
      RECT MASK 2 24.806 99.54 24.866 100.59 ;
      RECT MASK 2 25.08 99.54 25.14 100.59 ;
      RECT MASK 2 25.354 99.54 25.414 100.59 ;
      RECT MASK 2 25.628 99.54 25.688 100.59 ;
      RECT MASK 2 25.902 99.54 25.962 100.59 ;
      RECT MASK 2 26.176 99.54 26.236 100.59 ;
      RECT MASK 2 26.45 99.54 26.51 100.59 ;
      RECT MASK 2 26.724 99.54 26.784 100.59 ;
      RECT MASK 2 26.998 99.54 27.058 100.59 ;
      RECT MASK 2 27.272 99.54 27.332 100.59 ;
      RECT MASK 2 27.546 99.54 27.606 100.59 ;
      RECT MASK 2 27.82 99.54 27.88 100.59 ;
      RECT MASK 2 28.094 99.54 28.154 100.59 ;
      RECT MASK 2 28.368 99.54 28.428 100.59 ;
      RECT MASK 2 28.642 99.54 28.702 100.59 ;
      RECT MASK 2 28.916 99.54 28.976 100.59 ;
      RECT MASK 2 29.19 99.54 29.25 100.59 ;
      RECT MASK 2 29.464 99.54 29.524 100.59 ;
      RECT MASK 2 29.738 99.54 29.798 100.59 ;
      RECT MASK 2 30.012 99.54 30.072 100.59 ;
      RECT MASK 2 30.286 99.54 30.346 100.59 ;
      RECT MASK 2 30.56 99.54 30.62 100.59 ;
      RECT MASK 2 30.834 99.54 30.894 100.59 ;
      RECT MASK 2 31.108 99.54 31.168 100.59 ;
      RECT MASK 2 31.382 99.54 31.442 100.59 ;
      RECT MASK 2 31.656 99.54 31.716 100.59 ;
      RECT MASK 2 31.93 99.54 31.99 100.59 ;
      RECT MASK 2 32.204 99.54 32.264 100.59 ;
      RECT MASK 2 32.478 99.54 32.538 100.59 ;
      RECT MASK 2 32.752 99.54 32.812 100.59 ;
      RECT MASK 2 33.026 99.54 33.086 100.59 ;
      RECT MASK 2 33.3 99.54 33.36 100.59 ;
      RECT MASK 2 33.574 99.54 33.634 100.59 ;
      RECT MASK 2 33.848 99.54 33.908 100.59 ;
      RECT MASK 2 34.122 99.54 34.182 100.59 ;
      RECT MASK 2 34.396 99.54 34.456 100.59 ;
      RECT MASK 2 34.67 99.54 34.73 100.59 ;
      RECT MASK 2 34.944 99.54 35.004 100.59 ;
      RECT MASK 2 35.218 99.54 35.278 100.59 ;
      RECT MASK 2 35.492 99.54 35.552 100.59 ;
      RECT MASK 2 35.766 99.54 35.826 100.59 ;
      RECT MASK 2 36.04 99.54 36.1 100.59 ;
      RECT MASK 2 36.314 99.54 36.374 100.59 ;
      RECT MASK 2 36.588 99.54 36.648 100.59 ;
      RECT MASK 2 36.862 99.54 36.922 100.59 ;
      RECT MASK 2 37.136 99.54 37.196 100.59 ;
      RECT MASK 2 37.41 99.54 37.47 100.59 ;
      RECT MASK 2 37.684 99.54 37.744 100.59 ;
      RECT MASK 2 37.958 99.54 38.018 100.59 ;
      RECT MASK 2 38.232 99.54 38.292 100.59 ;
      RECT MASK 2 38.506 99.54 38.566 100.59 ;
      RECT MASK 2 38.78 99.54 38.84 100.59 ;
      RECT MASK 2 39.054 99.54 39.114 100.59 ;
      RECT MASK 2 39.328 99.54 39.388 100.59 ;
      RECT MASK 2 39.602 99.54 39.662 100.59 ;
      RECT MASK 2 39.876 99.54 39.936 100.59 ;
      RECT MASK 2 40.15 99.54 40.21 100.59 ;
      RECT MASK 2 40.424 99.54 40.484 100.59 ;
      RECT MASK 2 40.698 99.54 40.758 100.59 ;
      RECT MASK 2 40.972 99.54 41.032 100.59 ;
      RECT MASK 2 41.246 99.54 41.306 100.59 ;
      RECT MASK 2 41.52 99.54 41.58 100.59 ;
      RECT MASK 2 41.794 99.54 41.854 100.59 ;
      RECT MASK 2 42.068 99.54 42.128 100.59 ;
      RECT MASK 2 42.342 99.54 42.402 100.59 ;
      RECT MASK 2 42.616 99.54 42.676 100.59 ;
      RECT MASK 2 42.89 99.54 42.95 100.59 ;
      RECT MASK 2 43.164 99.54 43.224 100.59 ;
      RECT MASK 2 43.438 99.54 43.498 100.59 ;
      RECT MASK 2 45.73 99.54 45.79 100.59 ;
      RECT MASK 2 46.004 99.54 46.064 100.59 ;
      RECT MASK 2 46.278 99.54 46.338 100.59 ;
      RECT MASK 2 46.552 99.54 46.612 100.59 ;
      RECT MASK 2 46.826 99.54 46.886 100.59 ;
      RECT MASK 2 47.1 99.54 47.16 100.59 ;
      RECT MASK 2 47.374 99.54 47.434 100.59 ;
      RECT MASK 2 47.648 99.54 47.708 100.59 ;
      RECT MASK 2 47.922 99.54 47.982 100.59 ;
      RECT MASK 2 48.196 99.54 48.256 100.59 ;
      RECT MASK 2 48.47 99.54 48.53 100.59 ;
      RECT MASK 2 48.744 99.54 48.804 100.59 ;
      RECT MASK 2 49.018 99.54 49.078 100.59 ;
      RECT MASK 2 49.292 99.54 49.352 100.59 ;
      RECT MASK 2 49.566 99.54 49.626 100.59 ;
      RECT MASK 2 49.84 99.54 49.9 100.59 ;
      RECT MASK 2 50.114 99.54 50.174 100.59 ;
      RECT MASK 2 50.388 99.54 50.448 100.59 ;
      RECT MASK 2 50.662 99.54 50.722 100.59 ;
      RECT MASK 2 50.936 99.54 50.996 100.59 ;
      RECT MASK 2 51.21 99.54 51.27 100.59 ;
      RECT MASK 2 51.484 99.54 51.544 100.59 ;
      RECT MASK 2 51.758 99.54 51.818 100.59 ;
      RECT MASK 2 52.032 99.54 52.092 100.59 ;
      RECT MASK 2 52.306 99.54 52.366 100.59 ;
      RECT MASK 2 52.58 99.54 52.64 100.59 ;
      RECT MASK 2 52.854 99.54 52.914 100.59 ;
      RECT MASK 2 53.128 99.54 53.188 100.59 ;
      RECT MASK 2 53.402 99.54 53.462 100.59 ;
      RECT MASK 2 53.676 99.54 53.736 100.59 ;
      RECT MASK 2 53.95 99.54 54.01 100.59 ;
      RECT MASK 2 54.224 99.54 54.284 100.59 ;
      RECT MASK 2 54.498 99.54 54.558 100.59 ;
      RECT MASK 2 54.772 99.54 54.832 100.59 ;
      RECT MASK 2 55.046 99.54 55.106 100.59 ;
      RECT MASK 2 55.32 99.54 55.38 100.59 ;
      RECT MASK 2 55.594 99.54 55.654 100.59 ;
      RECT MASK 2 55.868 99.54 55.928 100.59 ;
      RECT MASK 2 56.142 99.54 56.202 100.59 ;
      RECT MASK 2 56.416 99.54 56.476 100.59 ;
      RECT MASK 2 56.69 99.54 56.75 100.59 ;
      RECT MASK 2 56.964 99.54 57.024 100.59 ;
      RECT MASK 2 57.238 99.54 57.298 100.59 ;
      RECT MASK 2 57.512 99.54 57.572 100.59 ;
      RECT MASK 2 57.786 99.54 57.846 100.59 ;
      RECT MASK 2 58.06 99.54 58.12 100.59 ;
      RECT MASK 2 58.334 99.54 58.394 100.59 ;
      RECT MASK 2 58.608 99.54 58.668 100.59 ;
      RECT MASK 2 58.882 99.54 58.942 100.59 ;
      RECT MASK 2 59.156 99.54 59.216 100.59 ;
      RECT MASK 2 59.43 99.54 59.49 100.59 ;
      RECT MASK 2 59.704 99.54 59.764 100.59 ;
      RECT MASK 2 59.978 99.54 60.038 100.59 ;
      RECT MASK 2 60.252 99.54 60.312 100.59 ;
      RECT MASK 2 60.526 99.54 60.586 100.59 ;
      RECT MASK 2 60.8 99.54 60.86 100.59 ;
      RECT MASK 2 61.074 99.54 61.134 100.59 ;
      RECT MASK 2 61.348 99.54 61.408 100.59 ;
      RECT MASK 2 61.622 99.54 61.682 100.59 ;
      RECT MASK 2 61.896 99.54 61.956 100.59 ;
      RECT MASK 2 62.17 99.54 62.23 100.59 ;
      RECT MASK 2 62.444 99.54 62.504 100.59 ;
      RECT MASK 2 62.718 99.54 62.778 100.59 ;
      RECT MASK 2 62.992 99.54 63.052 100.59 ;
      RECT MASK 2 63.266 99.54 63.326 100.59 ;
      RECT MASK 2 63.54 99.54 63.6 100.59 ;
      RECT MASK 2 63.814 99.54 63.874 100.59 ;
      RECT MASK 2 64.088 99.54 64.148 100.59 ;
      RECT MASK 2 64.362 99.54 64.422 100.59 ;
      RECT MASK 2 64.636 99.54 64.696 100.59 ;
      RECT MASK 2 64.91 99.54 64.97 100.59 ;
      RECT MASK 2 65.184 99.54 65.244 100.59 ;
      RECT MASK 2 65.458 99.54 65.518 100.59 ;
      RECT MASK 2 65.732 99.54 65.792 100.59 ;
      RECT MASK 2 66.006 99.54 66.066 100.59 ;
      RECT MASK 2 66.28 99.54 66.34 100.59 ;
      RECT MASK 2 66.554 99.54 66.614 100.59 ;
      RECT MASK 2 66.828 99.54 66.888 100.59 ;
      RECT MASK 2 67.102 99.54 67.162 100.59 ;
      RECT MASK 2 67.376 99.54 67.436 100.59 ;
      RECT MASK 2 67.65 99.54 67.71 100.59 ;
      RECT MASK 2 67.924 99.54 67.984 100.59 ;
      RECT MASK 2 68.198 99.54 68.258 100.59 ;
      RECT MASK 2 68.472 99.54 68.532 100.59 ;
      RECT MASK 2 68.746 99.54 68.806 100.59 ;
      RECT MASK 2 69.02 99.54 69.08 100.59 ;
      RECT MASK 2 69.294 99.54 69.354 100.59 ;
      RECT MASK 2 69.568 99.54 69.628 100.59 ;
      RECT MASK 2 69.842 99.54 69.902 100.59 ;
      RECT MASK 2 70.116 99.54 70.176 100.59 ;
      RECT MASK 2 70.39 99.54 70.45 100.59 ;
      RECT MASK 2 70.664 99.54 70.724 100.59 ;
      RECT MASK 2 70.938 99.54 70.998 100.59 ;
      RECT MASK 2 71.212 99.54 71.272 100.59 ;
      RECT MASK 2 71.486 99.54 71.546 100.59 ;
      RECT MASK 2 71.76 99.54 71.82 100.59 ;
      RECT MASK 2 72.034 99.54 72.094 100.59 ;
      RECT MASK 2 72.308 99.54 72.368 100.59 ;
      RECT MASK 2 72.582 99.54 72.642 100.59 ;
      RECT MASK 2 72.856 99.54 72.916 100.59 ;
      RECT MASK 2 73.13 99.54 73.19 100.59 ;
      RECT MASK 2 73.404 99.54 73.464 100.59 ;
      RECT MASK 2 73.678 99.54 73.738 100.59 ;
      RECT MASK 2 73.952 99.54 74.012 100.59 ;
      RECT MASK 2 74.226 99.54 74.286 100.59 ;
      RECT MASK 2 74.5 99.54 74.56 100.59 ;
      RECT MASK 2 74.774 99.54 74.834 100.59 ;
      RECT MASK 2 75.048 99.54 75.108 100.59 ;
      RECT MASK 2 75.322 99.54 75.382 100.59 ;
      RECT MASK 2 75.596 99.54 75.656 100.59 ;
      RECT MASK 2 75.87 99.54 75.93 100.59 ;
      RECT MASK 2 76.144 99.54 76.204 100.59 ;
      RECT MASK 2 76.418 99.54 76.478 100.59 ;
      RECT MASK 2 76.692 99.54 76.752 100.59 ;
      RECT MASK 2 76.966 99.54 77.026 100.59 ;
      RECT MASK 2 77.24 99.54 77.3 100.59 ;
      RECT MASK 2 77.514 99.54 77.574 100.59 ;
      RECT MASK 2 77.788 99.54 77.848 100.59 ;
      RECT MASK 2 78.062 99.54 78.122 100.59 ;
      RECT MASK 2 78.336 99.54 78.396 100.59 ;
      RECT MASK 2 78.61 99.54 78.67 100.59 ;
      RECT MASK 2 78.884 99.54 78.944 100.59 ;
      RECT MASK 2 79.158 99.54 79.218 100.59 ;
      RECT MASK 2 79.432 99.54 79.492 100.59 ;
      RECT MASK 2 79.706 99.54 79.766 100.59 ;
      RECT MASK 2 79.98 99.54 80.04 100.59 ;
      RECT MASK 2 80.254 99.54 80.314 100.59 ;
      RECT MASK 2 80.528 99.54 80.588 100.59 ;
      RECT MASK 2 80.802 99.54 80.862 100.59 ;
      RECT MASK 2 81.076 99.54 81.136 100.59 ;
      RECT MASK 2 81.35 99.54 81.41 100.59 ;
      RECT MASK 2 81.624 99.54 81.684 100.59 ;
      RECT MASK 2 81.898 99.54 81.958 100.59 ;
      RECT MASK 2 82.172 99.54 82.232 100.59 ;
      RECT MASK 2 82.446 99.54 82.506 100.59 ;
      RECT MASK 2 82.72 99.54 82.78 100.59 ;
      RECT MASK 2 82.994 99.54 83.054 100.59 ;
      RECT MASK 2 83.268 99.54 83.328 100.59 ;
      RECT MASK 2 83.542 99.54 83.602 100.59 ;
      RECT MASK 2 83.816 99.54 83.876 100.59 ;
      RECT MASK 2 84.09 99.54 84.15 100.59 ;
      RECT MASK 2 84.364 99.54 84.424 100.59 ;
      RECT MASK 2 84.638 99.54 84.698 100.59 ;
      RECT MASK 2 84.912 99.54 84.972 100.59 ;
      RECT MASK 2 85.186 99.54 85.246 100.59 ;
      RECT MASK 2 85.46 99.54 85.52 100.59 ;
      RECT MASK 2 85.734 99.54 85.794 100.59 ;
      RECT MASK 2 86.008 99.54 86.068 100.59 ;
      RECT MASK 2 86.282 99.54 86.342 100.59 ;
      RECT MASK 2 86.556 99.54 86.616 100.59 ;
      RECT MASK 2 86.83 99.54 86.89 100.59 ;
      RECT MASK 2 89.089 99.54 89.149 100.59 ;
      RECT MASK 2 89.363 99.54 89.423 100.59 ;
      RECT MASK 2 89.637 99.54 89.697 100.59 ;
      RECT MASK 2 89.911 99.54 89.971 100.59 ;
      RECT MASK 2 90.185 99.54 90.245 100.59 ;
      RECT MASK 2 90.459 99.54 90.519 100.59 ;
      RECT MASK 2 90.733 99.54 90.793 100.59 ;
      RECT MASK 2 91.007 99.54 91.067 100.59 ;
      RECT MASK 2 91.281 99.54 91.341 100.59 ;
      RECT MASK 2 91.555 99.54 91.615 100.59 ;
      RECT MASK 2 91.829 99.54 91.889 100.59 ;
      RECT MASK 2 92.103 99.54 92.163 100.59 ;
      RECT MASK 2 92.377 99.54 92.437 100.59 ;
      RECT MASK 2 92.651 99.54 92.711 100.59 ;
      RECT MASK 2 92.925 99.54 92.985 100.59 ;
      RECT MASK 2 93.199 99.54 93.259 100.59 ;
      RECT MASK 2 93.473 99.54 93.533 100.59 ;
      RECT MASK 2 93.747 99.54 93.807 100.59 ;
      RECT MASK 2 94.021 99.54 94.081 100.59 ;
      RECT MASK 2 94.295 99.54 94.355 100.59 ;
      RECT MASK 2 94.569 99.54 94.629 100.59 ;
      RECT MASK 2 94.843 99.54 94.903 100.59 ;
      RECT MASK 2 95.117 99.54 95.177 100.59 ;
      RECT MASK 2 95.391 99.54 95.451 100.59 ;
      RECT MASK 2 95.665 99.54 95.725 100.59 ;
      RECT MASK 2 95.939 99.54 95.999 100.59 ;
      RECT MASK 2 96.213 99.54 96.273 100.59 ;
      RECT MASK 2 96.487 99.54 96.547 100.59 ;
      RECT MASK 2 96.761 99.54 96.821 100.59 ;
      RECT MASK 2 97.035 99.54 97.095 100.59 ;
      RECT MASK 2 97.309 99.54 97.369 100.59 ;
      RECT MASK 2 97.583 99.54 97.643 100.59 ;
      RECT MASK 2 97.857 99.54 97.917 100.59 ;
      RECT MASK 2 98.131 99.54 98.191 100.59 ;
      RECT MASK 2 98.405 99.54 98.465 100.59 ;
      RECT MASK 2 98.679 99.54 98.739 100.59 ;
      RECT MASK 2 98.953 99.54 99.013 100.59 ;
      RECT MASK 2 99.227 99.54 99.287 100.59 ;
      RECT MASK 2 99.501 99.54 99.561 100.59 ;
      RECT MASK 2 99.775 99.54 99.835 100.59 ;
      RECT MASK 2 100.049 99.54 100.109 100.59 ;
      RECT MASK 2 100.323 99.54 100.383 100.59 ;
      RECT MASK 2 100.597 99.54 100.657 100.59 ;
      RECT MASK 2 100.871 99.54 100.931 100.59 ;
      RECT MASK 2 101.145 99.54 101.205 100.59 ;
      RECT MASK 2 101.419 99.54 101.479 100.59 ;
      RECT MASK 2 101.693 99.54 101.753 100.59 ;
      RECT MASK 2 101.967 99.54 102.027 100.59 ;
      RECT MASK 2 102.241 99.54 102.301 100.59 ;
      RECT MASK 2 102.515 99.54 102.575 100.59 ;
      RECT MASK 2 102.789 99.54 102.849 100.59 ;
      RECT MASK 2 103.063 99.54 103.123 100.59 ;
      RECT MASK 2 103.337 99.54 103.397 100.59 ;
      RECT MASK 2 103.611 99.54 103.671 100.59 ;
      RECT MASK 2 103.885 99.54 103.945 100.59 ;
      RECT MASK 2 104.159 99.54 104.219 100.59 ;
      RECT MASK 2 104.433 99.54 104.493 100.59 ;
      RECT MASK 2 104.707 99.54 104.767 100.59 ;
      RECT MASK 2 104.981 99.54 105.041 100.59 ;
      RECT MASK 2 105.255 99.54 105.315 100.59 ;
      RECT MASK 2 105.529 99.54 105.589 100.59 ;
      RECT MASK 2 105.803 99.54 105.863 100.59 ;
      RECT MASK 2 106.077 99.54 106.137 100.59 ;
      RECT MASK 2 106.351 99.54 106.411 100.59 ;
      RECT MASK 2 106.625 99.54 106.685 100.59 ;
      RECT MASK 2 106.899 99.54 106.959 100.59 ;
      RECT MASK 2 107.173 99.54 107.233 100.59 ;
      RECT MASK 2 107.447 99.54 107.507 100.59 ;
      RECT MASK 2 107.721 99.54 107.781 100.59 ;
      RECT MASK 2 107.995 99.54 108.055 100.59 ;
      RECT MASK 2 108.269 99.54 108.329 100.59 ;
      RECT MASK 2 108.543 99.54 108.603 100.59 ;
      RECT MASK 2 108.817 99.54 108.877 100.59 ;
      RECT MASK 2 109.091 99.54 109.151 100.59 ;
      RECT MASK 2 109.365 99.54 109.425 100.59 ;
      RECT MASK 2 109.639 99.54 109.699 100.59 ;
      RECT MASK 2 109.913 99.54 109.973 100.59 ;
      RECT MASK 2 110.187 99.54 110.247 100.59 ;
      RECT MASK 2 110.461 99.54 110.521 100.59 ;
      RECT MASK 2 110.735 99.54 110.795 100.59 ;
      RECT MASK 2 111.009 99.54 111.069 100.59 ;
      RECT MASK 2 111.283 99.54 111.343 100.59 ;
      RECT MASK 2 111.557 99.54 111.617 100.59 ;
      RECT MASK 2 111.831 99.54 111.891 100.59 ;
      RECT MASK 2 112.105 99.54 112.165 100.59 ;
      RECT MASK 2 112.379 99.54 112.439 100.59 ;
      RECT MASK 2 112.653 99.54 112.713 100.59 ;
      RECT MASK 2 112.927 99.54 112.987 100.59 ;
      RECT MASK 2 113.201 99.54 113.261 100.59 ;
      RECT MASK 2 113.475 99.54 113.535 100.59 ;
      RECT MASK 2 113.749 99.54 113.809 100.59 ;
      RECT MASK 2 114.023 99.54 114.083 100.59 ;
      RECT MASK 2 114.297 99.54 114.357 100.59 ;
      RECT MASK 2 114.571 99.54 114.631 100.59 ;
      RECT MASK 2 114.845 99.54 114.905 100.59 ;
      RECT MASK 2 115.119 99.54 115.179 100.59 ;
      RECT MASK 2 115.393 99.54 115.453 100.59 ;
      RECT MASK 2 115.667 99.54 115.727 100.59 ;
      RECT MASK 2 115.941 99.54 116.001 100.59 ;
      RECT MASK 2 116.215 99.54 116.275 100.59 ;
      RECT MASK 2 116.489 99.54 116.549 100.59 ;
      RECT MASK 2 116.763 99.54 116.823 100.59 ;
      RECT MASK 2 117.037 99.54 117.097 100.59 ;
      RECT MASK 2 117.311 99.54 117.371 100.59 ;
      RECT MASK 2 117.585 99.54 117.645 100.59 ;
      RECT MASK 2 117.859 99.54 117.919 100.59 ;
      RECT MASK 2 118.133 99.54 118.193 100.59 ;
      RECT MASK 2 118.407 99.54 118.467 100.59 ;
      RECT MASK 2 118.681 99.54 118.741 100.59 ;
      RECT MASK 2 118.955 99.54 119.015 100.59 ;
      RECT MASK 2 119.229 99.54 119.289 100.59 ;
      RECT MASK 2 119.503 99.54 119.563 100.59 ;
      RECT MASK 2 119.777 99.54 119.837 100.59 ;
      RECT MASK 2 120.051 99.54 120.111 100.59 ;
      RECT MASK 2 120.325 99.54 120.385 100.59 ;
      RECT MASK 2 120.599 99.54 120.659 100.59 ;
      RECT MASK 2 120.873 99.54 120.933 100.59 ;
      RECT MASK 2 121.147 99.54 121.207 100.59 ;
      RECT MASK 2 121.421 99.54 121.481 100.59 ;
      RECT MASK 2 121.695 99.54 121.755 100.59 ;
      RECT MASK 2 121.969 99.54 122.029 100.59 ;
      RECT MASK 2 122.243 99.54 122.303 100.59 ;
      RECT MASK 2 122.517 99.54 122.577 100.59 ;
      RECT MASK 2 122.791 99.54 122.851 100.59 ;
      RECT MASK 2 123.065 99.54 123.125 100.59 ;
      RECT MASK 2 123.339 99.54 123.399 100.59 ;
      RECT MASK 2 123.613 99.54 123.673 100.59 ;
      RECT MASK 2 123.887 99.54 123.947 100.59 ;
      RECT MASK 2 124.161 99.54 124.221 100.59 ;
      RECT MASK 2 124.435 99.54 124.495 100.59 ;
      RECT MASK 2 124.709 99.54 124.769 100.59 ;
      RECT MASK 2 124.983 99.54 125.043 100.59 ;
      RECT MASK 2 125.257 99.54 125.317 100.59 ;
      RECT MASK 2 125.531 99.54 125.591 100.59 ;
      RECT MASK 2 125.805 99.54 125.865 100.59 ;
      RECT MASK 2 126.079 99.54 126.139 100.59 ;
      RECT MASK 2 126.353 99.54 126.413 100.59 ;
      RECT MASK 2 126.627 99.54 126.687 100.59 ;
      RECT MASK 2 126.901 99.54 126.961 100.59 ;
      RECT MASK 2 127.175 99.54 127.235 100.59 ;
      RECT MASK 2 127.449 99.54 127.509 100.59 ;
      RECT MASK 2 2.338 101.25 2.398 102.3 ;
      RECT MASK 2 2.612 101.25 2.672 102.3 ;
      RECT MASK 2 2.886 101.25 2.946 102.3 ;
      RECT MASK 2 3.16 101.25 3.22 102.3 ;
      RECT MASK 2 3.434 101.25 3.494 102.3 ;
      RECT MASK 2 3.708 101.25 3.768 102.3 ;
      RECT MASK 2 3.982 101.25 4.042 102.3 ;
      RECT MASK 2 4.256 101.25 4.316 102.3 ;
      RECT MASK 2 4.53 101.25 4.59 102.3 ;
      RECT MASK 2 4.804 101.25 4.864 102.3 ;
      RECT MASK 2 5.078 101.25 5.138 102.3 ;
      RECT MASK 2 5.352 101.25 5.412 102.3 ;
      RECT MASK 2 5.626 101.25 5.686 102.3 ;
      RECT MASK 2 5.9 101.25 5.96 102.3 ;
      RECT MASK 2 6.174 101.25 6.234 102.3 ;
      RECT MASK 2 6.448 101.25 6.508 102.3 ;
      RECT MASK 2 6.722 101.25 6.782 102.3 ;
      RECT MASK 2 6.996 101.25 7.056 102.3 ;
      RECT MASK 2 7.27 101.25 7.33 102.3 ;
      RECT MASK 2 7.544 101.25 7.604 102.3 ;
      RECT MASK 2 7.818 101.25 7.878 102.3 ;
      RECT MASK 2 8.092 101.25 8.152 102.3 ;
      RECT MASK 2 8.366 101.25 8.426 102.3 ;
      RECT MASK 2 8.64 101.25 8.7 102.3 ;
      RECT MASK 2 8.914 101.25 8.974 102.3 ;
      RECT MASK 2 9.188 101.25 9.248 102.3 ;
      RECT MASK 2 9.462 101.25 9.522 102.3 ;
      RECT MASK 2 9.736 101.25 9.796 102.3 ;
      RECT MASK 2 10.01 101.25 10.07 102.3 ;
      RECT MASK 2 10.284 101.25 10.344 102.3 ;
      RECT MASK 2 10.558 101.25 10.618 102.3 ;
      RECT MASK 2 10.832 101.25 10.892 102.3 ;
      RECT MASK 2 11.106 101.25 11.166 102.3 ;
      RECT MASK 2 11.38 101.25 11.44 102.3 ;
      RECT MASK 2 11.654 101.25 11.714 102.3 ;
      RECT MASK 2 11.928 101.25 11.988 102.3 ;
      RECT MASK 2 12.202 101.25 12.262 102.3 ;
      RECT MASK 2 12.476 101.25 12.536 102.3 ;
      RECT MASK 2 12.75 101.25 12.81 102.3 ;
      RECT MASK 2 13.024 101.25 13.084 102.3 ;
      RECT MASK 2 13.298 101.25 13.358 102.3 ;
      RECT MASK 2 13.572 101.25 13.632 102.3 ;
      RECT MASK 2 13.846 101.25 13.906 102.3 ;
      RECT MASK 2 14.12 101.25 14.18 102.3 ;
      RECT MASK 2 14.394 101.25 14.454 102.3 ;
      RECT MASK 2 14.668 101.25 14.728 102.3 ;
      RECT MASK 2 14.942 101.25 15.002 102.3 ;
      RECT MASK 2 15.216 101.25 15.276 102.3 ;
      RECT MASK 2 15.49 101.25 15.55 102.3 ;
      RECT MASK 2 15.764 101.25 15.824 102.3 ;
      RECT MASK 2 16.038 101.25 16.098 102.3 ;
      RECT MASK 2 16.312 101.25 16.372 102.3 ;
      RECT MASK 2 16.586 101.25 16.646 102.3 ;
      RECT MASK 2 16.86 101.25 16.92 102.3 ;
      RECT MASK 2 17.134 101.25 17.194 102.3 ;
      RECT MASK 2 17.408 101.25 17.468 102.3 ;
      RECT MASK 2 17.682 101.25 17.742 102.3 ;
      RECT MASK 2 17.956 101.25 18.016 102.3 ;
      RECT MASK 2 18.23 101.25 18.29 102.3 ;
      RECT MASK 2 18.504 101.25 18.564 102.3 ;
      RECT MASK 2 18.778 101.25 18.838 102.3 ;
      RECT MASK 2 19.052 101.25 19.112 102.3 ;
      RECT MASK 2 19.326 101.25 19.386 102.3 ;
      RECT MASK 2 19.6 101.25 19.66 102.3 ;
      RECT MASK 2 19.874 101.25 19.934 102.3 ;
      RECT MASK 2 20.148 101.25 20.208 102.3 ;
      RECT MASK 2 20.422 101.25 20.482 102.3 ;
      RECT MASK 2 20.696 101.25 20.756 102.3 ;
      RECT MASK 2 20.97 101.25 21.03 102.3 ;
      RECT MASK 2 21.244 101.25 21.304 102.3 ;
      RECT MASK 2 21.518 101.25 21.578 102.3 ;
      RECT MASK 2 21.792 101.25 21.852 102.3 ;
      RECT MASK 2 22.066 101.25 22.126 102.3 ;
      RECT MASK 2 22.34 101.25 22.4 102.3 ;
      RECT MASK 2 22.614 101.25 22.674 102.3 ;
      RECT MASK 2 22.888 101.25 22.948 102.3 ;
      RECT MASK 2 23.162 101.25 23.222 102.3 ;
      RECT MASK 2 23.436 101.25 23.496 102.3 ;
      RECT MASK 2 23.71 101.25 23.77 102.3 ;
      RECT MASK 2 23.984 101.25 24.044 102.3 ;
      RECT MASK 2 24.258 101.25 24.318 102.3 ;
      RECT MASK 2 24.532 101.25 24.592 102.3 ;
      RECT MASK 2 24.806 101.25 24.866 102.3 ;
      RECT MASK 2 25.08 101.25 25.14 102.3 ;
      RECT MASK 2 25.354 101.25 25.414 102.3 ;
      RECT MASK 2 25.628 101.25 25.688 102.3 ;
      RECT MASK 2 25.902 101.25 25.962 102.3 ;
      RECT MASK 2 26.176 101.25 26.236 102.3 ;
      RECT MASK 2 26.45 101.25 26.51 102.3 ;
      RECT MASK 2 26.724 101.25 26.784 102.3 ;
      RECT MASK 2 26.998 101.25 27.058 102.3 ;
      RECT MASK 2 27.272 101.25 27.332 102.3 ;
      RECT MASK 2 27.546 101.25 27.606 102.3 ;
      RECT MASK 2 27.82 101.25 27.88 102.3 ;
      RECT MASK 2 28.094 101.25 28.154 102.3 ;
      RECT MASK 2 28.368 101.25 28.428 102.3 ;
      RECT MASK 2 28.642 101.25 28.702 102.3 ;
      RECT MASK 2 28.916 101.25 28.976 102.3 ;
      RECT MASK 2 29.19 101.25 29.25 102.3 ;
      RECT MASK 2 29.464 101.25 29.524 102.3 ;
      RECT MASK 2 29.738 101.25 29.798 102.3 ;
      RECT MASK 2 30.012 101.25 30.072 102.3 ;
      RECT MASK 2 30.286 101.25 30.346 102.3 ;
      RECT MASK 2 30.56 101.25 30.62 102.3 ;
      RECT MASK 2 30.834 101.25 30.894 102.3 ;
      RECT MASK 2 31.108 101.25 31.168 102.3 ;
      RECT MASK 2 31.382 101.25 31.442 102.3 ;
      RECT MASK 2 31.656 101.25 31.716 102.3 ;
      RECT MASK 2 31.93 101.25 31.99 102.3 ;
      RECT MASK 2 32.204 101.25 32.264 102.3 ;
      RECT MASK 2 32.478 101.25 32.538 102.3 ;
      RECT MASK 2 32.752 101.25 32.812 102.3 ;
      RECT MASK 2 33.026 101.25 33.086 102.3 ;
      RECT MASK 2 33.3 101.25 33.36 102.3 ;
      RECT MASK 2 33.574 101.25 33.634 102.3 ;
      RECT MASK 2 33.848 101.25 33.908 102.3 ;
      RECT MASK 2 34.122 101.25 34.182 102.3 ;
      RECT MASK 2 34.396 101.25 34.456 102.3 ;
      RECT MASK 2 34.67 101.25 34.73 102.3 ;
      RECT MASK 2 34.944 101.25 35.004 102.3 ;
      RECT MASK 2 35.218 101.25 35.278 102.3 ;
      RECT MASK 2 35.492 101.25 35.552 102.3 ;
      RECT MASK 2 35.766 101.25 35.826 102.3 ;
      RECT MASK 2 36.04 101.25 36.1 102.3 ;
      RECT MASK 2 36.314 101.25 36.374 102.3 ;
      RECT MASK 2 36.588 101.25 36.648 102.3 ;
      RECT MASK 2 36.862 101.25 36.922 102.3 ;
      RECT MASK 2 37.136 101.25 37.196 102.3 ;
      RECT MASK 2 37.41 101.25 37.47 102.3 ;
      RECT MASK 2 37.684 101.25 37.744 102.3 ;
      RECT MASK 2 37.958 101.25 38.018 102.3 ;
      RECT MASK 2 38.232 101.25 38.292 102.3 ;
      RECT MASK 2 38.506 101.25 38.566 102.3 ;
      RECT MASK 2 38.78 101.25 38.84 102.3 ;
      RECT MASK 2 39.054 101.25 39.114 102.3 ;
      RECT MASK 2 39.328 101.25 39.388 102.3 ;
      RECT MASK 2 39.602 101.25 39.662 102.3 ;
      RECT MASK 2 39.876 101.25 39.936 102.3 ;
      RECT MASK 2 40.15 101.25 40.21 102.3 ;
      RECT MASK 2 40.424 101.25 40.484 102.3 ;
      RECT MASK 2 40.698 101.25 40.758 102.3 ;
      RECT MASK 2 40.972 101.25 41.032 102.3 ;
      RECT MASK 2 41.246 101.25 41.306 102.3 ;
      RECT MASK 2 41.52 101.25 41.58 102.3 ;
      RECT MASK 2 41.794 101.25 41.854 102.3 ;
      RECT MASK 2 42.068 101.25 42.128 102.3 ;
      RECT MASK 2 42.342 101.25 42.402 102.3 ;
      RECT MASK 2 42.616 101.25 42.676 102.3 ;
      RECT MASK 2 42.89 101.25 42.95 102.3 ;
      RECT MASK 2 43.164 101.25 43.224 102.3 ;
      RECT MASK 2 43.438 101.25 43.498 102.3 ;
      RECT MASK 2 45.73 101.25 45.79 102.3 ;
      RECT MASK 2 46.004 101.25 46.064 102.3 ;
      RECT MASK 2 46.278 101.25 46.338 102.3 ;
      RECT MASK 2 46.552 101.25 46.612 102.3 ;
      RECT MASK 2 46.826 101.25 46.886 102.3 ;
      RECT MASK 2 47.1 101.25 47.16 102.3 ;
      RECT MASK 2 47.374 101.25 47.434 102.3 ;
      RECT MASK 2 47.648 101.25 47.708 102.3 ;
      RECT MASK 2 47.922 101.25 47.982 102.3 ;
      RECT MASK 2 48.196 101.25 48.256 102.3 ;
      RECT MASK 2 48.47 101.25 48.53 102.3 ;
      RECT MASK 2 48.744 101.25 48.804 102.3 ;
      RECT MASK 2 49.018 101.25 49.078 102.3 ;
      RECT MASK 2 49.292 101.25 49.352 102.3 ;
      RECT MASK 2 49.566 101.25 49.626 102.3 ;
      RECT MASK 2 49.84 101.25 49.9 102.3 ;
      RECT MASK 2 50.114 101.25 50.174 102.3 ;
      RECT MASK 2 50.388 101.25 50.448 102.3 ;
      RECT MASK 2 50.662 101.25 50.722 102.3 ;
      RECT MASK 2 50.936 101.25 50.996 102.3 ;
      RECT MASK 2 51.21 101.25 51.27 102.3 ;
      RECT MASK 2 51.484 101.25 51.544 102.3 ;
      RECT MASK 2 51.758 101.25 51.818 102.3 ;
      RECT MASK 2 52.032 101.25 52.092 102.3 ;
      RECT MASK 2 52.306 101.25 52.366 102.3 ;
      RECT MASK 2 52.58 101.25 52.64 102.3 ;
      RECT MASK 2 52.854 101.25 52.914 102.3 ;
      RECT MASK 2 53.128 101.25 53.188 102.3 ;
      RECT MASK 2 53.402 101.25 53.462 102.3 ;
      RECT MASK 2 53.676 101.25 53.736 102.3 ;
      RECT MASK 2 53.95 101.25 54.01 102.3 ;
      RECT MASK 2 54.224 101.25 54.284 102.3 ;
      RECT MASK 2 54.498 101.25 54.558 102.3 ;
      RECT MASK 2 54.772 101.25 54.832 102.3 ;
      RECT MASK 2 55.046 101.25 55.106 102.3 ;
      RECT MASK 2 55.32 101.25 55.38 102.3 ;
      RECT MASK 2 55.594 101.25 55.654 102.3 ;
      RECT MASK 2 55.868 101.25 55.928 102.3 ;
      RECT MASK 2 56.142 101.25 56.202 102.3 ;
      RECT MASK 2 56.416 101.25 56.476 102.3 ;
      RECT MASK 2 56.69 101.25 56.75 102.3 ;
      RECT MASK 2 56.964 101.25 57.024 102.3 ;
      RECT MASK 2 57.238 101.25 57.298 102.3 ;
      RECT MASK 2 57.512 101.25 57.572 102.3 ;
      RECT MASK 2 57.786 101.25 57.846 102.3 ;
      RECT MASK 2 58.06 101.25 58.12 102.3 ;
      RECT MASK 2 58.334 101.25 58.394 102.3 ;
      RECT MASK 2 58.608 101.25 58.668 102.3 ;
      RECT MASK 2 58.882 101.25 58.942 102.3 ;
      RECT MASK 2 59.156 101.25 59.216 102.3 ;
      RECT MASK 2 59.43 101.25 59.49 102.3 ;
      RECT MASK 2 59.704 101.25 59.764 102.3 ;
      RECT MASK 2 59.978 101.25 60.038 102.3 ;
      RECT MASK 2 60.252 101.25 60.312 102.3 ;
      RECT MASK 2 60.526 101.25 60.586 102.3 ;
      RECT MASK 2 60.8 101.25 60.86 102.3 ;
      RECT MASK 2 61.074 101.25 61.134 102.3 ;
      RECT MASK 2 61.348 101.25 61.408 102.3 ;
      RECT MASK 2 61.622 101.25 61.682 102.3 ;
      RECT MASK 2 61.896 101.25 61.956 102.3 ;
      RECT MASK 2 62.17 101.25 62.23 102.3 ;
      RECT MASK 2 62.444 101.25 62.504 102.3 ;
      RECT MASK 2 62.718 101.25 62.778 102.3 ;
      RECT MASK 2 62.992 101.25 63.052 102.3 ;
      RECT MASK 2 63.266 101.25 63.326 102.3 ;
      RECT MASK 2 63.54 101.25 63.6 102.3 ;
      RECT MASK 2 63.814 101.25 63.874 102.3 ;
      RECT MASK 2 64.088 101.25 64.148 102.3 ;
      RECT MASK 2 64.362 101.25 64.422 102.3 ;
      RECT MASK 2 64.636 101.25 64.696 102.3 ;
      RECT MASK 2 64.91 101.25 64.97 102.3 ;
      RECT MASK 2 65.184 101.25 65.244 102.3 ;
      RECT MASK 2 65.458 101.25 65.518 102.3 ;
      RECT MASK 2 65.732 101.25 65.792 102.3 ;
      RECT MASK 2 66.006 101.25 66.066 102.3 ;
      RECT MASK 2 66.28 101.25 66.34 102.3 ;
      RECT MASK 2 66.554 101.25 66.614 102.3 ;
      RECT MASK 2 66.828 101.25 66.888 102.3 ;
      RECT MASK 2 67.102 101.25 67.162 102.3 ;
      RECT MASK 2 67.376 101.25 67.436 102.3 ;
      RECT MASK 2 67.65 101.25 67.71 102.3 ;
      RECT MASK 2 67.924 101.25 67.984 102.3 ;
      RECT MASK 2 68.198 101.25 68.258 102.3 ;
      RECT MASK 2 68.472 101.25 68.532 102.3 ;
      RECT MASK 2 68.746 101.25 68.806 102.3 ;
      RECT MASK 2 69.02 101.25 69.08 102.3 ;
      RECT MASK 2 69.294 101.25 69.354 102.3 ;
      RECT MASK 2 69.568 101.25 69.628 102.3 ;
      RECT MASK 2 69.842 101.25 69.902 102.3 ;
      RECT MASK 2 70.116 101.25 70.176 102.3 ;
      RECT MASK 2 70.39 101.25 70.45 102.3 ;
      RECT MASK 2 70.664 101.25 70.724 102.3 ;
      RECT MASK 2 70.938 101.25 70.998 102.3 ;
      RECT MASK 2 71.212 101.25 71.272 102.3 ;
      RECT MASK 2 71.486 101.25 71.546 102.3 ;
      RECT MASK 2 71.76 101.25 71.82 102.3 ;
      RECT MASK 2 72.034 101.25 72.094 102.3 ;
      RECT MASK 2 72.308 101.25 72.368 102.3 ;
      RECT MASK 2 72.582 101.25 72.642 102.3 ;
      RECT MASK 2 72.856 101.25 72.916 102.3 ;
      RECT MASK 2 73.13 101.25 73.19 102.3 ;
      RECT MASK 2 73.404 101.25 73.464 102.3 ;
      RECT MASK 2 73.678 101.25 73.738 102.3 ;
      RECT MASK 2 73.952 101.25 74.012 102.3 ;
      RECT MASK 2 74.226 101.25 74.286 102.3 ;
      RECT MASK 2 74.5 101.25 74.56 102.3 ;
      RECT MASK 2 74.774 101.25 74.834 102.3 ;
      RECT MASK 2 75.048 101.25 75.108 102.3 ;
      RECT MASK 2 75.322 101.25 75.382 102.3 ;
      RECT MASK 2 75.596 101.25 75.656 102.3 ;
      RECT MASK 2 75.87 101.25 75.93 102.3 ;
      RECT MASK 2 76.144 101.25 76.204 102.3 ;
      RECT MASK 2 76.418 101.25 76.478 102.3 ;
      RECT MASK 2 76.692 101.25 76.752 102.3 ;
      RECT MASK 2 76.966 101.25 77.026 102.3 ;
      RECT MASK 2 77.24 101.25 77.3 102.3 ;
      RECT MASK 2 77.514 101.25 77.574 102.3 ;
      RECT MASK 2 77.788 101.25 77.848 102.3 ;
      RECT MASK 2 78.062 101.25 78.122 102.3 ;
      RECT MASK 2 78.336 101.25 78.396 102.3 ;
      RECT MASK 2 78.61 101.25 78.67 102.3 ;
      RECT MASK 2 78.884 101.25 78.944 102.3 ;
      RECT MASK 2 79.158 101.25 79.218 102.3 ;
      RECT MASK 2 79.432 101.25 79.492 102.3 ;
      RECT MASK 2 79.706 101.25 79.766 102.3 ;
      RECT MASK 2 79.98 101.25 80.04 102.3 ;
      RECT MASK 2 80.254 101.25 80.314 102.3 ;
      RECT MASK 2 80.528 101.25 80.588 102.3 ;
      RECT MASK 2 80.802 101.25 80.862 102.3 ;
      RECT MASK 2 81.076 101.25 81.136 102.3 ;
      RECT MASK 2 81.35 101.25 81.41 102.3 ;
      RECT MASK 2 81.624 101.25 81.684 102.3 ;
      RECT MASK 2 81.898 101.25 81.958 102.3 ;
      RECT MASK 2 82.172 101.25 82.232 102.3 ;
      RECT MASK 2 82.446 101.25 82.506 102.3 ;
      RECT MASK 2 82.72 101.25 82.78 102.3 ;
      RECT MASK 2 82.994 101.25 83.054 102.3 ;
      RECT MASK 2 83.268 101.25 83.328 102.3 ;
      RECT MASK 2 83.542 101.25 83.602 102.3 ;
      RECT MASK 2 83.816 101.25 83.876 102.3 ;
      RECT MASK 2 84.09 101.25 84.15 102.3 ;
      RECT MASK 2 84.364 101.25 84.424 102.3 ;
      RECT MASK 2 84.638 101.25 84.698 102.3 ;
      RECT MASK 2 84.912 101.25 84.972 102.3 ;
      RECT MASK 2 85.186 101.25 85.246 102.3 ;
      RECT MASK 2 85.46 101.25 85.52 102.3 ;
      RECT MASK 2 85.734 101.25 85.794 102.3 ;
      RECT MASK 2 86.008 101.25 86.068 102.3 ;
      RECT MASK 2 86.282 101.25 86.342 102.3 ;
      RECT MASK 2 86.556 101.25 86.616 102.3 ;
      RECT MASK 2 86.83 101.25 86.89 102.3 ;
      RECT MASK 2 89.089 101.25 89.149 102.3 ;
      RECT MASK 2 89.363 101.25 89.423 102.3 ;
      RECT MASK 2 89.637 101.25 89.697 102.3 ;
      RECT MASK 2 89.911 101.25 89.971 102.3 ;
      RECT MASK 2 90.185 101.25 90.245 102.3 ;
      RECT MASK 2 90.459 101.25 90.519 102.3 ;
      RECT MASK 2 90.733 101.25 90.793 102.3 ;
      RECT MASK 2 91.007 101.25 91.067 102.3 ;
      RECT MASK 2 91.281 101.25 91.341 102.3 ;
      RECT MASK 2 91.555 101.25 91.615 102.3 ;
      RECT MASK 2 91.829 101.25 91.889 102.3 ;
      RECT MASK 2 92.103 101.25 92.163 102.3 ;
      RECT MASK 2 92.377 101.25 92.437 102.3 ;
      RECT MASK 2 92.651 101.25 92.711 102.3 ;
      RECT MASK 2 92.925 101.25 92.985 102.3 ;
      RECT MASK 2 93.199 101.25 93.259 102.3 ;
      RECT MASK 2 93.473 101.25 93.533 102.3 ;
      RECT MASK 2 93.747 101.25 93.807 102.3 ;
      RECT MASK 2 94.021 101.25 94.081 102.3 ;
      RECT MASK 2 94.295 101.25 94.355 102.3 ;
      RECT MASK 2 94.569 101.25 94.629 102.3 ;
      RECT MASK 2 94.843 101.25 94.903 102.3 ;
      RECT MASK 2 95.117 101.25 95.177 102.3 ;
      RECT MASK 2 95.391 101.25 95.451 102.3 ;
      RECT MASK 2 95.665 101.25 95.725 102.3 ;
      RECT MASK 2 95.939 101.25 95.999 102.3 ;
      RECT MASK 2 96.213 101.25 96.273 102.3 ;
      RECT MASK 2 96.487 101.25 96.547 102.3 ;
      RECT MASK 2 96.761 101.25 96.821 102.3 ;
      RECT MASK 2 97.035 101.25 97.095 102.3 ;
      RECT MASK 2 97.309 101.25 97.369 102.3 ;
      RECT MASK 2 97.583 101.25 97.643 102.3 ;
      RECT MASK 2 97.857 101.25 97.917 102.3 ;
      RECT MASK 2 98.131 101.25 98.191 102.3 ;
      RECT MASK 2 98.405 101.25 98.465 102.3 ;
      RECT MASK 2 98.679 101.25 98.739 102.3 ;
      RECT MASK 2 98.953 101.25 99.013 102.3 ;
      RECT MASK 2 99.227 101.25 99.287 102.3 ;
      RECT MASK 2 99.501 101.25 99.561 102.3 ;
      RECT MASK 2 99.775 101.25 99.835 102.3 ;
      RECT MASK 2 100.049 101.25 100.109 102.3 ;
      RECT MASK 2 100.323 101.25 100.383 102.3 ;
      RECT MASK 2 100.597 101.25 100.657 102.3 ;
      RECT MASK 2 100.871 101.25 100.931 102.3 ;
      RECT MASK 2 101.145 101.25 101.205 102.3 ;
      RECT MASK 2 101.419 101.25 101.479 102.3 ;
      RECT MASK 2 101.693 101.25 101.753 102.3 ;
      RECT MASK 2 101.967 101.25 102.027 102.3 ;
      RECT MASK 2 102.241 101.25 102.301 102.3 ;
      RECT MASK 2 102.515 101.25 102.575 102.3 ;
      RECT MASK 2 102.789 101.25 102.849 102.3 ;
      RECT MASK 2 103.063 101.25 103.123 102.3 ;
      RECT MASK 2 103.337 101.25 103.397 102.3 ;
      RECT MASK 2 103.611 101.25 103.671 102.3 ;
      RECT MASK 2 103.885 101.25 103.945 102.3 ;
      RECT MASK 2 104.159 101.25 104.219 102.3 ;
      RECT MASK 2 104.433 101.25 104.493 102.3 ;
      RECT MASK 2 104.707 101.25 104.767 102.3 ;
      RECT MASK 2 104.981 101.25 105.041 102.3 ;
      RECT MASK 2 105.255 101.25 105.315 102.3 ;
      RECT MASK 2 105.529 101.25 105.589 102.3 ;
      RECT MASK 2 105.803 101.25 105.863 102.3 ;
      RECT MASK 2 106.077 101.25 106.137 102.3 ;
      RECT MASK 2 106.351 101.25 106.411 102.3 ;
      RECT MASK 2 106.625 101.25 106.685 102.3 ;
      RECT MASK 2 106.899 101.25 106.959 102.3 ;
      RECT MASK 2 107.173 101.25 107.233 102.3 ;
      RECT MASK 2 107.447 101.25 107.507 102.3 ;
      RECT MASK 2 107.721 101.25 107.781 102.3 ;
      RECT MASK 2 107.995 101.25 108.055 102.3 ;
      RECT MASK 2 108.269 101.25 108.329 102.3 ;
      RECT MASK 2 108.543 101.25 108.603 102.3 ;
      RECT MASK 2 108.817 101.25 108.877 102.3 ;
      RECT MASK 2 109.091 101.25 109.151 102.3 ;
      RECT MASK 2 109.365 101.25 109.425 102.3 ;
      RECT MASK 2 109.639 101.25 109.699 102.3 ;
      RECT MASK 2 109.913 101.25 109.973 102.3 ;
      RECT MASK 2 110.187 101.25 110.247 102.3 ;
      RECT MASK 2 110.461 101.25 110.521 102.3 ;
      RECT MASK 2 110.735 101.25 110.795 102.3 ;
      RECT MASK 2 111.009 101.25 111.069 102.3 ;
      RECT MASK 2 111.283 101.25 111.343 102.3 ;
      RECT MASK 2 111.557 101.25 111.617 102.3 ;
      RECT MASK 2 111.831 101.25 111.891 102.3 ;
      RECT MASK 2 112.105 101.25 112.165 102.3 ;
      RECT MASK 2 112.379 101.25 112.439 102.3 ;
      RECT MASK 2 112.653 101.25 112.713 102.3 ;
      RECT MASK 2 112.927 101.25 112.987 102.3 ;
      RECT MASK 2 113.201 101.25 113.261 102.3 ;
      RECT MASK 2 113.475 101.25 113.535 102.3 ;
      RECT MASK 2 113.749 101.25 113.809 102.3 ;
      RECT MASK 2 114.023 101.25 114.083 102.3 ;
      RECT MASK 2 114.297 101.25 114.357 102.3 ;
      RECT MASK 2 114.571 101.25 114.631 102.3 ;
      RECT MASK 2 114.845 101.25 114.905 102.3 ;
      RECT MASK 2 115.119 101.25 115.179 102.3 ;
      RECT MASK 2 115.393 101.25 115.453 102.3 ;
      RECT MASK 2 115.667 101.25 115.727 102.3 ;
      RECT MASK 2 115.941 101.25 116.001 102.3 ;
      RECT MASK 2 116.215 101.25 116.275 102.3 ;
      RECT MASK 2 116.489 101.25 116.549 102.3 ;
      RECT MASK 2 116.763 101.25 116.823 102.3 ;
      RECT MASK 2 117.037 101.25 117.097 102.3 ;
      RECT MASK 2 117.311 101.25 117.371 102.3 ;
      RECT MASK 2 117.585 101.25 117.645 102.3 ;
      RECT MASK 2 117.859 101.25 117.919 102.3 ;
      RECT MASK 2 118.133 101.25 118.193 102.3 ;
      RECT MASK 2 118.407 101.25 118.467 102.3 ;
      RECT MASK 2 118.681 101.25 118.741 102.3 ;
      RECT MASK 2 118.955 101.25 119.015 102.3 ;
      RECT MASK 2 119.229 101.25 119.289 102.3 ;
      RECT MASK 2 119.503 101.25 119.563 102.3 ;
      RECT MASK 2 119.777 101.25 119.837 102.3 ;
      RECT MASK 2 120.051 101.25 120.111 102.3 ;
      RECT MASK 2 120.325 101.25 120.385 102.3 ;
      RECT MASK 2 120.599 101.25 120.659 102.3 ;
      RECT MASK 2 120.873 101.25 120.933 102.3 ;
      RECT MASK 2 121.147 101.25 121.207 102.3 ;
      RECT MASK 2 121.421 101.25 121.481 102.3 ;
      RECT MASK 2 121.695 101.25 121.755 102.3 ;
      RECT MASK 2 121.969 101.25 122.029 102.3 ;
      RECT MASK 2 122.243 101.25 122.303 102.3 ;
      RECT MASK 2 122.517 101.25 122.577 102.3 ;
      RECT MASK 2 122.791 101.25 122.851 102.3 ;
      RECT MASK 2 123.065 101.25 123.125 102.3 ;
      RECT MASK 2 123.339 101.25 123.399 102.3 ;
      RECT MASK 2 123.613 101.25 123.673 102.3 ;
      RECT MASK 2 123.887 101.25 123.947 102.3 ;
      RECT MASK 2 124.161 101.25 124.221 102.3 ;
      RECT MASK 2 124.435 101.25 124.495 102.3 ;
      RECT MASK 2 124.709 101.25 124.769 102.3 ;
      RECT MASK 2 124.983 101.25 125.043 102.3 ;
      RECT MASK 2 125.257 101.25 125.317 102.3 ;
      RECT MASK 2 125.531 101.25 125.591 102.3 ;
      RECT MASK 2 125.805 101.25 125.865 102.3 ;
      RECT MASK 2 126.079 101.25 126.139 102.3 ;
      RECT MASK 2 126.353 101.25 126.413 102.3 ;
      RECT MASK 2 126.627 101.25 126.687 102.3 ;
      RECT MASK 2 126.901 101.25 126.961 102.3 ;
      RECT MASK 2 127.175 101.25 127.235 102.3 ;
      RECT MASK 2 127.449 101.25 127.509 102.3 ;
      RECT MASK 2 2.338 102.96 2.398 104.01 ;
      RECT MASK 2 2.612 102.96 2.672 104.01 ;
      RECT MASK 2 2.886 102.96 2.946 104.01 ;
      RECT MASK 2 3.16 102.96 3.22 104.01 ;
      RECT MASK 2 3.434 102.96 3.494 104.01 ;
      RECT MASK 2 3.708 102.96 3.768 104.01 ;
      RECT MASK 2 3.982 102.96 4.042 104.01 ;
      RECT MASK 2 4.256 102.96 4.316 104.01 ;
      RECT MASK 2 4.53 102.96 4.59 104.01 ;
      RECT MASK 2 4.804 102.96 4.864 104.01 ;
      RECT MASK 2 5.078 102.96 5.138 104.01 ;
      RECT MASK 2 5.352 102.96 5.412 104.01 ;
      RECT MASK 2 5.626 102.96 5.686 104.01 ;
      RECT MASK 2 5.9 102.96 5.96 104.01 ;
      RECT MASK 2 6.174 102.96 6.234 104.01 ;
      RECT MASK 2 6.448 102.96 6.508 104.01 ;
      RECT MASK 2 6.722 102.96 6.782 104.01 ;
      RECT MASK 2 6.996 102.96 7.056 104.01 ;
      RECT MASK 2 7.27 102.96 7.33 104.01 ;
      RECT MASK 2 7.544 102.96 7.604 104.01 ;
      RECT MASK 2 7.818 102.96 7.878 104.01 ;
      RECT MASK 2 8.092 102.96 8.152 104.01 ;
      RECT MASK 2 8.366 102.96 8.426 104.01 ;
      RECT MASK 2 8.64 102.96 8.7 104.01 ;
      RECT MASK 2 8.914 102.96 8.974 104.01 ;
      RECT MASK 2 9.188 102.96 9.248 104.01 ;
      RECT MASK 2 9.462 102.96 9.522 104.01 ;
      RECT MASK 2 9.736 102.96 9.796 104.01 ;
      RECT MASK 2 10.01 102.96 10.07 104.01 ;
      RECT MASK 2 10.284 102.96 10.344 104.01 ;
      RECT MASK 2 10.558 102.96 10.618 104.01 ;
      RECT MASK 2 10.832 102.96 10.892 104.01 ;
      RECT MASK 2 11.106 102.96 11.166 104.01 ;
      RECT MASK 2 11.38 102.96 11.44 104.01 ;
      RECT MASK 2 11.654 102.96 11.714 104.01 ;
      RECT MASK 2 11.928 102.96 11.988 104.01 ;
      RECT MASK 2 12.202 102.96 12.262 104.01 ;
      RECT MASK 2 12.476 102.96 12.536 104.01 ;
      RECT MASK 2 12.75 102.96 12.81 104.01 ;
      RECT MASK 2 13.024 102.96 13.084 104.01 ;
      RECT MASK 2 13.298 102.96 13.358 104.01 ;
      RECT MASK 2 13.572 102.96 13.632 104.01 ;
      RECT MASK 2 13.846 102.96 13.906 104.01 ;
      RECT MASK 2 14.12 102.96 14.18 104.01 ;
      RECT MASK 2 14.394 102.96 14.454 104.01 ;
      RECT MASK 2 14.668 102.96 14.728 104.01 ;
      RECT MASK 2 14.942 102.96 15.002 104.01 ;
      RECT MASK 2 15.216 102.96 15.276 104.01 ;
      RECT MASK 2 15.49 102.96 15.55 104.01 ;
      RECT MASK 2 15.764 102.96 15.824 104.01 ;
      RECT MASK 2 16.038 102.96 16.098 104.01 ;
      RECT MASK 2 16.312 102.96 16.372 104.01 ;
      RECT MASK 2 16.586 102.96 16.646 104.01 ;
      RECT MASK 2 16.86 102.96 16.92 104.01 ;
      RECT MASK 2 17.134 102.96 17.194 104.01 ;
      RECT MASK 2 17.408 102.96 17.468 104.01 ;
      RECT MASK 2 17.682 102.96 17.742 104.01 ;
      RECT MASK 2 17.956 102.96 18.016 104.01 ;
      RECT MASK 2 18.23 102.96 18.29 104.01 ;
      RECT MASK 2 18.504 102.96 18.564 104.01 ;
      RECT MASK 2 18.778 102.96 18.838 104.01 ;
      RECT MASK 2 19.052 102.96 19.112 104.01 ;
      RECT MASK 2 19.326 102.96 19.386 104.01 ;
      RECT MASK 2 19.6 102.96 19.66 104.01 ;
      RECT MASK 2 19.874 102.96 19.934 104.01 ;
      RECT MASK 2 20.148 102.96 20.208 104.01 ;
      RECT MASK 2 20.422 102.96 20.482 104.01 ;
      RECT MASK 2 20.696 102.96 20.756 104.01 ;
      RECT MASK 2 20.97 102.96 21.03 104.01 ;
      RECT MASK 2 21.244 102.96 21.304 104.01 ;
      RECT MASK 2 21.518 102.96 21.578 104.01 ;
      RECT MASK 2 21.792 102.96 21.852 104.01 ;
      RECT MASK 2 22.066 102.96 22.126 104.01 ;
      RECT MASK 2 22.34 102.96 22.4 104.01 ;
      RECT MASK 2 22.614 102.96 22.674 104.01 ;
      RECT MASK 2 22.888 102.96 22.948 104.01 ;
      RECT MASK 2 23.162 102.96 23.222 104.01 ;
      RECT MASK 2 23.436 102.96 23.496 104.01 ;
      RECT MASK 2 23.71 102.96 23.77 104.01 ;
      RECT MASK 2 23.984 102.96 24.044 104.01 ;
      RECT MASK 2 24.258 102.96 24.318 104.01 ;
      RECT MASK 2 24.532 102.96 24.592 104.01 ;
      RECT MASK 2 24.806 102.96 24.866 104.01 ;
      RECT MASK 2 25.08 102.96 25.14 104.01 ;
      RECT MASK 2 25.354 102.96 25.414 104.01 ;
      RECT MASK 2 25.628 102.96 25.688 104.01 ;
      RECT MASK 2 25.902 102.96 25.962 104.01 ;
      RECT MASK 2 26.176 102.96 26.236 104.01 ;
      RECT MASK 2 26.45 102.96 26.51 104.01 ;
      RECT MASK 2 26.724 102.96 26.784 104.01 ;
      RECT MASK 2 26.998 102.96 27.058 104.01 ;
      RECT MASK 2 27.272 102.96 27.332 104.01 ;
      RECT MASK 2 27.546 102.96 27.606 104.01 ;
      RECT MASK 2 27.82 102.96 27.88 104.01 ;
      RECT MASK 2 28.094 102.96 28.154 104.01 ;
      RECT MASK 2 28.368 102.96 28.428 104.01 ;
      RECT MASK 2 28.642 102.96 28.702 104.01 ;
      RECT MASK 2 28.916 102.96 28.976 104.01 ;
      RECT MASK 2 29.19 102.96 29.25 104.01 ;
      RECT MASK 2 29.464 102.96 29.524 104.01 ;
      RECT MASK 2 29.738 102.96 29.798 104.01 ;
      RECT MASK 2 30.012 102.96 30.072 104.01 ;
      RECT MASK 2 30.286 102.96 30.346 104.01 ;
      RECT MASK 2 30.56 102.96 30.62 104.01 ;
      RECT MASK 2 30.834 102.96 30.894 104.01 ;
      RECT MASK 2 31.108 102.96 31.168 104.01 ;
      RECT MASK 2 31.382 102.96 31.442 104.01 ;
      RECT MASK 2 31.656 102.96 31.716 104.01 ;
      RECT MASK 2 31.93 102.96 31.99 104.01 ;
      RECT MASK 2 32.204 102.96 32.264 104.01 ;
      RECT MASK 2 32.478 102.96 32.538 104.01 ;
      RECT MASK 2 32.752 102.96 32.812 104.01 ;
      RECT MASK 2 33.026 102.96 33.086 104.01 ;
      RECT MASK 2 33.3 102.96 33.36 104.01 ;
      RECT MASK 2 33.574 102.96 33.634 104.01 ;
      RECT MASK 2 33.848 102.96 33.908 104.01 ;
      RECT MASK 2 34.122 102.96 34.182 104.01 ;
      RECT MASK 2 34.396 102.96 34.456 104.01 ;
      RECT MASK 2 34.67 102.96 34.73 104.01 ;
      RECT MASK 2 34.944 102.96 35.004 104.01 ;
      RECT MASK 2 35.218 102.96 35.278 104.01 ;
      RECT MASK 2 35.492 102.96 35.552 104.01 ;
      RECT MASK 2 35.766 102.96 35.826 104.01 ;
      RECT MASK 2 36.04 102.96 36.1 104.01 ;
      RECT MASK 2 36.314 102.96 36.374 104.01 ;
      RECT MASK 2 36.588 102.96 36.648 104.01 ;
      RECT MASK 2 36.862 102.96 36.922 104.01 ;
      RECT MASK 2 37.136 102.96 37.196 104.01 ;
      RECT MASK 2 37.41 102.96 37.47 104.01 ;
      RECT MASK 2 37.684 102.96 37.744 104.01 ;
      RECT MASK 2 37.958 102.96 38.018 104.01 ;
      RECT MASK 2 38.232 102.96 38.292 104.01 ;
      RECT MASK 2 38.506 102.96 38.566 104.01 ;
      RECT MASK 2 38.78 102.96 38.84 104.01 ;
      RECT MASK 2 39.054 102.96 39.114 104.01 ;
      RECT MASK 2 39.328 102.96 39.388 104.01 ;
      RECT MASK 2 39.602 102.96 39.662 104.01 ;
      RECT MASK 2 39.876 102.96 39.936 104.01 ;
      RECT MASK 2 40.15 102.96 40.21 104.01 ;
      RECT MASK 2 40.424 102.96 40.484 104.01 ;
      RECT MASK 2 40.698 102.96 40.758 104.01 ;
      RECT MASK 2 40.972 102.96 41.032 104.01 ;
      RECT MASK 2 41.246 102.96 41.306 104.01 ;
      RECT MASK 2 41.52 102.96 41.58 104.01 ;
      RECT MASK 2 41.794 102.96 41.854 104.01 ;
      RECT MASK 2 42.068 102.96 42.128 104.01 ;
      RECT MASK 2 42.342 102.96 42.402 104.01 ;
      RECT MASK 2 42.616 102.96 42.676 104.01 ;
      RECT MASK 2 42.89 102.96 42.95 104.01 ;
      RECT MASK 2 43.164 102.96 43.224 104.01 ;
      RECT MASK 2 43.438 102.96 43.498 104.01 ;
      RECT MASK 2 45.73 102.96 45.79 104.01 ;
      RECT MASK 2 46.004 102.96 46.064 104.01 ;
      RECT MASK 2 46.278 102.96 46.338 104.01 ;
      RECT MASK 2 46.552 102.96 46.612 104.01 ;
      RECT MASK 2 46.826 102.96 46.886 104.01 ;
      RECT MASK 2 47.1 102.96 47.16 104.01 ;
      RECT MASK 2 47.374 102.96 47.434 104.01 ;
      RECT MASK 2 47.648 102.96 47.708 104.01 ;
      RECT MASK 2 47.922 102.96 47.982 104.01 ;
      RECT MASK 2 48.196 102.96 48.256 104.01 ;
      RECT MASK 2 48.47 102.96 48.53 104.01 ;
      RECT MASK 2 48.744 102.96 48.804 104.01 ;
      RECT MASK 2 49.018 102.96 49.078 104.01 ;
      RECT MASK 2 49.292 102.96 49.352 104.01 ;
      RECT MASK 2 49.566 102.96 49.626 104.01 ;
      RECT MASK 2 49.84 102.96 49.9 104.01 ;
      RECT MASK 2 50.114 102.96 50.174 104.01 ;
      RECT MASK 2 50.388 102.96 50.448 104.01 ;
      RECT MASK 2 50.662 102.96 50.722 104.01 ;
      RECT MASK 2 50.936 102.96 50.996 104.01 ;
      RECT MASK 2 51.21 102.96 51.27 104.01 ;
      RECT MASK 2 51.484 102.96 51.544 104.01 ;
      RECT MASK 2 51.758 102.96 51.818 104.01 ;
      RECT MASK 2 52.032 102.96 52.092 104.01 ;
      RECT MASK 2 52.306 102.96 52.366 104.01 ;
      RECT MASK 2 52.58 102.96 52.64 104.01 ;
      RECT MASK 2 52.854 102.96 52.914 104.01 ;
      RECT MASK 2 53.128 102.96 53.188 104.01 ;
      RECT MASK 2 53.402 102.96 53.462 104.01 ;
      RECT MASK 2 53.676 102.96 53.736 104.01 ;
      RECT MASK 2 53.95 102.96 54.01 104.01 ;
      RECT MASK 2 54.224 102.96 54.284 104.01 ;
      RECT MASK 2 54.498 102.96 54.558 104.01 ;
      RECT MASK 2 54.772 102.96 54.832 104.01 ;
      RECT MASK 2 55.046 102.96 55.106 104.01 ;
      RECT MASK 2 55.32 102.96 55.38 104.01 ;
      RECT MASK 2 55.594 102.96 55.654 104.01 ;
      RECT MASK 2 55.868 102.96 55.928 104.01 ;
      RECT MASK 2 56.142 102.96 56.202 104.01 ;
      RECT MASK 2 56.416 102.96 56.476 104.01 ;
      RECT MASK 2 56.69 102.96 56.75 104.01 ;
      RECT MASK 2 56.964 102.96 57.024 104.01 ;
      RECT MASK 2 57.238 102.96 57.298 104.01 ;
      RECT MASK 2 57.512 102.96 57.572 104.01 ;
      RECT MASK 2 57.786 102.96 57.846 104.01 ;
      RECT MASK 2 58.06 102.96 58.12 104.01 ;
      RECT MASK 2 58.334 102.96 58.394 104.01 ;
      RECT MASK 2 58.608 102.96 58.668 104.01 ;
      RECT MASK 2 58.882 102.96 58.942 104.01 ;
      RECT MASK 2 59.156 102.96 59.216 104.01 ;
      RECT MASK 2 59.43 102.96 59.49 104.01 ;
      RECT MASK 2 59.704 102.96 59.764 104.01 ;
      RECT MASK 2 59.978 102.96 60.038 104.01 ;
      RECT MASK 2 60.252 102.96 60.312 104.01 ;
      RECT MASK 2 60.526 102.96 60.586 104.01 ;
      RECT MASK 2 60.8 102.96 60.86 104.01 ;
      RECT MASK 2 61.074 102.96 61.134 104.01 ;
      RECT MASK 2 61.348 102.96 61.408 104.01 ;
      RECT MASK 2 61.622 102.96 61.682 104.01 ;
      RECT MASK 2 61.896 102.96 61.956 104.01 ;
      RECT MASK 2 62.17 102.96 62.23 104.01 ;
      RECT MASK 2 62.444 102.96 62.504 104.01 ;
      RECT MASK 2 62.718 102.96 62.778 104.01 ;
      RECT MASK 2 62.992 102.96 63.052 104.01 ;
      RECT MASK 2 63.266 102.96 63.326 104.01 ;
      RECT MASK 2 63.54 102.96 63.6 104.01 ;
      RECT MASK 2 63.814 102.96 63.874 104.01 ;
      RECT MASK 2 64.088 102.96 64.148 104.01 ;
      RECT MASK 2 64.362 102.96 64.422 104.01 ;
      RECT MASK 2 64.636 102.96 64.696 104.01 ;
      RECT MASK 2 64.91 102.96 64.97 104.01 ;
      RECT MASK 2 65.184 102.96 65.244 104.01 ;
      RECT MASK 2 65.458 102.96 65.518 104.01 ;
      RECT MASK 2 65.732 102.96 65.792 104.01 ;
      RECT MASK 2 66.006 102.96 66.066 104.01 ;
      RECT MASK 2 66.28 102.96 66.34 104.01 ;
      RECT MASK 2 66.554 102.96 66.614 104.01 ;
      RECT MASK 2 66.828 102.96 66.888 104.01 ;
      RECT MASK 2 67.102 102.96 67.162 104.01 ;
      RECT MASK 2 67.376 102.96 67.436 104.01 ;
      RECT MASK 2 67.65 102.96 67.71 104.01 ;
      RECT MASK 2 67.924 102.96 67.984 104.01 ;
      RECT MASK 2 68.198 102.96 68.258 104.01 ;
      RECT MASK 2 68.472 102.96 68.532 104.01 ;
      RECT MASK 2 68.746 102.96 68.806 104.01 ;
      RECT MASK 2 69.02 102.96 69.08 104.01 ;
      RECT MASK 2 69.294 102.96 69.354 104.01 ;
      RECT MASK 2 69.568 102.96 69.628 104.01 ;
      RECT MASK 2 69.842 102.96 69.902 104.01 ;
      RECT MASK 2 70.116 102.96 70.176 104.01 ;
      RECT MASK 2 70.39 102.96 70.45 104.01 ;
      RECT MASK 2 70.664 102.96 70.724 104.01 ;
      RECT MASK 2 70.938 102.96 70.998 104.01 ;
      RECT MASK 2 71.212 102.96 71.272 104.01 ;
      RECT MASK 2 71.486 102.96 71.546 104.01 ;
      RECT MASK 2 71.76 102.96 71.82 104.01 ;
      RECT MASK 2 72.034 102.96 72.094 104.01 ;
      RECT MASK 2 72.308 102.96 72.368 104.01 ;
      RECT MASK 2 72.582 102.96 72.642 104.01 ;
      RECT MASK 2 72.856 102.96 72.916 104.01 ;
      RECT MASK 2 73.13 102.96 73.19 104.01 ;
      RECT MASK 2 73.404 102.96 73.464 104.01 ;
      RECT MASK 2 73.678 102.96 73.738 104.01 ;
      RECT MASK 2 73.952 102.96 74.012 104.01 ;
      RECT MASK 2 74.226 102.96 74.286 104.01 ;
      RECT MASK 2 74.5 102.96 74.56 104.01 ;
      RECT MASK 2 74.774 102.96 74.834 104.01 ;
      RECT MASK 2 75.048 102.96 75.108 104.01 ;
      RECT MASK 2 75.322 102.96 75.382 104.01 ;
      RECT MASK 2 75.596 102.96 75.656 104.01 ;
      RECT MASK 2 75.87 102.96 75.93 104.01 ;
      RECT MASK 2 76.144 102.96 76.204 104.01 ;
      RECT MASK 2 76.418 102.96 76.478 104.01 ;
      RECT MASK 2 76.692 102.96 76.752 104.01 ;
      RECT MASK 2 76.966 102.96 77.026 104.01 ;
      RECT MASK 2 77.24 102.96 77.3 104.01 ;
      RECT MASK 2 77.514 102.96 77.574 104.01 ;
      RECT MASK 2 77.788 102.96 77.848 104.01 ;
      RECT MASK 2 78.062 102.96 78.122 104.01 ;
      RECT MASK 2 78.336 102.96 78.396 104.01 ;
      RECT MASK 2 78.61 102.96 78.67 104.01 ;
      RECT MASK 2 78.884 102.96 78.944 104.01 ;
      RECT MASK 2 79.158 102.96 79.218 104.01 ;
      RECT MASK 2 79.432 102.96 79.492 104.01 ;
      RECT MASK 2 79.706 102.96 79.766 104.01 ;
      RECT MASK 2 79.98 102.96 80.04 104.01 ;
      RECT MASK 2 80.254 102.96 80.314 104.01 ;
      RECT MASK 2 80.528 102.96 80.588 104.01 ;
      RECT MASK 2 80.802 102.96 80.862 104.01 ;
      RECT MASK 2 81.076 102.96 81.136 104.01 ;
      RECT MASK 2 81.35 102.96 81.41 104.01 ;
      RECT MASK 2 81.624 102.96 81.684 104.01 ;
      RECT MASK 2 81.898 102.96 81.958 104.01 ;
      RECT MASK 2 82.172 102.96 82.232 104.01 ;
      RECT MASK 2 82.446 102.96 82.506 104.01 ;
      RECT MASK 2 82.72 102.96 82.78 104.01 ;
      RECT MASK 2 82.994 102.96 83.054 104.01 ;
      RECT MASK 2 83.268 102.96 83.328 104.01 ;
      RECT MASK 2 83.542 102.96 83.602 104.01 ;
      RECT MASK 2 83.816 102.96 83.876 104.01 ;
      RECT MASK 2 84.09 102.96 84.15 104.01 ;
      RECT MASK 2 84.364 102.96 84.424 104.01 ;
      RECT MASK 2 84.638 102.96 84.698 104.01 ;
      RECT MASK 2 84.912 102.96 84.972 104.01 ;
      RECT MASK 2 85.186 102.96 85.246 104.01 ;
      RECT MASK 2 85.46 102.96 85.52 104.01 ;
      RECT MASK 2 85.734 102.96 85.794 104.01 ;
      RECT MASK 2 86.008 102.96 86.068 104.01 ;
      RECT MASK 2 86.282 102.96 86.342 104.01 ;
      RECT MASK 2 86.556 102.96 86.616 104.01 ;
      RECT MASK 2 86.83 102.96 86.89 104.01 ;
      RECT MASK 2 89.089 102.96 89.149 104.01 ;
      RECT MASK 2 89.363 102.96 89.423 104.01 ;
      RECT MASK 2 89.637 102.96 89.697 104.01 ;
      RECT MASK 2 89.911 102.96 89.971 104.01 ;
      RECT MASK 2 90.185 102.96 90.245 104.01 ;
      RECT MASK 2 90.459 102.96 90.519 104.01 ;
      RECT MASK 2 90.733 102.96 90.793 104.01 ;
      RECT MASK 2 91.007 102.96 91.067 104.01 ;
      RECT MASK 2 91.281 102.96 91.341 104.01 ;
      RECT MASK 2 91.555 102.96 91.615 104.01 ;
      RECT MASK 2 91.829 102.96 91.889 104.01 ;
      RECT MASK 2 92.103 102.96 92.163 104.01 ;
      RECT MASK 2 92.377 102.96 92.437 104.01 ;
      RECT MASK 2 92.651 102.96 92.711 104.01 ;
      RECT MASK 2 92.925 102.96 92.985 104.01 ;
      RECT MASK 2 93.199 102.96 93.259 104.01 ;
      RECT MASK 2 93.473 102.96 93.533 104.01 ;
      RECT MASK 2 93.747 102.96 93.807 104.01 ;
      RECT MASK 2 94.021 102.96 94.081 104.01 ;
      RECT MASK 2 94.295 102.96 94.355 104.01 ;
      RECT MASK 2 94.569 102.96 94.629 104.01 ;
      RECT MASK 2 94.843 102.96 94.903 104.01 ;
      RECT MASK 2 95.117 102.96 95.177 104.01 ;
      RECT MASK 2 95.391 102.96 95.451 104.01 ;
      RECT MASK 2 95.665 102.96 95.725 104.01 ;
      RECT MASK 2 95.939 102.96 95.999 104.01 ;
      RECT MASK 2 96.213 102.96 96.273 104.01 ;
      RECT MASK 2 96.487 102.96 96.547 104.01 ;
      RECT MASK 2 96.761 102.96 96.821 104.01 ;
      RECT MASK 2 97.035 102.96 97.095 104.01 ;
      RECT MASK 2 97.309 102.96 97.369 104.01 ;
      RECT MASK 2 97.583 102.96 97.643 104.01 ;
      RECT MASK 2 97.857 102.96 97.917 104.01 ;
      RECT MASK 2 98.131 102.96 98.191 104.01 ;
      RECT MASK 2 98.405 102.96 98.465 104.01 ;
      RECT MASK 2 98.679 102.96 98.739 104.01 ;
      RECT MASK 2 98.953 102.96 99.013 104.01 ;
      RECT MASK 2 99.227 102.96 99.287 104.01 ;
      RECT MASK 2 99.501 102.96 99.561 104.01 ;
      RECT MASK 2 99.775 102.96 99.835 104.01 ;
      RECT MASK 2 100.049 102.96 100.109 104.01 ;
      RECT MASK 2 100.323 102.96 100.383 104.01 ;
      RECT MASK 2 100.597 102.96 100.657 104.01 ;
      RECT MASK 2 100.871 102.96 100.931 104.01 ;
      RECT MASK 2 101.145 102.96 101.205 104.01 ;
      RECT MASK 2 101.419 102.96 101.479 104.01 ;
      RECT MASK 2 101.693 102.96 101.753 104.01 ;
      RECT MASK 2 101.967 102.96 102.027 104.01 ;
      RECT MASK 2 102.241 102.96 102.301 104.01 ;
      RECT MASK 2 102.515 102.96 102.575 104.01 ;
      RECT MASK 2 102.789 102.96 102.849 104.01 ;
      RECT MASK 2 103.063 102.96 103.123 104.01 ;
      RECT MASK 2 103.337 102.96 103.397 104.01 ;
      RECT MASK 2 103.611 102.96 103.671 104.01 ;
      RECT MASK 2 103.885 102.96 103.945 104.01 ;
      RECT MASK 2 104.159 102.96 104.219 104.01 ;
      RECT MASK 2 104.433 102.96 104.493 104.01 ;
      RECT MASK 2 104.707 102.96 104.767 104.01 ;
      RECT MASK 2 104.981 102.96 105.041 104.01 ;
      RECT MASK 2 105.255 102.96 105.315 104.01 ;
      RECT MASK 2 105.529 102.96 105.589 104.01 ;
      RECT MASK 2 105.803 102.96 105.863 104.01 ;
      RECT MASK 2 106.077 102.96 106.137 104.01 ;
      RECT MASK 2 106.351 102.96 106.411 104.01 ;
      RECT MASK 2 106.625 102.96 106.685 104.01 ;
      RECT MASK 2 106.899 102.96 106.959 104.01 ;
      RECT MASK 2 107.173 102.96 107.233 104.01 ;
      RECT MASK 2 107.447 102.96 107.507 104.01 ;
      RECT MASK 2 107.721 102.96 107.781 104.01 ;
      RECT MASK 2 107.995 102.96 108.055 104.01 ;
      RECT MASK 2 108.269 102.96 108.329 104.01 ;
      RECT MASK 2 108.543 102.96 108.603 104.01 ;
      RECT MASK 2 108.817 102.96 108.877 104.01 ;
      RECT MASK 2 109.091 102.96 109.151 104.01 ;
      RECT MASK 2 109.365 102.96 109.425 104.01 ;
      RECT MASK 2 109.639 102.96 109.699 104.01 ;
      RECT MASK 2 109.913 102.96 109.973 104.01 ;
      RECT MASK 2 110.187 102.96 110.247 104.01 ;
      RECT MASK 2 110.461 102.96 110.521 104.01 ;
      RECT MASK 2 110.735 102.96 110.795 104.01 ;
      RECT MASK 2 111.009 102.96 111.069 104.01 ;
      RECT MASK 2 111.283 102.96 111.343 104.01 ;
      RECT MASK 2 111.557 102.96 111.617 104.01 ;
      RECT MASK 2 111.831 102.96 111.891 104.01 ;
      RECT MASK 2 112.105 102.96 112.165 104.01 ;
      RECT MASK 2 112.379 102.96 112.439 104.01 ;
      RECT MASK 2 112.653 102.96 112.713 104.01 ;
      RECT MASK 2 112.927 102.96 112.987 104.01 ;
      RECT MASK 2 113.201 102.96 113.261 104.01 ;
      RECT MASK 2 113.475 102.96 113.535 104.01 ;
      RECT MASK 2 113.749 102.96 113.809 104.01 ;
      RECT MASK 2 114.023 102.96 114.083 104.01 ;
      RECT MASK 2 114.297 102.96 114.357 104.01 ;
      RECT MASK 2 114.571 102.96 114.631 104.01 ;
      RECT MASK 2 114.845 102.96 114.905 104.01 ;
      RECT MASK 2 115.119 102.96 115.179 104.01 ;
      RECT MASK 2 115.393 102.96 115.453 104.01 ;
      RECT MASK 2 115.667 102.96 115.727 104.01 ;
      RECT MASK 2 115.941 102.96 116.001 104.01 ;
      RECT MASK 2 116.215 102.96 116.275 104.01 ;
      RECT MASK 2 116.489 102.96 116.549 104.01 ;
      RECT MASK 2 116.763 102.96 116.823 104.01 ;
      RECT MASK 2 117.037 102.96 117.097 104.01 ;
      RECT MASK 2 117.311 102.96 117.371 104.01 ;
      RECT MASK 2 117.585 102.96 117.645 104.01 ;
      RECT MASK 2 117.859 102.96 117.919 104.01 ;
      RECT MASK 2 118.133 102.96 118.193 104.01 ;
      RECT MASK 2 118.407 102.96 118.467 104.01 ;
      RECT MASK 2 118.681 102.96 118.741 104.01 ;
      RECT MASK 2 118.955 102.96 119.015 104.01 ;
      RECT MASK 2 119.229 102.96 119.289 104.01 ;
      RECT MASK 2 119.503 102.96 119.563 104.01 ;
      RECT MASK 2 119.777 102.96 119.837 104.01 ;
      RECT MASK 2 120.051 102.96 120.111 104.01 ;
      RECT MASK 2 120.325 102.96 120.385 104.01 ;
      RECT MASK 2 120.599 102.96 120.659 104.01 ;
      RECT MASK 2 120.873 102.96 120.933 104.01 ;
      RECT MASK 2 121.147 102.96 121.207 104.01 ;
      RECT MASK 2 121.421 102.96 121.481 104.01 ;
      RECT MASK 2 121.695 102.96 121.755 104.01 ;
      RECT MASK 2 121.969 102.96 122.029 104.01 ;
      RECT MASK 2 122.243 102.96 122.303 104.01 ;
      RECT MASK 2 122.517 102.96 122.577 104.01 ;
      RECT MASK 2 122.791 102.96 122.851 104.01 ;
      RECT MASK 2 123.065 102.96 123.125 104.01 ;
      RECT MASK 2 123.339 102.96 123.399 104.01 ;
      RECT MASK 2 123.613 102.96 123.673 104.01 ;
      RECT MASK 2 123.887 102.96 123.947 104.01 ;
      RECT MASK 2 124.161 102.96 124.221 104.01 ;
      RECT MASK 2 124.435 102.96 124.495 104.01 ;
      RECT MASK 2 124.709 102.96 124.769 104.01 ;
      RECT MASK 2 124.983 102.96 125.043 104.01 ;
      RECT MASK 2 125.257 102.96 125.317 104.01 ;
      RECT MASK 2 125.531 102.96 125.591 104.01 ;
      RECT MASK 2 125.805 102.96 125.865 104.01 ;
      RECT MASK 2 126.079 102.96 126.139 104.01 ;
      RECT MASK 2 126.353 102.96 126.413 104.01 ;
      RECT MASK 2 126.627 102.96 126.687 104.01 ;
      RECT MASK 2 126.901 102.96 126.961 104.01 ;
      RECT MASK 2 127.175 102.96 127.235 104.01 ;
      RECT MASK 2 127.449 102.96 127.509 104.01 ;
      RECT MASK 2 2.338 104.67 2.398 105.72 ;
      RECT MASK 2 2.612 104.67 2.672 105.72 ;
      RECT MASK 2 2.886 104.67 2.946 105.72 ;
      RECT MASK 2 3.16 104.67 3.22 105.72 ;
      RECT MASK 2 3.434 104.67 3.494 105.72 ;
      RECT MASK 2 3.708 104.67 3.768 105.72 ;
      RECT MASK 2 3.982 104.67 4.042 105.72 ;
      RECT MASK 2 4.256 104.67 4.316 105.72 ;
      RECT MASK 2 4.53 104.67 4.59 105.72 ;
      RECT MASK 2 4.804 104.67 4.864 105.72 ;
      RECT MASK 2 5.078 104.67 5.138 105.72 ;
      RECT MASK 2 5.352 104.67 5.412 105.72 ;
      RECT MASK 2 5.626 104.67 5.686 105.72 ;
      RECT MASK 2 5.9 104.67 5.96 105.72 ;
      RECT MASK 2 6.174 104.67 6.234 105.72 ;
      RECT MASK 2 6.448 104.67 6.508 105.72 ;
      RECT MASK 2 6.722 104.67 6.782 105.72 ;
      RECT MASK 2 6.996 104.67 7.056 105.72 ;
      RECT MASK 2 7.27 104.67 7.33 105.72 ;
      RECT MASK 2 7.544 104.67 7.604 105.72 ;
      RECT MASK 2 7.818 104.67 7.878 105.72 ;
      RECT MASK 2 8.092 104.67 8.152 105.72 ;
      RECT MASK 2 8.366 104.67 8.426 105.72 ;
      RECT MASK 2 8.64 104.67 8.7 105.72 ;
      RECT MASK 2 8.914 104.67 8.974 105.72 ;
      RECT MASK 2 9.188 104.67 9.248 105.72 ;
      RECT MASK 2 9.462 104.67 9.522 105.72 ;
      RECT MASK 2 9.736 104.67 9.796 105.72 ;
      RECT MASK 2 10.01 104.67 10.07 105.72 ;
      RECT MASK 2 10.284 104.67 10.344 105.72 ;
      RECT MASK 2 10.558 104.67 10.618 105.72 ;
      RECT MASK 2 10.832 104.67 10.892 105.72 ;
      RECT MASK 2 11.106 104.67 11.166 105.72 ;
      RECT MASK 2 11.38 104.67 11.44 105.72 ;
      RECT MASK 2 11.654 104.67 11.714 105.72 ;
      RECT MASK 2 11.928 104.67 11.988 105.72 ;
      RECT MASK 2 12.202 104.67 12.262 105.72 ;
      RECT MASK 2 12.476 104.67 12.536 105.72 ;
      RECT MASK 2 12.75 104.67 12.81 105.72 ;
      RECT MASK 2 13.024 104.67 13.084 105.72 ;
      RECT MASK 2 13.298 104.67 13.358 105.72 ;
      RECT MASK 2 13.572 104.67 13.632 105.72 ;
      RECT MASK 2 13.846 104.67 13.906 105.72 ;
      RECT MASK 2 14.12 104.67 14.18 105.72 ;
      RECT MASK 2 14.394 104.67 14.454 105.72 ;
      RECT MASK 2 14.668 104.67 14.728 105.72 ;
      RECT MASK 2 14.942 104.67 15.002 105.72 ;
      RECT MASK 2 15.216 104.67 15.276 105.72 ;
      RECT MASK 2 15.49 104.67 15.55 105.72 ;
      RECT MASK 2 15.764 104.67 15.824 105.72 ;
      RECT MASK 2 16.038 104.67 16.098 105.72 ;
      RECT MASK 2 16.312 104.67 16.372 105.72 ;
      RECT MASK 2 16.586 104.67 16.646 105.72 ;
      RECT MASK 2 16.86 104.67 16.92 105.72 ;
      RECT MASK 2 17.134 104.67 17.194 105.72 ;
      RECT MASK 2 17.408 104.67 17.468 105.72 ;
      RECT MASK 2 17.682 104.67 17.742 105.72 ;
      RECT MASK 2 17.956 104.67 18.016 105.72 ;
      RECT MASK 2 18.23 104.67 18.29 105.72 ;
      RECT MASK 2 18.504 104.67 18.564 105.72 ;
      RECT MASK 2 18.778 104.67 18.838 105.72 ;
      RECT MASK 2 19.052 104.67 19.112 105.72 ;
      RECT MASK 2 19.326 104.67 19.386 105.72 ;
      RECT MASK 2 19.6 104.67 19.66 105.72 ;
      RECT MASK 2 19.874 104.67 19.934 105.72 ;
      RECT MASK 2 20.148 104.67 20.208 105.72 ;
      RECT MASK 2 20.422 104.67 20.482 105.72 ;
      RECT MASK 2 20.696 104.67 20.756 105.72 ;
      RECT MASK 2 20.97 104.67 21.03 105.72 ;
      RECT MASK 2 21.244 104.67 21.304 105.72 ;
      RECT MASK 2 21.518 104.67 21.578 105.72 ;
      RECT MASK 2 21.792 104.67 21.852 105.72 ;
      RECT MASK 2 22.066 104.67 22.126 105.72 ;
      RECT MASK 2 22.34 104.67 22.4 105.72 ;
      RECT MASK 2 22.614 104.67 22.674 105.72 ;
      RECT MASK 2 22.888 104.67 22.948 105.72 ;
      RECT MASK 2 23.162 104.67 23.222 105.72 ;
      RECT MASK 2 23.436 104.67 23.496 105.72 ;
      RECT MASK 2 23.71 104.67 23.77 105.72 ;
      RECT MASK 2 23.984 104.67 24.044 105.72 ;
      RECT MASK 2 24.258 104.67 24.318 105.72 ;
      RECT MASK 2 24.532 104.67 24.592 105.72 ;
      RECT MASK 2 24.806 104.67 24.866 105.72 ;
      RECT MASK 2 25.08 104.67 25.14 105.72 ;
      RECT MASK 2 25.354 104.67 25.414 105.72 ;
      RECT MASK 2 25.628 104.67 25.688 105.72 ;
      RECT MASK 2 25.902 104.67 25.962 105.72 ;
      RECT MASK 2 26.176 104.67 26.236 105.72 ;
      RECT MASK 2 26.45 104.67 26.51 105.72 ;
      RECT MASK 2 26.724 104.67 26.784 105.72 ;
      RECT MASK 2 26.998 104.67 27.058 105.72 ;
      RECT MASK 2 27.272 104.67 27.332 105.72 ;
      RECT MASK 2 27.546 104.67 27.606 105.72 ;
      RECT MASK 2 27.82 104.67 27.88 105.72 ;
      RECT MASK 2 28.094 104.67 28.154 105.72 ;
      RECT MASK 2 28.368 104.67 28.428 105.72 ;
      RECT MASK 2 28.642 104.67 28.702 105.72 ;
      RECT MASK 2 28.916 104.67 28.976 105.72 ;
      RECT MASK 2 29.19 104.67 29.25 105.72 ;
      RECT MASK 2 29.464 104.67 29.524 105.72 ;
      RECT MASK 2 29.738 104.67 29.798 105.72 ;
      RECT MASK 2 30.012 104.67 30.072 105.72 ;
      RECT MASK 2 30.286 104.67 30.346 105.72 ;
      RECT MASK 2 30.56 104.67 30.62 105.72 ;
      RECT MASK 2 30.834 104.67 30.894 105.72 ;
      RECT MASK 2 31.108 104.67 31.168 105.72 ;
      RECT MASK 2 31.382 104.67 31.442 105.72 ;
      RECT MASK 2 31.656 104.67 31.716 105.72 ;
      RECT MASK 2 31.93 104.67 31.99 105.72 ;
      RECT MASK 2 32.204 104.67 32.264 105.72 ;
      RECT MASK 2 32.478 104.67 32.538 105.72 ;
      RECT MASK 2 32.752 104.67 32.812 105.72 ;
      RECT MASK 2 33.026 104.67 33.086 105.72 ;
      RECT MASK 2 33.3 104.67 33.36 105.72 ;
      RECT MASK 2 33.574 104.67 33.634 105.72 ;
      RECT MASK 2 33.848 104.67 33.908 105.72 ;
      RECT MASK 2 34.122 104.67 34.182 105.72 ;
      RECT MASK 2 34.396 104.67 34.456 105.72 ;
      RECT MASK 2 34.67 104.67 34.73 105.72 ;
      RECT MASK 2 34.944 104.67 35.004 105.72 ;
      RECT MASK 2 35.218 104.67 35.278 105.72 ;
      RECT MASK 2 35.492 104.67 35.552 105.72 ;
      RECT MASK 2 35.766 104.67 35.826 105.72 ;
      RECT MASK 2 36.04 104.67 36.1 105.72 ;
      RECT MASK 2 36.314 104.67 36.374 105.72 ;
      RECT MASK 2 36.588 104.67 36.648 105.72 ;
      RECT MASK 2 36.862 104.67 36.922 105.72 ;
      RECT MASK 2 37.136 104.67 37.196 105.72 ;
      RECT MASK 2 37.41 104.67 37.47 105.72 ;
      RECT MASK 2 37.684 104.67 37.744 105.72 ;
      RECT MASK 2 37.958 104.67 38.018 105.72 ;
      RECT MASK 2 38.232 104.67 38.292 105.72 ;
      RECT MASK 2 38.506 104.67 38.566 105.72 ;
      RECT MASK 2 38.78 104.67 38.84 105.72 ;
      RECT MASK 2 39.054 104.67 39.114 105.72 ;
      RECT MASK 2 39.328 104.67 39.388 105.72 ;
      RECT MASK 2 39.602 104.67 39.662 105.72 ;
      RECT MASK 2 39.876 104.67 39.936 105.72 ;
      RECT MASK 2 40.15 104.67 40.21 105.72 ;
      RECT MASK 2 40.424 104.67 40.484 105.72 ;
      RECT MASK 2 40.698 104.67 40.758 105.72 ;
      RECT MASK 2 40.972 104.67 41.032 105.72 ;
      RECT MASK 2 41.246 104.67 41.306 105.72 ;
      RECT MASK 2 41.52 104.67 41.58 105.72 ;
      RECT MASK 2 41.794 104.67 41.854 105.72 ;
      RECT MASK 2 42.068 104.67 42.128 105.72 ;
      RECT MASK 2 42.342 104.67 42.402 105.72 ;
      RECT MASK 2 42.616 104.67 42.676 105.72 ;
      RECT MASK 2 42.89 104.67 42.95 105.72 ;
      RECT MASK 2 43.164 104.67 43.224 105.72 ;
      RECT MASK 2 43.438 104.67 43.498 105.72 ;
      RECT MASK 2 45.73 104.67 45.79 105.72 ;
      RECT MASK 2 46.004 104.67 46.064 105.72 ;
      RECT MASK 2 46.278 104.67 46.338 105.72 ;
      RECT MASK 2 46.552 104.67 46.612 105.72 ;
      RECT MASK 2 46.826 104.67 46.886 105.72 ;
      RECT MASK 2 47.1 104.67 47.16 105.72 ;
      RECT MASK 2 47.374 104.67 47.434 105.72 ;
      RECT MASK 2 47.648 104.67 47.708 105.72 ;
      RECT MASK 2 47.922 104.67 47.982 105.72 ;
      RECT MASK 2 48.196 104.67 48.256 105.72 ;
      RECT MASK 2 48.47 104.67 48.53 105.72 ;
      RECT MASK 2 48.744 104.67 48.804 105.72 ;
      RECT MASK 2 49.018 104.67 49.078 105.72 ;
      RECT MASK 2 49.292 104.67 49.352 105.72 ;
      RECT MASK 2 49.566 104.67 49.626 105.72 ;
      RECT MASK 2 49.84 104.67 49.9 105.72 ;
      RECT MASK 2 50.114 104.67 50.174 105.72 ;
      RECT MASK 2 50.388 104.67 50.448 105.72 ;
      RECT MASK 2 50.662 104.67 50.722 105.72 ;
      RECT MASK 2 50.936 104.67 50.996 105.72 ;
      RECT MASK 2 51.21 104.67 51.27 105.72 ;
      RECT MASK 2 51.484 104.67 51.544 105.72 ;
      RECT MASK 2 51.758 104.67 51.818 105.72 ;
      RECT MASK 2 52.032 104.67 52.092 105.72 ;
      RECT MASK 2 52.306 104.67 52.366 105.72 ;
      RECT MASK 2 52.58 104.67 52.64 105.72 ;
      RECT MASK 2 52.854 104.67 52.914 105.72 ;
      RECT MASK 2 53.128 104.67 53.188 105.72 ;
      RECT MASK 2 53.402 104.67 53.462 105.72 ;
      RECT MASK 2 53.676 104.67 53.736 105.72 ;
      RECT MASK 2 53.95 104.67 54.01 105.72 ;
      RECT MASK 2 54.224 104.67 54.284 105.72 ;
      RECT MASK 2 54.498 104.67 54.558 105.72 ;
      RECT MASK 2 54.772 104.67 54.832 105.72 ;
      RECT MASK 2 55.046 104.67 55.106 105.72 ;
      RECT MASK 2 55.32 104.67 55.38 105.72 ;
      RECT MASK 2 55.594 104.67 55.654 105.72 ;
      RECT MASK 2 55.868 104.67 55.928 105.72 ;
      RECT MASK 2 56.142 104.67 56.202 105.72 ;
      RECT MASK 2 56.416 104.67 56.476 105.72 ;
      RECT MASK 2 56.69 104.67 56.75 105.72 ;
      RECT MASK 2 56.964 104.67 57.024 105.72 ;
      RECT MASK 2 57.238 104.67 57.298 105.72 ;
      RECT MASK 2 57.512 104.67 57.572 105.72 ;
      RECT MASK 2 57.786 104.67 57.846 105.72 ;
      RECT MASK 2 58.06 104.67 58.12 105.72 ;
      RECT MASK 2 58.334 104.67 58.394 105.72 ;
      RECT MASK 2 58.608 104.67 58.668 105.72 ;
      RECT MASK 2 58.882 104.67 58.942 105.72 ;
      RECT MASK 2 59.156 104.67 59.216 105.72 ;
      RECT MASK 2 59.43 104.67 59.49 105.72 ;
      RECT MASK 2 59.704 104.67 59.764 105.72 ;
      RECT MASK 2 59.978 104.67 60.038 105.72 ;
      RECT MASK 2 60.252 104.67 60.312 105.72 ;
      RECT MASK 2 60.526 104.67 60.586 105.72 ;
      RECT MASK 2 60.8 104.67 60.86 105.72 ;
      RECT MASK 2 61.074 104.67 61.134 105.72 ;
      RECT MASK 2 61.348 104.67 61.408 105.72 ;
      RECT MASK 2 61.622 104.67 61.682 105.72 ;
      RECT MASK 2 61.896 104.67 61.956 105.72 ;
      RECT MASK 2 62.17 104.67 62.23 105.72 ;
      RECT MASK 2 62.444 104.67 62.504 105.72 ;
      RECT MASK 2 62.718 104.67 62.778 105.72 ;
      RECT MASK 2 62.992 104.67 63.052 105.72 ;
      RECT MASK 2 63.266 104.67 63.326 105.72 ;
      RECT MASK 2 63.54 104.67 63.6 105.72 ;
      RECT MASK 2 63.814 104.67 63.874 105.72 ;
      RECT MASK 2 64.088 104.67 64.148 105.72 ;
      RECT MASK 2 64.362 104.67 64.422 105.72 ;
      RECT MASK 2 64.636 104.67 64.696 105.72 ;
      RECT MASK 2 64.91 104.67 64.97 105.72 ;
      RECT MASK 2 65.184 104.67 65.244 105.72 ;
      RECT MASK 2 65.458 104.67 65.518 105.72 ;
      RECT MASK 2 65.732 104.67 65.792 105.72 ;
      RECT MASK 2 66.006 104.67 66.066 105.72 ;
      RECT MASK 2 66.28 104.67 66.34 105.72 ;
      RECT MASK 2 66.554 104.67 66.614 105.72 ;
      RECT MASK 2 66.828 104.67 66.888 105.72 ;
      RECT MASK 2 67.102 104.67 67.162 105.72 ;
      RECT MASK 2 67.376 104.67 67.436 105.72 ;
      RECT MASK 2 67.65 104.67 67.71 105.72 ;
      RECT MASK 2 67.924 104.67 67.984 105.72 ;
      RECT MASK 2 68.198 104.67 68.258 105.72 ;
      RECT MASK 2 68.472 104.67 68.532 105.72 ;
      RECT MASK 2 68.746 104.67 68.806 105.72 ;
      RECT MASK 2 69.02 104.67 69.08 105.72 ;
      RECT MASK 2 69.294 104.67 69.354 105.72 ;
      RECT MASK 2 69.568 104.67 69.628 105.72 ;
      RECT MASK 2 69.842 104.67 69.902 105.72 ;
      RECT MASK 2 70.116 104.67 70.176 105.72 ;
      RECT MASK 2 70.39 104.67 70.45 105.72 ;
      RECT MASK 2 70.664 104.67 70.724 105.72 ;
      RECT MASK 2 70.938 104.67 70.998 105.72 ;
      RECT MASK 2 71.212 104.67 71.272 105.72 ;
      RECT MASK 2 71.486 104.67 71.546 105.72 ;
      RECT MASK 2 71.76 104.67 71.82 105.72 ;
      RECT MASK 2 72.034 104.67 72.094 105.72 ;
      RECT MASK 2 72.308 104.67 72.368 105.72 ;
      RECT MASK 2 72.582 104.67 72.642 105.72 ;
      RECT MASK 2 72.856 104.67 72.916 105.72 ;
      RECT MASK 2 73.13 104.67 73.19 105.72 ;
      RECT MASK 2 73.404 104.67 73.464 105.72 ;
      RECT MASK 2 73.678 104.67 73.738 105.72 ;
      RECT MASK 2 73.952 104.67 74.012 105.72 ;
      RECT MASK 2 74.226 104.67 74.286 105.72 ;
      RECT MASK 2 74.5 104.67 74.56 105.72 ;
      RECT MASK 2 74.774 104.67 74.834 105.72 ;
      RECT MASK 2 75.048 104.67 75.108 105.72 ;
      RECT MASK 2 75.322 104.67 75.382 105.72 ;
      RECT MASK 2 75.596 104.67 75.656 105.72 ;
      RECT MASK 2 75.87 104.67 75.93 105.72 ;
      RECT MASK 2 76.144 104.67 76.204 105.72 ;
      RECT MASK 2 76.418 104.67 76.478 105.72 ;
      RECT MASK 2 76.692 104.67 76.752 105.72 ;
      RECT MASK 2 76.966 104.67 77.026 105.72 ;
      RECT MASK 2 77.24 104.67 77.3 105.72 ;
      RECT MASK 2 77.514 104.67 77.574 105.72 ;
      RECT MASK 2 77.788 104.67 77.848 105.72 ;
      RECT MASK 2 78.062 104.67 78.122 105.72 ;
      RECT MASK 2 78.336 104.67 78.396 105.72 ;
      RECT MASK 2 78.61 104.67 78.67 105.72 ;
      RECT MASK 2 78.884 104.67 78.944 105.72 ;
      RECT MASK 2 79.158 104.67 79.218 105.72 ;
      RECT MASK 2 79.432 104.67 79.492 105.72 ;
      RECT MASK 2 79.706 104.67 79.766 105.72 ;
      RECT MASK 2 79.98 104.67 80.04 105.72 ;
      RECT MASK 2 80.254 104.67 80.314 105.72 ;
      RECT MASK 2 80.528 104.67 80.588 105.72 ;
      RECT MASK 2 80.802 104.67 80.862 105.72 ;
      RECT MASK 2 81.076 104.67 81.136 105.72 ;
      RECT MASK 2 81.35 104.67 81.41 105.72 ;
      RECT MASK 2 81.624 104.67 81.684 105.72 ;
      RECT MASK 2 81.898 104.67 81.958 105.72 ;
      RECT MASK 2 82.172 104.67 82.232 105.72 ;
      RECT MASK 2 82.446 104.67 82.506 105.72 ;
      RECT MASK 2 82.72 104.67 82.78 105.72 ;
      RECT MASK 2 82.994 104.67 83.054 105.72 ;
      RECT MASK 2 83.268 104.67 83.328 105.72 ;
      RECT MASK 2 83.542 104.67 83.602 105.72 ;
      RECT MASK 2 83.816 104.67 83.876 105.72 ;
      RECT MASK 2 84.09 104.67 84.15 105.72 ;
      RECT MASK 2 84.364 104.67 84.424 105.72 ;
      RECT MASK 2 84.638 104.67 84.698 105.72 ;
      RECT MASK 2 84.912 104.67 84.972 105.72 ;
      RECT MASK 2 85.186 104.67 85.246 105.72 ;
      RECT MASK 2 85.46 104.67 85.52 105.72 ;
      RECT MASK 2 85.734 104.67 85.794 105.72 ;
      RECT MASK 2 86.008 104.67 86.068 105.72 ;
      RECT MASK 2 86.282 104.67 86.342 105.72 ;
      RECT MASK 2 86.556 104.67 86.616 105.72 ;
      RECT MASK 2 86.83 104.67 86.89 105.72 ;
      RECT MASK 2 89.089 104.67 89.149 105.72 ;
      RECT MASK 2 89.363 104.67 89.423 105.72 ;
      RECT MASK 2 89.637 104.67 89.697 105.72 ;
      RECT MASK 2 89.911 104.67 89.971 105.72 ;
      RECT MASK 2 90.185 104.67 90.245 105.72 ;
      RECT MASK 2 90.459 104.67 90.519 105.72 ;
      RECT MASK 2 90.733 104.67 90.793 105.72 ;
      RECT MASK 2 91.007 104.67 91.067 105.72 ;
      RECT MASK 2 91.281 104.67 91.341 105.72 ;
      RECT MASK 2 91.555 104.67 91.615 105.72 ;
      RECT MASK 2 91.829 104.67 91.889 105.72 ;
      RECT MASK 2 92.103 104.67 92.163 105.72 ;
      RECT MASK 2 92.377 104.67 92.437 105.72 ;
      RECT MASK 2 92.651 104.67 92.711 105.72 ;
      RECT MASK 2 92.925 104.67 92.985 105.72 ;
      RECT MASK 2 93.199 104.67 93.259 105.72 ;
      RECT MASK 2 93.473 104.67 93.533 105.72 ;
      RECT MASK 2 93.747 104.67 93.807 105.72 ;
      RECT MASK 2 94.021 104.67 94.081 105.72 ;
      RECT MASK 2 94.295 104.67 94.355 105.72 ;
      RECT MASK 2 94.569 104.67 94.629 105.72 ;
      RECT MASK 2 94.843 104.67 94.903 105.72 ;
      RECT MASK 2 95.117 104.67 95.177 105.72 ;
      RECT MASK 2 95.391 104.67 95.451 105.72 ;
      RECT MASK 2 95.665 104.67 95.725 105.72 ;
      RECT MASK 2 95.939 104.67 95.999 105.72 ;
      RECT MASK 2 96.213 104.67 96.273 105.72 ;
      RECT MASK 2 96.487 104.67 96.547 105.72 ;
      RECT MASK 2 96.761 104.67 96.821 105.72 ;
      RECT MASK 2 97.035 104.67 97.095 105.72 ;
      RECT MASK 2 97.309 104.67 97.369 105.72 ;
      RECT MASK 2 97.583 104.67 97.643 105.72 ;
      RECT MASK 2 97.857 104.67 97.917 105.72 ;
      RECT MASK 2 98.131 104.67 98.191 105.72 ;
      RECT MASK 2 98.405 104.67 98.465 105.72 ;
      RECT MASK 2 98.679 104.67 98.739 105.72 ;
      RECT MASK 2 98.953 104.67 99.013 105.72 ;
      RECT MASK 2 99.227 104.67 99.287 105.72 ;
      RECT MASK 2 99.501 104.67 99.561 105.72 ;
      RECT MASK 2 99.775 104.67 99.835 105.72 ;
      RECT MASK 2 100.049 104.67 100.109 105.72 ;
      RECT MASK 2 100.323 104.67 100.383 105.72 ;
      RECT MASK 2 100.597 104.67 100.657 105.72 ;
      RECT MASK 2 100.871 104.67 100.931 105.72 ;
      RECT MASK 2 101.145 104.67 101.205 105.72 ;
      RECT MASK 2 101.419 104.67 101.479 105.72 ;
      RECT MASK 2 101.693 104.67 101.753 105.72 ;
      RECT MASK 2 101.967 104.67 102.027 105.72 ;
      RECT MASK 2 102.241 104.67 102.301 105.72 ;
      RECT MASK 2 102.515 104.67 102.575 105.72 ;
      RECT MASK 2 102.789 104.67 102.849 105.72 ;
      RECT MASK 2 103.063 104.67 103.123 105.72 ;
      RECT MASK 2 103.337 104.67 103.397 105.72 ;
      RECT MASK 2 103.611 104.67 103.671 105.72 ;
      RECT MASK 2 103.885 104.67 103.945 105.72 ;
      RECT MASK 2 104.159 104.67 104.219 105.72 ;
      RECT MASK 2 104.433 104.67 104.493 105.72 ;
      RECT MASK 2 104.707 104.67 104.767 105.72 ;
      RECT MASK 2 104.981 104.67 105.041 105.72 ;
      RECT MASK 2 105.255 104.67 105.315 105.72 ;
      RECT MASK 2 105.529 104.67 105.589 105.72 ;
      RECT MASK 2 105.803 104.67 105.863 105.72 ;
      RECT MASK 2 106.077 104.67 106.137 105.72 ;
      RECT MASK 2 106.351 104.67 106.411 105.72 ;
      RECT MASK 2 106.625 104.67 106.685 105.72 ;
      RECT MASK 2 106.899 104.67 106.959 105.72 ;
      RECT MASK 2 107.173 104.67 107.233 105.72 ;
      RECT MASK 2 107.447 104.67 107.507 105.72 ;
      RECT MASK 2 107.721 104.67 107.781 105.72 ;
      RECT MASK 2 107.995 104.67 108.055 105.72 ;
      RECT MASK 2 108.269 104.67 108.329 105.72 ;
      RECT MASK 2 108.543 104.67 108.603 105.72 ;
      RECT MASK 2 108.817 104.67 108.877 105.72 ;
      RECT MASK 2 109.091 104.67 109.151 105.72 ;
      RECT MASK 2 109.365 104.67 109.425 105.72 ;
      RECT MASK 2 109.639 104.67 109.699 105.72 ;
      RECT MASK 2 109.913 104.67 109.973 105.72 ;
      RECT MASK 2 110.187 104.67 110.247 105.72 ;
      RECT MASK 2 110.461 104.67 110.521 105.72 ;
      RECT MASK 2 110.735 104.67 110.795 105.72 ;
      RECT MASK 2 111.009 104.67 111.069 105.72 ;
      RECT MASK 2 111.283 104.67 111.343 105.72 ;
      RECT MASK 2 111.557 104.67 111.617 105.72 ;
      RECT MASK 2 111.831 104.67 111.891 105.72 ;
      RECT MASK 2 112.105 104.67 112.165 105.72 ;
      RECT MASK 2 112.379 104.67 112.439 105.72 ;
      RECT MASK 2 112.653 104.67 112.713 105.72 ;
      RECT MASK 2 112.927 104.67 112.987 105.72 ;
      RECT MASK 2 113.201 104.67 113.261 105.72 ;
      RECT MASK 2 113.475 104.67 113.535 105.72 ;
      RECT MASK 2 113.749 104.67 113.809 105.72 ;
      RECT MASK 2 114.023 104.67 114.083 105.72 ;
      RECT MASK 2 114.297 104.67 114.357 105.72 ;
      RECT MASK 2 114.571 104.67 114.631 105.72 ;
      RECT MASK 2 114.845 104.67 114.905 105.72 ;
      RECT MASK 2 115.119 104.67 115.179 105.72 ;
      RECT MASK 2 115.393 104.67 115.453 105.72 ;
      RECT MASK 2 115.667 104.67 115.727 105.72 ;
      RECT MASK 2 115.941 104.67 116.001 105.72 ;
      RECT MASK 2 116.215 104.67 116.275 105.72 ;
      RECT MASK 2 116.489 104.67 116.549 105.72 ;
      RECT MASK 2 116.763 104.67 116.823 105.72 ;
      RECT MASK 2 117.037 104.67 117.097 105.72 ;
      RECT MASK 2 117.311 104.67 117.371 105.72 ;
      RECT MASK 2 117.585 104.67 117.645 105.72 ;
      RECT MASK 2 117.859 104.67 117.919 105.72 ;
      RECT MASK 2 118.133 104.67 118.193 105.72 ;
      RECT MASK 2 118.407 104.67 118.467 105.72 ;
      RECT MASK 2 118.681 104.67 118.741 105.72 ;
      RECT MASK 2 118.955 104.67 119.015 105.72 ;
      RECT MASK 2 119.229 104.67 119.289 105.72 ;
      RECT MASK 2 119.503 104.67 119.563 105.72 ;
      RECT MASK 2 119.777 104.67 119.837 105.72 ;
      RECT MASK 2 120.051 104.67 120.111 105.72 ;
      RECT MASK 2 120.325 104.67 120.385 105.72 ;
      RECT MASK 2 120.599 104.67 120.659 105.72 ;
      RECT MASK 2 120.873 104.67 120.933 105.72 ;
      RECT MASK 2 121.147 104.67 121.207 105.72 ;
      RECT MASK 2 121.421 104.67 121.481 105.72 ;
      RECT MASK 2 121.695 104.67 121.755 105.72 ;
      RECT MASK 2 121.969 104.67 122.029 105.72 ;
      RECT MASK 2 122.243 104.67 122.303 105.72 ;
      RECT MASK 2 122.517 104.67 122.577 105.72 ;
      RECT MASK 2 122.791 104.67 122.851 105.72 ;
      RECT MASK 2 123.065 104.67 123.125 105.72 ;
      RECT MASK 2 123.339 104.67 123.399 105.72 ;
      RECT MASK 2 123.613 104.67 123.673 105.72 ;
      RECT MASK 2 123.887 104.67 123.947 105.72 ;
      RECT MASK 2 124.161 104.67 124.221 105.72 ;
      RECT MASK 2 124.435 104.67 124.495 105.72 ;
      RECT MASK 2 124.709 104.67 124.769 105.72 ;
      RECT MASK 2 124.983 104.67 125.043 105.72 ;
      RECT MASK 2 125.257 104.67 125.317 105.72 ;
      RECT MASK 2 125.531 104.67 125.591 105.72 ;
      RECT MASK 2 125.805 104.67 125.865 105.72 ;
      RECT MASK 2 126.079 104.67 126.139 105.72 ;
      RECT MASK 2 126.353 104.67 126.413 105.72 ;
      RECT MASK 2 126.627 104.67 126.687 105.72 ;
      RECT MASK 2 126.901 104.67 126.961 105.72 ;
      RECT MASK 2 127.175 104.67 127.235 105.72 ;
      RECT MASK 2 127.449 104.67 127.509 105.72 ;
      RECT MASK 2 2.338 106.38 2.398 107.43 ;
      RECT MASK 2 2.612 106.38 2.672 107.43 ;
      RECT MASK 2 2.886 106.38 2.946 107.43 ;
      RECT MASK 2 3.16 106.38 3.22 107.43 ;
      RECT MASK 2 3.434 106.38 3.494 107.43 ;
      RECT MASK 2 3.708 106.38 3.768 107.43 ;
      RECT MASK 2 3.982 106.38 4.042 107.43 ;
      RECT MASK 2 4.256 106.38 4.316 107.43 ;
      RECT MASK 2 4.53 106.38 4.59 107.43 ;
      RECT MASK 2 4.804 106.38 4.864 107.43 ;
      RECT MASK 2 5.078 106.38 5.138 107.43 ;
      RECT MASK 2 5.352 106.38 5.412 107.43 ;
      RECT MASK 2 5.626 106.38 5.686 107.43 ;
      RECT MASK 2 5.9 106.38 5.96 107.43 ;
      RECT MASK 2 6.174 106.38 6.234 107.43 ;
      RECT MASK 2 6.448 106.38 6.508 107.43 ;
      RECT MASK 2 6.722 106.38 6.782 107.43 ;
      RECT MASK 2 6.996 106.38 7.056 107.43 ;
      RECT MASK 2 7.27 106.38 7.33 107.43 ;
      RECT MASK 2 7.544 106.38 7.604 107.43 ;
      RECT MASK 2 7.818 106.38 7.878 107.43 ;
      RECT MASK 2 8.092 106.38 8.152 107.43 ;
      RECT MASK 2 8.366 106.38 8.426 107.43 ;
      RECT MASK 2 8.64 106.38 8.7 107.43 ;
      RECT MASK 2 8.914 106.38 8.974 107.43 ;
      RECT MASK 2 9.188 106.38 9.248 107.43 ;
      RECT MASK 2 9.462 106.38 9.522 107.43 ;
      RECT MASK 2 9.736 106.38 9.796 107.43 ;
      RECT MASK 2 10.01 106.38 10.07 107.43 ;
      RECT MASK 2 10.284 106.38 10.344 107.43 ;
      RECT MASK 2 10.558 106.38 10.618 107.43 ;
      RECT MASK 2 10.832 106.38 10.892 107.43 ;
      RECT MASK 2 11.106 106.38 11.166 107.43 ;
      RECT MASK 2 11.38 106.38 11.44 107.43 ;
      RECT MASK 2 11.654 106.38 11.714 107.43 ;
      RECT MASK 2 11.928 106.38 11.988 107.43 ;
      RECT MASK 2 12.202 106.38 12.262 107.43 ;
      RECT MASK 2 12.476 106.38 12.536 107.43 ;
      RECT MASK 2 12.75 106.38 12.81 107.43 ;
      RECT MASK 2 13.024 106.38 13.084 107.43 ;
      RECT MASK 2 13.298 106.38 13.358 107.43 ;
      RECT MASK 2 13.572 106.38 13.632 107.43 ;
      RECT MASK 2 13.846 106.38 13.906 107.43 ;
      RECT MASK 2 14.12 106.38 14.18 107.43 ;
      RECT MASK 2 14.394 106.38 14.454 107.43 ;
      RECT MASK 2 14.668 106.38 14.728 107.43 ;
      RECT MASK 2 14.942 106.38 15.002 107.43 ;
      RECT MASK 2 15.216 106.38 15.276 107.43 ;
      RECT MASK 2 15.49 106.38 15.55 107.43 ;
      RECT MASK 2 15.764 106.38 15.824 107.43 ;
      RECT MASK 2 16.038 106.38 16.098 107.43 ;
      RECT MASK 2 16.312 106.38 16.372 107.43 ;
      RECT MASK 2 16.586 106.38 16.646 107.43 ;
      RECT MASK 2 16.86 106.38 16.92 107.43 ;
      RECT MASK 2 17.134 106.38 17.194 107.43 ;
      RECT MASK 2 17.408 106.38 17.468 107.43 ;
      RECT MASK 2 17.682 106.38 17.742 107.43 ;
      RECT MASK 2 17.956 106.38 18.016 107.43 ;
      RECT MASK 2 18.23 106.38 18.29 107.43 ;
      RECT MASK 2 18.504 106.38 18.564 107.43 ;
      RECT MASK 2 18.778 106.38 18.838 107.43 ;
      RECT MASK 2 19.052 106.38 19.112 107.43 ;
      RECT MASK 2 19.326 106.38 19.386 107.43 ;
      RECT MASK 2 19.6 106.38 19.66 107.43 ;
      RECT MASK 2 19.874 106.38 19.934 107.43 ;
      RECT MASK 2 20.148 106.38 20.208 107.43 ;
      RECT MASK 2 20.422 106.38 20.482 107.43 ;
      RECT MASK 2 20.696 106.38 20.756 107.43 ;
      RECT MASK 2 20.97 106.38 21.03 107.43 ;
      RECT MASK 2 21.244 106.38 21.304 107.43 ;
      RECT MASK 2 21.518 106.38 21.578 107.43 ;
      RECT MASK 2 21.792 106.38 21.852 107.43 ;
      RECT MASK 2 22.066 106.38 22.126 107.43 ;
      RECT MASK 2 22.34 106.38 22.4 107.43 ;
      RECT MASK 2 22.614 106.38 22.674 107.43 ;
      RECT MASK 2 22.888 106.38 22.948 107.43 ;
      RECT MASK 2 23.162 106.38 23.222 107.43 ;
      RECT MASK 2 23.436 106.38 23.496 107.43 ;
      RECT MASK 2 23.71 106.38 23.77 107.43 ;
      RECT MASK 2 23.984 106.38 24.044 107.43 ;
      RECT MASK 2 24.258 106.38 24.318 107.43 ;
      RECT MASK 2 24.532 106.38 24.592 107.43 ;
      RECT MASK 2 24.806 106.38 24.866 107.43 ;
      RECT MASK 2 25.08 106.38 25.14 107.43 ;
      RECT MASK 2 25.354 106.38 25.414 107.43 ;
      RECT MASK 2 25.628 106.38 25.688 107.43 ;
      RECT MASK 2 25.902 106.38 25.962 107.43 ;
      RECT MASK 2 26.176 106.38 26.236 107.43 ;
      RECT MASK 2 26.45 106.38 26.51 107.43 ;
      RECT MASK 2 26.724 106.38 26.784 107.43 ;
      RECT MASK 2 26.998 106.38 27.058 107.43 ;
      RECT MASK 2 27.272 106.38 27.332 107.43 ;
      RECT MASK 2 27.546 106.38 27.606 107.43 ;
      RECT MASK 2 27.82 106.38 27.88 107.43 ;
      RECT MASK 2 28.094 106.38 28.154 107.43 ;
      RECT MASK 2 28.368 106.38 28.428 107.43 ;
      RECT MASK 2 28.642 106.38 28.702 107.43 ;
      RECT MASK 2 28.916 106.38 28.976 107.43 ;
      RECT MASK 2 29.19 106.38 29.25 107.43 ;
      RECT MASK 2 29.464 106.38 29.524 107.43 ;
      RECT MASK 2 29.738 106.38 29.798 107.43 ;
      RECT MASK 2 30.012 106.38 30.072 107.43 ;
      RECT MASK 2 30.286 106.38 30.346 107.43 ;
      RECT MASK 2 30.56 106.38 30.62 107.43 ;
      RECT MASK 2 30.834 106.38 30.894 107.43 ;
      RECT MASK 2 31.108 106.38 31.168 107.43 ;
      RECT MASK 2 31.382 106.38 31.442 107.43 ;
      RECT MASK 2 31.656 106.38 31.716 107.43 ;
      RECT MASK 2 31.93 106.38 31.99 107.43 ;
      RECT MASK 2 32.204 106.38 32.264 107.43 ;
      RECT MASK 2 32.478 106.38 32.538 107.43 ;
      RECT MASK 2 32.752 106.38 32.812 107.43 ;
      RECT MASK 2 33.026 106.38 33.086 107.43 ;
      RECT MASK 2 33.3 106.38 33.36 107.43 ;
      RECT MASK 2 33.574 106.38 33.634 107.43 ;
      RECT MASK 2 33.848 106.38 33.908 107.43 ;
      RECT MASK 2 34.122 106.38 34.182 107.43 ;
      RECT MASK 2 34.396 106.38 34.456 107.43 ;
      RECT MASK 2 34.67 106.38 34.73 107.43 ;
      RECT MASK 2 34.944 106.38 35.004 107.43 ;
      RECT MASK 2 35.218 106.38 35.278 107.43 ;
      RECT MASK 2 35.492 106.38 35.552 107.43 ;
      RECT MASK 2 35.766 106.38 35.826 107.43 ;
      RECT MASK 2 36.04 106.38 36.1 107.43 ;
      RECT MASK 2 36.314 106.38 36.374 107.43 ;
      RECT MASK 2 36.588 106.38 36.648 107.43 ;
      RECT MASK 2 36.862 106.38 36.922 107.43 ;
      RECT MASK 2 37.136 106.38 37.196 107.43 ;
      RECT MASK 2 37.41 106.38 37.47 107.43 ;
      RECT MASK 2 37.684 106.38 37.744 107.43 ;
      RECT MASK 2 37.958 106.38 38.018 107.43 ;
      RECT MASK 2 38.232 106.38 38.292 107.43 ;
      RECT MASK 2 38.506 106.38 38.566 107.43 ;
      RECT MASK 2 38.78 106.38 38.84 107.43 ;
      RECT MASK 2 39.054 106.38 39.114 107.43 ;
      RECT MASK 2 39.328 106.38 39.388 107.43 ;
      RECT MASK 2 39.602 106.38 39.662 107.43 ;
      RECT MASK 2 39.876 106.38 39.936 107.43 ;
      RECT MASK 2 40.15 106.38 40.21 107.43 ;
      RECT MASK 2 40.424 106.38 40.484 107.43 ;
      RECT MASK 2 40.698 106.38 40.758 107.43 ;
      RECT MASK 2 40.972 106.38 41.032 107.43 ;
      RECT MASK 2 41.246 106.38 41.306 107.43 ;
      RECT MASK 2 41.52 106.38 41.58 107.43 ;
      RECT MASK 2 41.794 106.38 41.854 107.43 ;
      RECT MASK 2 42.068 106.38 42.128 107.43 ;
      RECT MASK 2 42.342 106.38 42.402 107.43 ;
      RECT MASK 2 42.616 106.38 42.676 107.43 ;
      RECT MASK 2 42.89 106.38 42.95 107.43 ;
      RECT MASK 2 43.164 106.38 43.224 107.43 ;
      RECT MASK 2 43.438 106.38 43.498 107.43 ;
      RECT MASK 2 45.73 106.38 45.79 107.43 ;
      RECT MASK 2 46.004 106.38 46.064 107.43 ;
      RECT MASK 2 46.278 106.38 46.338 107.43 ;
      RECT MASK 2 46.552 106.38 46.612 107.43 ;
      RECT MASK 2 46.826 106.38 46.886 107.43 ;
      RECT MASK 2 47.1 106.38 47.16 107.43 ;
      RECT MASK 2 47.374 106.38 47.434 107.43 ;
      RECT MASK 2 47.648 106.38 47.708 107.43 ;
      RECT MASK 2 47.922 106.38 47.982 107.43 ;
      RECT MASK 2 48.196 106.38 48.256 107.43 ;
      RECT MASK 2 48.47 106.38 48.53 107.43 ;
      RECT MASK 2 48.744 106.38 48.804 107.43 ;
      RECT MASK 2 49.018 106.38 49.078 107.43 ;
      RECT MASK 2 49.292 106.38 49.352 107.43 ;
      RECT MASK 2 49.566 106.38 49.626 107.43 ;
      RECT MASK 2 49.84 106.38 49.9 107.43 ;
      RECT MASK 2 50.114 106.38 50.174 107.43 ;
      RECT MASK 2 50.388 106.38 50.448 107.43 ;
      RECT MASK 2 50.662 106.38 50.722 107.43 ;
      RECT MASK 2 50.936 106.38 50.996 107.43 ;
      RECT MASK 2 51.21 106.38 51.27 107.43 ;
      RECT MASK 2 51.484 106.38 51.544 107.43 ;
      RECT MASK 2 51.758 106.38 51.818 107.43 ;
      RECT MASK 2 52.032 106.38 52.092 107.43 ;
      RECT MASK 2 52.306 106.38 52.366 107.43 ;
      RECT MASK 2 52.58 106.38 52.64 107.43 ;
      RECT MASK 2 52.854 106.38 52.914 107.43 ;
      RECT MASK 2 53.128 106.38 53.188 107.43 ;
      RECT MASK 2 53.402 106.38 53.462 107.43 ;
      RECT MASK 2 53.676 106.38 53.736 107.43 ;
      RECT MASK 2 53.95 106.38 54.01 107.43 ;
      RECT MASK 2 54.224 106.38 54.284 107.43 ;
      RECT MASK 2 54.498 106.38 54.558 107.43 ;
      RECT MASK 2 54.772 106.38 54.832 107.43 ;
      RECT MASK 2 55.046 106.38 55.106 107.43 ;
      RECT MASK 2 55.32 106.38 55.38 107.43 ;
      RECT MASK 2 55.594 106.38 55.654 107.43 ;
      RECT MASK 2 55.868 106.38 55.928 107.43 ;
      RECT MASK 2 56.142 106.38 56.202 107.43 ;
      RECT MASK 2 56.416 106.38 56.476 107.43 ;
      RECT MASK 2 56.69 106.38 56.75 107.43 ;
      RECT MASK 2 56.964 106.38 57.024 107.43 ;
      RECT MASK 2 57.238 106.38 57.298 107.43 ;
      RECT MASK 2 57.512 106.38 57.572 107.43 ;
      RECT MASK 2 57.786 106.38 57.846 107.43 ;
      RECT MASK 2 58.06 106.38 58.12 107.43 ;
      RECT MASK 2 58.334 106.38 58.394 107.43 ;
      RECT MASK 2 58.608 106.38 58.668 107.43 ;
      RECT MASK 2 58.882 106.38 58.942 107.43 ;
      RECT MASK 2 59.156 106.38 59.216 107.43 ;
      RECT MASK 2 59.43 106.38 59.49 107.43 ;
      RECT MASK 2 59.704 106.38 59.764 107.43 ;
      RECT MASK 2 59.978 106.38 60.038 107.43 ;
      RECT MASK 2 60.252 106.38 60.312 107.43 ;
      RECT MASK 2 60.526 106.38 60.586 107.43 ;
      RECT MASK 2 60.8 106.38 60.86 107.43 ;
      RECT MASK 2 61.074 106.38 61.134 107.43 ;
      RECT MASK 2 61.348 106.38 61.408 107.43 ;
      RECT MASK 2 61.622 106.38 61.682 107.43 ;
      RECT MASK 2 61.896 106.38 61.956 107.43 ;
      RECT MASK 2 62.17 106.38 62.23 107.43 ;
      RECT MASK 2 62.444 106.38 62.504 107.43 ;
      RECT MASK 2 62.718 106.38 62.778 107.43 ;
      RECT MASK 2 62.992 106.38 63.052 107.43 ;
      RECT MASK 2 63.266 106.38 63.326 107.43 ;
      RECT MASK 2 63.54 106.38 63.6 107.43 ;
      RECT MASK 2 63.814 106.38 63.874 107.43 ;
      RECT MASK 2 64.088 106.38 64.148 107.43 ;
      RECT MASK 2 64.362 106.38 64.422 107.43 ;
      RECT MASK 2 64.636 106.38 64.696 107.43 ;
      RECT MASK 2 64.91 106.38 64.97 107.43 ;
      RECT MASK 2 65.184 106.38 65.244 107.43 ;
      RECT MASK 2 65.458 106.38 65.518 107.43 ;
      RECT MASK 2 65.732 106.38 65.792 107.43 ;
      RECT MASK 2 66.006 106.38 66.066 107.43 ;
      RECT MASK 2 66.28 106.38 66.34 107.43 ;
      RECT MASK 2 66.554 106.38 66.614 107.43 ;
      RECT MASK 2 66.828 106.38 66.888 107.43 ;
      RECT MASK 2 67.102 106.38 67.162 107.43 ;
      RECT MASK 2 67.376 106.38 67.436 107.43 ;
      RECT MASK 2 67.65 106.38 67.71 107.43 ;
      RECT MASK 2 67.924 106.38 67.984 107.43 ;
      RECT MASK 2 68.198 106.38 68.258 107.43 ;
      RECT MASK 2 68.472 106.38 68.532 107.43 ;
      RECT MASK 2 68.746 106.38 68.806 107.43 ;
      RECT MASK 2 69.02 106.38 69.08 107.43 ;
      RECT MASK 2 69.294 106.38 69.354 107.43 ;
      RECT MASK 2 69.568 106.38 69.628 107.43 ;
      RECT MASK 2 69.842 106.38 69.902 107.43 ;
      RECT MASK 2 70.116 106.38 70.176 107.43 ;
      RECT MASK 2 70.39 106.38 70.45 107.43 ;
      RECT MASK 2 70.664 106.38 70.724 107.43 ;
      RECT MASK 2 70.938 106.38 70.998 107.43 ;
      RECT MASK 2 71.212 106.38 71.272 107.43 ;
      RECT MASK 2 71.486 106.38 71.546 107.43 ;
      RECT MASK 2 71.76 106.38 71.82 107.43 ;
      RECT MASK 2 72.034 106.38 72.094 107.43 ;
      RECT MASK 2 72.308 106.38 72.368 107.43 ;
      RECT MASK 2 72.582 106.38 72.642 107.43 ;
      RECT MASK 2 72.856 106.38 72.916 107.43 ;
      RECT MASK 2 73.13 106.38 73.19 107.43 ;
      RECT MASK 2 73.404 106.38 73.464 107.43 ;
      RECT MASK 2 73.678 106.38 73.738 107.43 ;
      RECT MASK 2 73.952 106.38 74.012 107.43 ;
      RECT MASK 2 74.226 106.38 74.286 107.43 ;
      RECT MASK 2 74.5 106.38 74.56 107.43 ;
      RECT MASK 2 74.774 106.38 74.834 107.43 ;
      RECT MASK 2 75.048 106.38 75.108 107.43 ;
      RECT MASK 2 75.322 106.38 75.382 107.43 ;
      RECT MASK 2 75.596 106.38 75.656 107.43 ;
      RECT MASK 2 75.87 106.38 75.93 107.43 ;
      RECT MASK 2 76.144 106.38 76.204 107.43 ;
      RECT MASK 2 76.418 106.38 76.478 107.43 ;
      RECT MASK 2 76.692 106.38 76.752 107.43 ;
      RECT MASK 2 76.966 106.38 77.026 107.43 ;
      RECT MASK 2 77.24 106.38 77.3 107.43 ;
      RECT MASK 2 77.514 106.38 77.574 107.43 ;
      RECT MASK 2 77.788 106.38 77.848 107.43 ;
      RECT MASK 2 78.062 106.38 78.122 107.43 ;
      RECT MASK 2 78.336 106.38 78.396 107.43 ;
      RECT MASK 2 78.61 106.38 78.67 107.43 ;
      RECT MASK 2 78.884 106.38 78.944 107.43 ;
      RECT MASK 2 79.158 106.38 79.218 107.43 ;
      RECT MASK 2 79.432 106.38 79.492 107.43 ;
      RECT MASK 2 79.706 106.38 79.766 107.43 ;
      RECT MASK 2 79.98 106.38 80.04 107.43 ;
      RECT MASK 2 80.254 106.38 80.314 107.43 ;
      RECT MASK 2 80.528 106.38 80.588 107.43 ;
      RECT MASK 2 80.802 106.38 80.862 107.43 ;
      RECT MASK 2 81.076 106.38 81.136 107.43 ;
      RECT MASK 2 81.35 106.38 81.41 107.43 ;
      RECT MASK 2 81.624 106.38 81.684 107.43 ;
      RECT MASK 2 81.898 106.38 81.958 107.43 ;
      RECT MASK 2 82.172 106.38 82.232 107.43 ;
      RECT MASK 2 82.446 106.38 82.506 107.43 ;
      RECT MASK 2 82.72 106.38 82.78 107.43 ;
      RECT MASK 2 82.994 106.38 83.054 107.43 ;
      RECT MASK 2 83.268 106.38 83.328 107.43 ;
      RECT MASK 2 83.542 106.38 83.602 107.43 ;
      RECT MASK 2 83.816 106.38 83.876 107.43 ;
      RECT MASK 2 84.09 106.38 84.15 107.43 ;
      RECT MASK 2 84.364 106.38 84.424 107.43 ;
      RECT MASK 2 84.638 106.38 84.698 107.43 ;
      RECT MASK 2 84.912 106.38 84.972 107.43 ;
      RECT MASK 2 85.186 106.38 85.246 107.43 ;
      RECT MASK 2 85.46 106.38 85.52 107.43 ;
      RECT MASK 2 85.734 106.38 85.794 107.43 ;
      RECT MASK 2 86.008 106.38 86.068 107.43 ;
      RECT MASK 2 86.282 106.38 86.342 107.43 ;
      RECT MASK 2 86.556 106.38 86.616 107.43 ;
      RECT MASK 2 86.83 106.38 86.89 107.43 ;
      RECT MASK 2 89.089 106.38 89.149 107.43 ;
      RECT MASK 2 89.363 106.38 89.423 107.43 ;
      RECT MASK 2 89.637 106.38 89.697 107.43 ;
      RECT MASK 2 89.911 106.38 89.971 107.43 ;
      RECT MASK 2 90.185 106.38 90.245 107.43 ;
      RECT MASK 2 90.459 106.38 90.519 107.43 ;
      RECT MASK 2 90.733 106.38 90.793 107.43 ;
      RECT MASK 2 91.007 106.38 91.067 107.43 ;
      RECT MASK 2 91.281 106.38 91.341 107.43 ;
      RECT MASK 2 91.555 106.38 91.615 107.43 ;
      RECT MASK 2 91.829 106.38 91.889 107.43 ;
      RECT MASK 2 92.103 106.38 92.163 107.43 ;
      RECT MASK 2 92.377 106.38 92.437 107.43 ;
      RECT MASK 2 92.651 106.38 92.711 107.43 ;
      RECT MASK 2 92.925 106.38 92.985 107.43 ;
      RECT MASK 2 93.199 106.38 93.259 107.43 ;
      RECT MASK 2 93.473 106.38 93.533 107.43 ;
      RECT MASK 2 93.747 106.38 93.807 107.43 ;
      RECT MASK 2 94.021 106.38 94.081 107.43 ;
      RECT MASK 2 94.295 106.38 94.355 107.43 ;
      RECT MASK 2 94.569 106.38 94.629 107.43 ;
      RECT MASK 2 94.843 106.38 94.903 107.43 ;
      RECT MASK 2 95.117 106.38 95.177 107.43 ;
      RECT MASK 2 95.391 106.38 95.451 107.43 ;
      RECT MASK 2 95.665 106.38 95.725 107.43 ;
      RECT MASK 2 95.939 106.38 95.999 107.43 ;
      RECT MASK 2 96.213 106.38 96.273 107.43 ;
      RECT MASK 2 96.487 106.38 96.547 107.43 ;
      RECT MASK 2 96.761 106.38 96.821 107.43 ;
      RECT MASK 2 97.035 106.38 97.095 107.43 ;
      RECT MASK 2 97.309 106.38 97.369 107.43 ;
      RECT MASK 2 97.583 106.38 97.643 107.43 ;
      RECT MASK 2 97.857 106.38 97.917 107.43 ;
      RECT MASK 2 98.131 106.38 98.191 107.43 ;
      RECT MASK 2 98.405 106.38 98.465 107.43 ;
      RECT MASK 2 98.679 106.38 98.739 107.43 ;
      RECT MASK 2 98.953 106.38 99.013 107.43 ;
      RECT MASK 2 99.227 106.38 99.287 107.43 ;
      RECT MASK 2 99.501 106.38 99.561 107.43 ;
      RECT MASK 2 99.775 106.38 99.835 107.43 ;
      RECT MASK 2 100.049 106.38 100.109 107.43 ;
      RECT MASK 2 100.323 106.38 100.383 107.43 ;
      RECT MASK 2 100.597 106.38 100.657 107.43 ;
      RECT MASK 2 100.871 106.38 100.931 107.43 ;
      RECT MASK 2 101.145 106.38 101.205 107.43 ;
      RECT MASK 2 101.419 106.38 101.479 107.43 ;
      RECT MASK 2 101.693 106.38 101.753 107.43 ;
      RECT MASK 2 101.967 106.38 102.027 107.43 ;
      RECT MASK 2 102.241 106.38 102.301 107.43 ;
      RECT MASK 2 102.515 106.38 102.575 107.43 ;
      RECT MASK 2 102.789 106.38 102.849 107.43 ;
      RECT MASK 2 103.063 106.38 103.123 107.43 ;
      RECT MASK 2 103.337 106.38 103.397 107.43 ;
      RECT MASK 2 103.611 106.38 103.671 107.43 ;
      RECT MASK 2 103.885 106.38 103.945 107.43 ;
      RECT MASK 2 104.159 106.38 104.219 107.43 ;
      RECT MASK 2 104.433 106.38 104.493 107.43 ;
      RECT MASK 2 104.707 106.38 104.767 107.43 ;
      RECT MASK 2 104.981 106.38 105.041 107.43 ;
      RECT MASK 2 105.255 106.38 105.315 107.43 ;
      RECT MASK 2 105.529 106.38 105.589 107.43 ;
      RECT MASK 2 105.803 106.38 105.863 107.43 ;
      RECT MASK 2 106.077 106.38 106.137 107.43 ;
      RECT MASK 2 106.351 106.38 106.411 107.43 ;
      RECT MASK 2 106.625 106.38 106.685 107.43 ;
      RECT MASK 2 106.899 106.38 106.959 107.43 ;
      RECT MASK 2 107.173 106.38 107.233 107.43 ;
      RECT MASK 2 107.447 106.38 107.507 107.43 ;
      RECT MASK 2 107.721 106.38 107.781 107.43 ;
      RECT MASK 2 107.995 106.38 108.055 107.43 ;
      RECT MASK 2 108.269 106.38 108.329 107.43 ;
      RECT MASK 2 108.543 106.38 108.603 107.43 ;
      RECT MASK 2 108.817 106.38 108.877 107.43 ;
      RECT MASK 2 109.091 106.38 109.151 107.43 ;
      RECT MASK 2 109.365 106.38 109.425 107.43 ;
      RECT MASK 2 109.639 106.38 109.699 107.43 ;
      RECT MASK 2 109.913 106.38 109.973 107.43 ;
      RECT MASK 2 110.187 106.38 110.247 107.43 ;
      RECT MASK 2 110.461 106.38 110.521 107.43 ;
      RECT MASK 2 110.735 106.38 110.795 107.43 ;
      RECT MASK 2 111.009 106.38 111.069 107.43 ;
      RECT MASK 2 111.283 106.38 111.343 107.43 ;
      RECT MASK 2 111.557 106.38 111.617 107.43 ;
      RECT MASK 2 111.831 106.38 111.891 107.43 ;
      RECT MASK 2 112.105 106.38 112.165 107.43 ;
      RECT MASK 2 112.379 106.38 112.439 107.43 ;
      RECT MASK 2 112.653 106.38 112.713 107.43 ;
      RECT MASK 2 112.927 106.38 112.987 107.43 ;
      RECT MASK 2 113.201 106.38 113.261 107.43 ;
      RECT MASK 2 113.475 106.38 113.535 107.43 ;
      RECT MASK 2 113.749 106.38 113.809 107.43 ;
      RECT MASK 2 114.023 106.38 114.083 107.43 ;
      RECT MASK 2 114.297 106.38 114.357 107.43 ;
      RECT MASK 2 114.571 106.38 114.631 107.43 ;
      RECT MASK 2 114.845 106.38 114.905 107.43 ;
      RECT MASK 2 115.119 106.38 115.179 107.43 ;
      RECT MASK 2 115.393 106.38 115.453 107.43 ;
      RECT MASK 2 115.667 106.38 115.727 107.43 ;
      RECT MASK 2 115.941 106.38 116.001 107.43 ;
      RECT MASK 2 116.215 106.38 116.275 107.43 ;
      RECT MASK 2 116.489 106.38 116.549 107.43 ;
      RECT MASK 2 116.763 106.38 116.823 107.43 ;
      RECT MASK 2 117.037 106.38 117.097 107.43 ;
      RECT MASK 2 117.311 106.38 117.371 107.43 ;
      RECT MASK 2 117.585 106.38 117.645 107.43 ;
      RECT MASK 2 117.859 106.38 117.919 107.43 ;
      RECT MASK 2 118.133 106.38 118.193 107.43 ;
      RECT MASK 2 118.407 106.38 118.467 107.43 ;
      RECT MASK 2 118.681 106.38 118.741 107.43 ;
      RECT MASK 2 118.955 106.38 119.015 107.43 ;
      RECT MASK 2 119.229 106.38 119.289 107.43 ;
      RECT MASK 2 119.503 106.38 119.563 107.43 ;
      RECT MASK 2 119.777 106.38 119.837 107.43 ;
      RECT MASK 2 120.051 106.38 120.111 107.43 ;
      RECT MASK 2 120.325 106.38 120.385 107.43 ;
      RECT MASK 2 120.599 106.38 120.659 107.43 ;
      RECT MASK 2 120.873 106.38 120.933 107.43 ;
      RECT MASK 2 121.147 106.38 121.207 107.43 ;
      RECT MASK 2 121.421 106.38 121.481 107.43 ;
      RECT MASK 2 121.695 106.38 121.755 107.43 ;
      RECT MASK 2 121.969 106.38 122.029 107.43 ;
      RECT MASK 2 122.243 106.38 122.303 107.43 ;
      RECT MASK 2 122.517 106.38 122.577 107.43 ;
      RECT MASK 2 122.791 106.38 122.851 107.43 ;
      RECT MASK 2 123.065 106.38 123.125 107.43 ;
      RECT MASK 2 123.339 106.38 123.399 107.43 ;
      RECT MASK 2 123.613 106.38 123.673 107.43 ;
      RECT MASK 2 123.887 106.38 123.947 107.43 ;
      RECT MASK 2 124.161 106.38 124.221 107.43 ;
      RECT MASK 2 124.435 106.38 124.495 107.43 ;
      RECT MASK 2 124.709 106.38 124.769 107.43 ;
      RECT MASK 2 124.983 106.38 125.043 107.43 ;
      RECT MASK 2 125.257 106.38 125.317 107.43 ;
      RECT MASK 2 125.531 106.38 125.591 107.43 ;
      RECT MASK 2 125.805 106.38 125.865 107.43 ;
      RECT MASK 2 126.079 106.38 126.139 107.43 ;
      RECT MASK 2 126.353 106.38 126.413 107.43 ;
      RECT MASK 2 126.627 106.38 126.687 107.43 ;
      RECT MASK 2 126.901 106.38 126.961 107.43 ;
      RECT MASK 2 127.175 106.38 127.235 107.43 ;
      RECT MASK 2 127.449 106.38 127.509 107.43 ;
      RECT MASK 2 1.454 107.75 44.382 107.79 ;
      RECT MASK 2 44.846 107.75 87.774 107.79 ;
      RECT MASK 2 88.238 107.75 128.51 107.79 ;
      RECT MASK 2 1.454 107.94 44.382 107.98 ;
      RECT MASK 2 44.846 107.94 87.774 107.98 ;
      RECT MASK 2 88.238 107.94 128.51 107.98 ;
  END
END dwc_ddrphy_vrefglobal

END LIBRARY
