# LEF OUT API 
# Creation Date : Tue Mar 29 15:03:31 IST 2022
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_lpddr5xphy_lstx_acx2_ew
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_lpddr5xphy_lstx_acx2_ew 0 0 ;
  SYMMETRY X Y ;
  SIZE 72.369 BY 74.76 ;
  PIN csrLsTxSlewLPPU0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.07344 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 23.285 0.05 23.323 0.088 ;
    END
  END csrLsTxSlewLPPU0[0]
  PIN csrLsTxSlewLPPU1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.07344 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 23.361 0.05 23.399 0.088 ;
    END
  END csrLsTxSlewLPPU1[0]
  PIN csrLsTxSlewPD0{0}
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.07344 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 23.437 0.05 23.475 0.088 ;
    END
  END csrLsTxSlewPD0[0]
  PIN csrLsTxSlewPD3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.07344 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 23.665 0.05 23.703 0.088 ;
    END
  END csrLsTxSlewPD3[0]
  PIN csrLsTxSlewPD2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.07344 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 23.589 0.05 23.627 0.088 ;
    END
  END csrLsTxSlewPD2[0]
  PIN csrLsTxSlewPD1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.07344 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 23.513 0.05 23.551 0.088 ;
    END
  END csrLsTxSlewPD1[0]
  PIN csrLsTxCalCodePD0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 23.969 0.05 24.007 0.088 ;
    END
  END csrLsTxCalCodePD0[0]
  PIN csrLsTxCalCodePD1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.045 0.05 24.083 0.088 ;
    END
  END csrLsTxCalCodePD1[0]
  PIN csrLsTxCalCodePD2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.121 0.05 24.159 0.088 ;
    END
  END csrLsTxCalCodePD2[0]
  PIN csrLsTxCalCodeLPPU0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.653 74.672 24.691 74.71 ;
    END
  END csrLsTxCalCodeLPPU0[1]
  PIN csrLsTxCalCodeLPPU1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.729 74.672 24.767 74.71 ;
    END
  END csrLsTxCalCodeLPPU1[1]
  PIN csrLsTxCalCodeLPPU2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.805 74.672 24.843 74.71 ;
    END
  END csrLsTxCalCodeLPPU2[1]
  PIN csrLsTxCalCodeLPPU3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.881 74.672 24.919 74.71 ;
    END
  END csrLsTxCalCodeLPPU3[1]
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M10 ;
        RECT 7.2425 41.2625 23.317 41.8625 ;
    END
  END VDDQ
  PIN csrLsReservedP[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.35989775 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 28.165 0.04 28.203 ;
    END
  END csrLsReservedP[0]
  PIN csrLsReservedP[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.353989 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 28.317 0.04 28.355 ;
    END
  END csrLsReservedP[1]
  PIN csrLsReserved[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.310688 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 28.773 0.04 28.811 ;
    END
  END csrLsReserved[1]
  PIN csrLsReservedP[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.341601 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 28.621 0.04 28.659 ;
    END
  END csrLsReservedP[2]
  PIN csrLsReserved[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.293075 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 29.077 0.04 29.115 ;
    END
  END csrLsReserved[2]
  PIN csrLsReserved[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.299896 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 29.229 0.04 29.267 ;
    END
  END csrLsReserved[3]
  PIN VIO_PwrOk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3096 LAYER M10 ;
    ANTENNADIFFAREA 2.09563 LAYER M10 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 4.15908 LAYER M10 ;
      ANTENNAMAXAREACAR 5.3857 LAYER M10 ;
    PORT
      LAYER M10 ;
        RECT 20.104 46.9165 25.62 47.5165 ;
    END
  END VIO_PwrOk
  PIN csrReservedP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 413.493 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.181 0.038 33.219 ;
    END
  END csrReservedP[0]
  PIN csrReservedP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 425.63 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.333 0.038 33.371 ;
    END
  END csrReservedP[1]
  PIN csrReservedP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 411.915 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.485 0.038 33.523 ;
    END
  END csrReservedP[2]
  PIN csrReservedP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 409.296 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.637 0.038 33.675 ;
    END
  END csrReservedP[3]
  PIN csrReserved[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 385.591 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.789 0.038 33.827 ;
    END
  END csrReserved[2]
  PIN csrReserved[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 370.796 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 33.941 0.038 33.979 ;
    END
  END csrReserved[3]
  PIN csrReserved[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 370.561 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 34.397 0.038 34.435 ;
    END
  END csrReserved[1]
  PIN csrLsTxCalCodeLPPU4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.957 74.672 24.995 74.71 ;
    END
  END csrLsTxCalCodeLPPU4[1]
  PIN csrLsTxCalCodeLPPU5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 25.033 74.672 25.071 74.71 ;
    END
  END csrLsTxCalCodeLPPU5[1]
  PIN csrReserved[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 383.709 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 34.245 0.038 34.283 ;
    END
  END csrReserved[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M10 ;
        RECT 7.2425 44.8165 23.317 45.4165 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 35.9425 23.317 36.5425 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 34.1125 23.317 34.7125 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 37.7025 23.317 38.3025 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 46.9165 18.792 47.5165 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 39.4825 23.317 40.0825 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 43.0365 22.7485 43.6365 ;
    END
  END VDD
  PIN LsScan_mode
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.24795 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 34.701 0.038 34.739 ;
    END
  END LsScan_mode
  PIN LsIDDQ_mode
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.255987 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00305975 LAYER M6 ;
      ANTENNAMAXAREACAR 260.144 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.005 0.038 35.043 ;
    END
  END LsIDDQ_mode
  PIN csrLsReserved[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.304779 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 28.925 0.04 28.963 ;
    END
  END csrLsReserved[0]
  PIN csrLsReservedP[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34751 LAYER M6 ;
    ANTENNADIFFAREA 0.00305975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 28.469 0.04 28.507 ;
    END
  END csrLsReservedP[3]
  PIN csrTxSlewPD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 340.214 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.917 0.038 35.955 ;
    END
  END csrTxSlewPD[3]
  PIN csrTxSlewPD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 345.508 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.461 0.038 35.499 ;
    END
  END csrTxSlewPD[0]
  PIN csrTxSlewPD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 340.253 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.613 0.038 35.651 ;
    END
  END csrTxSlewPD[1]
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M10 ;
        RECT 7.2425 34.9925 23.317 35.5925 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 43.9165 23.317 44.5165 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 40.3625 23.317 40.9625 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 46.0165 23.317 46.6165 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 42.1365 23.317 42.7365 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 36.8225 23.317 37.4225 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 38.5825 23.317 39.1825 ;
    END
    PORT
      LAYER M10 ;
        RECT 7.2425 33.1625 23.317 33.7625 ;
    END
  END VSS
  PIN csrTxSlewPD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 348.449 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 35.765 0.038 35.803 ;
    END
  END csrTxSlewPD[2]
  PIN csrTxCalCodePD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 375.273 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.677 0.038 36.715 ;
    END
  END csrTxCalCodePD[2]
  PIN scan_shift
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 365.508 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.221 0.038 36.259 ;
    END
  END scan_shift
  PIN csrTxCalCodePD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 346.018 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.373 0.038 36.411 ;
    END
  END csrTxCalCodePD[0]
  PIN csrTxCalCodePD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 355.018 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.981 0.038 37.019 ;
    END
  END csrTxCalCodePD[3]
  PIN csrTxCalCodePD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 387.881 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.525 0.038 36.563 ;
    END
  END csrTxCalCodePD[1]
  PIN csrTxCalCodePD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 351.057 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 37.133 0.038 37.171 ;
    END
  END csrTxCalCodePD[4]
  PIN csrTxCalCodePD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 372.293 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 37.437 0.038 37.475 ;
    END
  END csrTxCalCodePD[6]
  PIN scan_shift_cg
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 352.279 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.045 0.038 38.083 ;
    END
  END scan_shift_cg
  PIN CalUpdate
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.248292 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 442.275 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 37.893 0.038 37.931 ;
    END
  END CalUpdate
  PIN scan_si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 387.103 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 40.477 0.038 40.515 ;
    END
  END scan_si
  PIN csrTxCalCodePU[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 380.668 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.653 0.038 38.691 ;
    END
  END csrTxCalCodePU[8]
  PIN csrTxSlewPU[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 348.567 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 41.389 0.038 41.427 ;
    END
  END csrTxSlewPU[3]
  PIN csrTxSlewPU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 340.665 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 41.237 0.038 41.275 ;
    END
  END csrTxSlewPU[2]
  PIN csrTxCalCodePU[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 362.038 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 39.413 0.038 39.451 ;
    END
  END csrTxCalCodePU[5]
  PIN csrTxCalCodePU[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 363.335 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.957 0.038 38.995 ;
    END
  END csrTxCalCodePU[7]
  PIN csrTxCalCodePU[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 358.096 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.805 0.038 38.843 ;
    END
  END csrTxCalCodePU[6]
  PIN csrTxCalCodePD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 384.685 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 37.285 0.038 37.323 ;
    END
  END csrTxCalCodePD[5]
  PIN Dficlk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 363.077 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.501 0.038 38.539 ;
    END
  END Dficlk
  PIN scan_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00611975 LAYER M6 ;
      ANTENNAMAXAREACAR 84.04059975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 36.069 0.038 36.107 ;
    END
  END scan_mode
  PIN scan_so
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNADIFFAREA 0.00611975 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.273 0.038 38.311 ;
    END
  END scan_so
  PIN csrTxCalCodePU[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 377.469 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 39.261 0.038 39.299 ;
    END
  END csrTxCalCodePU[4]
  PIN csrTxCalCodePU[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 370.469 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 39.717 0.038 39.755 ;
    END
  END csrTxCalCodePU[3]
  PIN csrTxCalCodePU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 350.978 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 40.325 0.038 40.363 ;
    END
  END csrTxCalCodePU[1]
  PIN ResetAsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00204 LAYER M6 ;
      ANTENNAMAXAREACAR 179.472 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.197 0.038 38.235 ;
    END
  END ResetAsync
  PIN IDDQ_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00408 LAYER M6 ;
      ANTENNAMAXAREACAR 173.92 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 40.629 0.038 40.667 ;
    END
  END IDDQ_mode
  PIN csrTxSlewPU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 350.743 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 40.781 0.038 40.819 ;
    END
  END csrTxSlewPU[0]
  PIN csrTxSlewPU[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 348.135 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 41.085 0.038 41.123 ;
    END
  END csrTxSlewPU[1]
  PIN csrTxCalCodePD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 352.707 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 37.741 0.038 37.779 ;
    END
  END csrTxCalCodePD[7]
  PIN csrTxCalCodePU[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 378.312 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 40.173 0.038 40.211 ;
    END
  END csrTxCalCodePU[0]
  PIN csrTxCalCodePU[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 370.939 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 39.565 0.038 39.603 ;
    END
  END csrTxCalCodePU[2]
  PIN csrTxCalCodePD[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.267254 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 351.883 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 38.349 0.038 38.387 ;
    END
  END csrTxCalCodePD[8]
  PIN csrLsTxCalCodeLPPU6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 25.109 74.672 25.147 74.71 ;
    END
  END csrLsTxCalCodeLPPU6[1]
  PIN csrLsTxCalCodePD3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.197 0.05 24.235 0.088 ;
    END
  END csrLsTxCalCodePD3[0]
  PIN csrLsTxCalCodePD4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.273 0.05 24.311 0.088 ;
    END
  END csrLsTxCalCodePD4[0]
  PIN csrLsTxCalCodePD5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.349 0.05 24.387 0.088 ;
    END
  END csrLsTxCalCodePD5[0]
  PIN csrLsTxCalCodePD6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.425 0.05 24.463 0.088 ;
    END
  END csrLsTxCalCodePD6[0]
  PIN csrLsTxCalCodePD7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.501 0.05 24.539 0.088 ;
    END
  END csrLsTxCalCodePD7[0]
  PIN csrLsTxCalCodePD8[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.577 0.05 24.615 0.088 ;
    END
  END csrLsTxCalCodePD8[0]
  PIN csrLsTxCalCodeLPPU7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 25.185 0.05 25.223 0.088 ;
    END
  END csrLsTxCalCodeLPPU7[0]
  PIN csrLsTxCalCodeLPPU8[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 25.261 0.05 25.299 0.088 ;
    END
  END csrLsTxCalCodeLPPU8[0]
  PIN csrLsTxCalCodeLPPU6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 25.109 0.05 25.147 0.088 ;
    END
  END csrLsTxCalCodeLPPU6[0]
  PIN csrLsTxCalCodeLPPU8[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 25.261 74.672 25.299 74.71 ;
    END
  END csrLsTxCalCodeLPPU8[1]
  PIN csrLsTxSlewPD1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 23.513 74.672 23.551 74.71 ;
    END
  END csrLsTxSlewPD1[1]
  PIN csrLsTxSlewPD2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 23.589 74.672 23.627 74.71 ;
    END
  END csrLsTxSlewPD2[1]
  PIN csrLsTxSlewPD3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 23.665 74.672 23.703 74.71 ;
    END
  END csrLsTxSlewPD3[1]
  PIN csrLsTxCalCodePD8[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.577 74.672 24.615 74.71 ;
    END
  END csrLsTxCalCodePD8[1]
  PIN csrLsTxCalCodePD7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.501 74.672 24.539 74.71 ;
    END
  END csrLsTxCalCodePD7[1]
  PIN csrLsTxCalCodePD1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.045 74.672 24.083 74.71 ;
    END
  END csrLsTxCalCodePD1[1]
  PIN csrLsTxCalCodePD2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.121 74.672 24.159 74.71 ;
    END
  END csrLsTxCalCodePD2[1]
  PIN csrLsTxCalCodePD3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.197 74.672 24.235 74.71 ;
    END
  END csrLsTxCalCodePD3[1]
  PIN csrLsTxCalCodePD4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.273 74.672 24.311 74.71 ;
    END
  END csrLsTxCalCodePD4[1]
  PIN csrLsTxCalCodePD5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.349 74.672 24.387 74.71 ;
    END
  END csrLsTxCalCodePD5[1]
  PIN csrLsTxCalCodePD6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 24.425 74.672 24.463 74.71 ;
    END
  END csrLsTxCalCodePD6[1]
  PIN csrLsTxCalCodeLPPU5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 25.033 0.05 25.071 0.088 ;
    END
  END csrLsTxCalCodeLPPU5[0]
  PIN csrLsTxCalCodeLPPU4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.957 0.05 24.995 0.088 ;
    END
  END csrLsTxCalCodeLPPU4[0]
  PIN csrLsTxCalCodeLPPU3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.881 0.05 24.919 0.088 ;
    END
  END csrLsTxCalCodeLPPU3[0]
  PIN csrLsTxCalCodeLPPU7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 25.185 74.672 25.223 74.71 ;
    END
  END csrLsTxCalCodeLPPU7[1]
  PIN BurnIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.457482 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.00102 LAYER M6 ;
      ANTENNAMAXAREACAR 739.753 LAYER M6 ;
    PORT
      LAYER M6 ;
        RECT 0 27.557 0.04 27.595 ;
    END
  END BurnIn
  PIN LsPwrOkVDD[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 22.905 74.672 22.943 74.71 ;
    END
  END LsPwrOkVDD[1]
  PIN csrLsTxCalCodeLPPU2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.805 0.05 24.843 0.088 ;
    END
  END csrLsTxCalCodeLPPU2[0]
  PIN csrLsTxSlewPD0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 23.437 74.672 23.475 74.71 ;
    END
  END csrLsTxSlewPD0[1]
  PIN csrLsTxCalCodeLPPU1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.729 0.05 24.767 0.088 ;
    END
  END csrLsTxCalCodeLPPU1[0]
  PIN csrLsTxSlewLPPU1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 23.361 74.672 23.399 74.71 ;
    END
  END csrLsTxSlewLPPU1[1]
  PIN csrLsTxCalCodeLPPU0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.11016 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 24.653 0.05 24.691 0.088 ;
    END
  END csrLsTxCalCodeLPPU0[0]
  PIN csrLsTxSlewLPPU0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 23.285 74.672 23.323 74.71 ;
    END
  END csrLsTxSlewLPPU0[1]
  PIN csrLsTxSlewLPPU2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.07344 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 23.209 0.05 23.247 0.088 ;
    END
  END csrLsTxSlewLPPU2[0]
  PIN csrLsTxSlewLPPU2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 23.209 74.672 23.247 74.71 ;
    END
  END csrLsTxSlewLPPU2[1]
  PIN LsPwrOkVDD[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83708 LAYER M7 ;
    ANTENNADIFFAREA 0.44064 LAYER M7 ;
    PORT
      LAYER M7 ;
        RECT 22.905 0.05 22.943 0.088 ;
    END
  END LsPwrOkVDD[0]
  PIN csrLsTxCalCodePD0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M7 ;
        RECT 23.969 74.672 24.007 74.71 ;
    END
  END csrLsTxCalCodePD0[1]
  OBS
    LAYER M0 SPACING 0 ;
      RECT MASK 1 0 0 72.369 74.76 ;
    LAYER M1 SPACING 0 ;
      RECT MASK 1 0 0 72.369 74.76 ;
    LAYER M0 SPACING 0 ;
      RECT MASK 2 0 0 72.369 74.76 ;
    LAYER M1 SPACING 0 ;
      RECT MASK 2 0 0 72.369 74.76 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 1 0 0 72.369 74.76 ;
    LAYER M3 SPACING 0 ;
      RECT MASK 1 0 0 72.369 74.76 ;
    LAYER M2 SPACING 0 ;
      RECT MASK 2 0 0 72.369 74.76 ;
    LAYER M5 SPACING 0 ;
      RECT 0 0 72.369 74.76 ;
    LAYER M3 SPACING 0 ;
      RECT MASK 2 0 0 72.369 74.76 ;
    LAYER M4 SPACING 0 ;
      RECT MASK 1 0 0 72.369 74.76 ;
    LAYER M6 SPACING 0 ;
      POLYGON 72.369 0 72.369 74.76 0 74.76 0 41.427 0.038 41.427 0.038 41.389 0 41.389 0 41.275 0.038 41.275 0.038 41.237 0 41.237 0 41.123 0.038 41.123 0.038 41.085 0 41.085 0 40.819 0.038 40.819 0.038 40.781 0 40.781 0 40.667 0.038 40.667 0.038 40.629 0 40.629 0 40.515 0.038 40.515 0.038 40.477 0 40.477 0 40.363 0.038 40.363 0.038 40.325 0 40.325 0 40.211 0.038 40.211 0.038 40.173 0 40.173 0 39.755 0.038 39.755 0.038 39.717 0 39.717 0 39.603 0.038 39.603 0.038 39.565 0 39.565 0 39.451 0.038 39.451 0.038 39.413 0 39.413 0 39.299 0.038 39.299 0.038 39.261 0 39.261 0 38.995 0.038 38.995 0.038 38.957 0 38.957 0 38.843 0.038 38.843 0.038 38.805 0 38.805 0 38.691 0.038 38.691 0.038 38.653 0 38.653 0 38.539 0.038 38.539 0.038 38.501 0 38.501 0 38.387 0.038 38.387 0.038 38.349 0 38.349 0 38.311 0.038 38.311 0.038 38.273 0 38.273 0 38.235 0.038 38.235 0.038 38.197 0 38.197 0 38.083 0.038 38.083 0.038 38.045 0 38.045 0 37.931 0.038 37.931 0.038 37.893 0 37.893 0 37.779 0.038 37.779 0.038 37.741 0 37.741 0 37.475 0.038 37.475 0.038 37.437 0 37.437 0 37.323 0.038 37.323 0.038 37.285 0 37.285 0 37.171 0.038 37.171 0.038 37.133 0 37.133 0 37.019 0.038 37.019 0.038 36.981 0 36.981 0 36.715 0.038 36.715 0.038 36.677 0 36.677 0 36.563 0.038 36.563 0.038 36.525 0 36.525 0 36.411 0.038 36.411 0.038 36.373 0 36.373 0 36.259 0.038 36.259 0.038 36.221 0 36.221 0 36.107 0.038 36.107 0.038 36.069 0 36.069 0 35.955 0.038 35.955 0.038 35.917 0 35.917 0 35.803 0.038 35.803 0.038 35.765 0 35.765 0 35.651 0.038 35.651 0.038 35.613 0 35.613 0 35.499 0.038 35.499 0.038 35.461 0 35.461 0 35.043 0.038 35.043 0.038 35.005 0 35.005 0 34.739 0.038 34.739 0.038 34.701 0 34.701 0 34.435 0.038 34.435 0.038 34.397 0 34.397 0 34.283 0.038 34.283 0.038 34.245 0 34.245 0 33.979 0.038 33.979 0.038 33.941 0 33.941 0 33.827 0.038 33.827 0.038 33.789 0 33.789 0 33.675 0.038 33.675 0.038 33.637 0 33.637 0 33.523 0.038 33.523 0.038 33.485 0 33.485 0 33.371 0.038 33.371 0.038 33.333 0 33.333 0 33.219 0.038 33.219 0.038 33.181 0 33.181 0 29.267 0.04 29.267 0.04 29.229 0 29.229 0 29.115 0.04 29.115 0.04 29.077 0 29.077 0 28.963 0.04 28.963 0.04 28.925 0 28.925 0 28.811 0.04 28.811 0.04 28.773 0 28.773 0 28.659 0.04 28.659 0.04 28.621 0 28.621 0 28.507 0.04 28.507 0.04 28.469 0 28.469 0 28.355 0.04 28.355 0.04 28.317 0 28.317 0 28.203 0.04 28.203 0.04 28.165 0 28.165 0 27.595 0.04 27.595 0.04 27.557 0 27.557 0 0 ;
    LAYER M4 SPACING 0 ;
      RECT MASK 2 0 0 72.369 74.76 ;
    LAYER M7 SPACING 0 ;
      POLYGON 0 0 0 74.76 72.369 74.76 72.369 74.71 22.905 74.71 22.905 74.672 22.943 74.672 22.943 74.71 23.209 74.71 23.209 74.672 23.247 74.672 23.247 74.71 23.285 74.71 23.285 74.672 23.323 74.672 23.323 74.71 23.361 74.71 23.361 74.672 23.399 74.672 23.399 74.71 23.437 74.71 23.437 74.672 23.475 74.672 23.475 74.71 23.513 74.71 23.513 74.672 23.551 74.672 23.551 74.71 23.589 74.71 23.589 74.672 23.627 74.672 23.627 74.71 23.665 74.71 23.665 74.672 23.703 74.672 23.703 74.71 23.969 74.71 23.969 74.672 24.007 74.672 24.007 74.71 24.045 74.71 24.045 74.672 24.083 74.672 24.083 74.71 24.121 74.71 24.121 74.672 24.159 74.672 24.159 74.71 24.197 74.71 24.197 74.672 24.235 74.672 24.235 74.71 24.273 74.71 24.273 74.672 24.311 74.672 24.311 74.71 24.349 74.71 24.349 74.672 24.387 74.672 24.387 74.71 24.425 74.71 24.425 74.672 24.463 74.672 24.463 74.71 24.501 74.71 24.501 74.672 24.539 74.672 24.539 74.71 24.577 74.71 24.577 74.672 24.615 74.672 24.615 74.71 24.653 74.71 24.653 74.672 24.691 74.672 24.691 74.71 24.729 74.71 24.729 74.672 24.767 74.672 24.767 74.71 24.805 74.71 24.805 74.672 24.843 74.672 24.843 74.71 24.881 74.71 24.881 74.672 24.919 74.672 24.919 74.71 24.957 74.71 24.957 74.672 24.995 74.672 24.995 74.71 25.033 74.71 25.033 74.672 25.071 74.672 25.071 74.71 25.109 74.71 25.109 74.672 25.147 74.672 25.147 74.71 25.185 74.71 25.185 74.672 25.223 74.672 25.223 74.71 25.261 74.71 25.261 74.672 25.299 74.672 25.299 74.71 72.369 74.71 72.369 0.088 22.905 0.088 22.905 0.05 22.943 0.05 22.943 0.088 23.209 0.088 23.209 0.05 23.247 0.05 23.247 0.088 23.285 0.088 23.285 0.05 23.323 0.05 23.323 0.088 23.361 0.088 23.361 0.05 23.399 0.05 23.399 0.088 23.437 0.088 23.437 0.05 23.475 0.05 23.475 0.088 23.513 0.088 23.513 0.05 23.551 0.05 23.551 0.088 23.589 0.088 23.589 0.05 23.627 0.05 23.627 0.088 23.665 0.088 23.665 0.05 23.703 0.05 23.703 0.088 23.969 0.088 23.969 0.05 24.007 0.05 24.007 0.088 24.045 0.088 24.045 0.05 24.083 0.05 24.083 0.088 24.121 0.088 24.121 0.05 24.159 0.05 24.159 0.088 24.197 0.088 24.197 0.05 24.235 0.05 24.235 0.088 24.273 0.088 24.273 0.05 24.311 0.05 24.311 0.088 24.349 0.088 24.349 0.05 24.387 0.05 24.387 0.088 24.425 0.088 24.425 0.05 24.463 0.05 24.463 0.088 24.501 0.088 24.501 0.05 24.539 0.05 24.539 0.088 24.577 0.088 24.577 0.05 24.615 0.05 24.615 0.088 24.653 0.088 24.653 0.05 24.691 0.05 24.691 0.088 24.729 0.088 24.729 0.05 24.767 0.05 24.767 0.088 24.805 0.088 24.805 0.05 24.843 0.05 24.843 0.088 24.881 0.088 24.881 0.05 24.919 0.05 24.919 0.088 24.957 0.088 24.957 0.05 24.995 0.05 24.995 0.088 25.033 0.088 25.033 0.05 25.071 0.05 25.071 0.088 25.109 0.088 25.109 0.05 25.147 0.05 25.147 0.088 25.185 0.088 25.185 0.05 25.223 0.05 25.223 0.088 25.261 0.088 25.261 0.05 25.299 0.05 25.299 0.088 72.369 0.088 72.369 0 ;
    LAYER M8 SPACING 0 ;
      RECT 0 0 72.369 74.76 ;
    LAYER M9 SPACING 0 ;
      RECT 0 0 72.369 74.76 ;
    LAYER M10 SPACING 0 ;
      POLYGON 0 0 0 74.76 72.369 74.76 72.369 47.5165 7.2425 47.5165 7.2425 46.9165 18.792 46.9165 18.792 47.5165 20.104 47.5165 20.104 46.9165 25.62 46.9165 25.62 47.5165 72.369 47.5165 72.369 46.6165 7.2425 46.6165 7.2425 46.0165 23.317 46.0165 23.317 46.6165 72.369 46.6165 72.369 45.4165 7.2425 45.4165 7.2425 44.8165 23.317 44.8165 23.317 45.4165 72.369 45.4165 72.369 44.5165 7.2425 44.5165 7.2425 43.9165 23.317 43.9165 23.317 44.5165 72.369 44.5165 72.369 43.6365 7.2425 43.6365 7.2425 43.0365 22.7485 43.0365 22.7485 43.6365 72.369 43.6365 72.369 42.7365 7.2425 42.7365 7.2425 42.1365 23.317 42.1365 23.317 42.7365 72.369 42.7365 72.369 41.8625 7.2425 41.8625 7.2425 41.2625 23.317 41.2625 23.317 41.8625 72.369 41.8625 72.369 40.9625 7.2425 40.9625 7.2425 40.3625 23.317 40.3625 23.317 40.9625 72.369 40.9625 72.369 40.0825 7.2425 40.0825 7.2425 39.4825 23.317 39.4825 23.317 40.0825 72.369 40.0825 72.369 39.1825 7.2425 39.1825 7.2425 38.5825 23.317 38.5825 23.317 39.1825 72.369 39.1825 72.369 38.3025 7.2425 38.3025 7.2425 37.7025 23.317 37.7025 23.317 38.3025 72.369 38.3025 72.369 37.4225 7.2425 37.4225 7.2425 36.8225 23.317 36.8225 23.317 37.4225 72.369 37.4225 72.369 36.5425 7.2425 36.5425 7.2425 35.9425 23.317 35.9425 23.317 36.5425 72.369 36.5425 72.369 35.5925 7.2425 35.5925 7.2425 34.9925 23.317 34.9925 23.317 35.5925 72.369 35.5925 72.369 34.7125 7.2425 34.7125 7.2425 34.1125 23.317 34.1125 23.317 34.7125 72.369 34.7125 72.369 33.7625 7.2425 33.7625 7.2425 33.1625 23.317 33.1625 23.317 33.7625 72.369 33.7625 72.369 0 ;
  END
END dwc_lpddr5xphy_lstx_acx2_ew

END LIBRARY
