.subckt abutment_acx4_a0_aM_aM_a0_ew
.ends abutment_acx4_a0_aM_aM_a0_ew
