# LEF OUT API 
# Creation Date : Thu May 12 04:30:06 PDT 2022
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO dwc_ddrphy_txrxac_ns
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dwc_ddrphy_txrxac_ns 0 0 ;
  SYMMETRY X Y ;
  SIZE 38.16 BY 241.65 ;
  PIN CsrTxChargeCancel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1206.6 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5408.68 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.813 37.98 213.853 ;
    END
  END CsrTxChargeCancel[3]
  PIN CsrTxChargeCancel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1199.89 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5380.21 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.653 37.98 213.693 ;
    END
  END CsrTxChargeCancel[2]
  PIN CsrTxChargeCancel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1201.11 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5385.56 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.493 37.98 213.533 ;
    END
  END CsrTxChargeCancel[1]
  PIN CsrTxChargeCancel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1185.47 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5328.31 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.333 37.98 213.373 ;
    END
  END CsrTxChargeCancel[0]
  PIN CsrTxCalBaseN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1260.31 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5640.32 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 202.508 37.98 202.548 ;
    END
  END CsrTxCalBaseN
  PIN atpg_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.24564 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.56709 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0375839375 LAYER D6 ;
      ANTENNAMAXAREACAR 275.845 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 652.01 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 20.3955 0 20.4755 0.08 ;
    END
  END atpg_mode
  PIN VREFA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.051 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 3.48196 LAYER D8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 23.3688 LAYER D8 ;
      ANTENNAMAXAREACAR 9.29188 LAYER D8 ;
      ANTENNAMAXSIDEAREACAR 5.42132 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 0.6 4.6 19.24425 5.3 ;
    END
  END VREFA
  PIN VIO_TIE_LO_VREFA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 1.026 LAYER D8 ;
    ANTENNADIFFAREA 0.08064 LAYER D8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0588 LAYER D8 ;
      ANTENNAMAXAREACAR 110.706 LAYER D8 ;
      ANTENNAMAXSIDEAREACAR 47.4331 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 19.6305 4.6 24.6305 5.3 ;
    END
  END VIO_TIE_LO_VREFA
  PIN RxRcvDataOdd
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.06518 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.161055 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 2.3135 0 2.3935 0.08 ;
    END
  END RxRcvDataOdd
  PIN RxRcvDataEven
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.08278 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.200655 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 2.4585 0 2.5385 0.08 ;
    END
  END RxRcvDataEven
  PIN RxPowerdown
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05638 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.141255 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 478.903 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 1191.04 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 2.7485 0 2.8285 0.08 ;
    END
  END RxPowerdown
  PIN RxCoreLoopEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.83 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8818999375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0518399375 LAYER D6 ;
      ANTENNAMAXAREACAR 224.698 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 781.095 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 20.2505 0 20.3305 0.08 ;
    END
  END RxCoreLoopEn
  PIN RxClkX
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.04758 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.121455 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D6 ;
      ANTENNAMAXAREACAR 241.383 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 574.417 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 2.6035 0 2.6835 0.08 ;
    END
  END RxClkX
  PIN RxClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.02998 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081855 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D6 ;
      ANTENNAMAXAREACAR 242.222 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 592.722 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 2.8935 0 2.9735 0.08 ;
    END
  END RxClk
  PIN FlyOverEnRx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07596 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.18531 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 161.414 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 355.875 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 7.616 0 7.696 0.08 ;
    END
  END FlyOverEnRx
  PIN FlyOverDataRx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.17208 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.65158 LAYER D6 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.0655 0 28.1455 0.08 ;
    END
  END FlyOverDataRx
  PIN TxPowerdown{1}
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18832 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.43812 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 175.297 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 451.445 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 29.1205 0 29.2005 0.08 ;
    END
  END TxPowerdown[1]
  PIN TxPowerdown[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 170.079 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 427.389 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.9755 0 29.0555 0.08 ;
    END
  END TxPowerdown[0]
  PIN TxEq
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.34552 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7918199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0259199375 LAYER D6 ;
      ANTENNAMAXAREACAR 24.9867 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 69.9385 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.6855 0 28.7655 0.08 ;
    END
  END TxEq
  PIN TxEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.30232 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.69462 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0259199375 LAYER D6 ;
      ANTENNAMAXAREACAR 20.5081 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 56.348 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.8305 0 28.9105 0.08 ;
    END
  END TxEn
  PIN TxDat
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.17272 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40302 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.020736 LAYER D6 ;
      ANTENNAMAXAREACAR 25.217 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 85.599 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.7755 0 25.8555 0.08 ;
    END
  END TxDat
  PIN TxClk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23752 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5488199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.011664 LAYER D6 ;
      ANTENNAMAXAREACAR 54.2725 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 163.442 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 28.2105 0 28.2905 0.08 ;
    END
  END TxClk
  PIN FlyOverTriTx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D6 ;
      ANTENNAMAXAREACAR 96.573099938 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 250.576 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.9205 0 28.0005 0.08 ;
    END
  END FlyOverTriTx
  PIN FlyOverEnTx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.17276 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40311 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 176.982 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 492.035 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 24.5755 0 24.6555 0.08 ;
    END
  END FlyOverEnTx
  PIN FlyOverDataTx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 191.853 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 498.611 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.7755 0 27.8555 0.08 ;
    END
  END FlyOverDataTx
  PIN Ctlpipe_ODT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1592399375 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.37269 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D6 ;
      ANTENNAMAXAREACAR 164.825 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 504.143 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 26.9755 0 27.0555 0.08 ;
    END
  END Ctlpipe_ODT
  PIN CsrTxStrenEqLo480Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18832 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.43812 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 101.298 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 224.406 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.4855 0 27.5655 0.08 ;
    END
  END CsrTxStrenEqLo480Pu
  PIN CsrTxStrenEqLo480Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.4983 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.922 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 29.4105 0 29.4905 0.08 ;
    END
  END CsrTxStrenEqLo480Pd
  PIN CsrTxStrenEqLo240Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18832 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.43812 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 101.298 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 224.406 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 26.2855 0 26.3655 0.08 ;
    END
  END CsrTxStrenEqLo240Pu
  PIN CsrTxStrenEqLo240Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.440399937 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.661 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 30.6105 0 30.6905 0.08 ;
    END
  END CsrTxStrenEqLo240Pd
  PIN CsrTxStrenEqLo120Pu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 101.183 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 224.146 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 21.4855 0 21.5655 0.08 ;
    END
  END CsrTxStrenEqLo120Pu[3]
  PIN CsrTxStrenEqLo120Pu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 101.183 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 224.146 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 22.6855 0 22.7655 0.08 ;
    END
  END CsrTxStrenEqLo120Pu[2]
  PIN CsrTxStrenEqLo120Pu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 101.183 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 224.146 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 23.8855 0 23.9655 0.08 ;
    END
  END CsrTxStrenEqLo120Pu[1]
  PIN CsrTxStrenEqLo120Pu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 101.183 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 224.146 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.0855 0 25.1655 0.08 ;
    END
  END CsrTxStrenEqLo120Pu[0]
  PIN CsrTxStrenEqLo120Pd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.440399937 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.661 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 35.4105 0 35.4905 0.08 ;
    END
  END CsrTxStrenEqLo120Pd[3]
  PIN CsrTxStrenEqLo120Pd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.440399937 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.661 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 34.2105 0 34.2905 0.08 ;
    END
  END CsrTxStrenEqLo120Pd[2]
  PIN CsrTxStrenEqLo120Pd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.440399937 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.661 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.0105 0 33.0905 0.08 ;
    END
  END CsrTxStrenEqLo120Pd[1]
  PIN CsrTxStrenEqLo120Pd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.440399937 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.661 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 31.8105 0 31.8905 0.08 ;
    END
  END CsrTxStrenEqLo120Pd[0]
  PIN CsrTxStrenEqHi480Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 103.595 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 237.906 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 26.8305 0 26.9105 0.08 ;
    END
  END CsrTxStrenEqHi480Pu
  PIN CsrTxStrenEqHi480Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.5827 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.305 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 29.2655 0 29.3455 0.08 ;
    END
  END CsrTxStrenEqHi480Pd
  PIN CsrTxStrenEqHi240Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 103.595 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 237.906 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.6305 0 25.7105 0.08 ;
    END
  END CsrTxStrenEqHi240Pu
  PIN CsrTxStrenEqHi240Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.5827 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.305 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 30.4655 0 30.5455 0.08 ;
    END
  END CsrTxStrenEqHi240Pd
  PIN CsrTxStrenEqHi120Pu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 103.595 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 237.906 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 20.8305 0 20.9105 0.08 ;
    END
  END CsrTxStrenEqHi120Pu[3]
  PIN CsrTxStrenEqHi120Pu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 103.595 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 237.906 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 22.0305 0 22.1105 0.08 ;
    END
  END CsrTxStrenEqHi120Pu[2]
  PIN CsrTxStrenEqHi120Pu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 103.595 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 237.906 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 23.2305 0 23.3105 0.08 ;
    END
  END CsrTxStrenEqHi120Pu[1]
  PIN CsrTxStrenEqHi120Pu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.003456 LAYER D6 ;
      ANTENNAMAXAREACAR 103.595 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 237.906 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 24.4305 0 24.5105 0.08 ;
    END
  END CsrTxStrenEqHi120Pu[0]
  PIN CsrTxStrenEqHi120Pd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.5827 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.305 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 35.2655 0 35.3455 0.08 ;
    END
  END CsrTxStrenEqHi120Pd[3]
  PIN CsrTxStrenEqHi120Pd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.5827 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.305 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 34.0655 0 34.1455 0.08 ;
    END
  END CsrTxStrenEqHi120Pd[2]
  PIN CsrTxStrenEqHi120Pd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.5827 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.305 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.8655 0 32.9455 0.08 ;
    END
  END CsrTxStrenEqHi120Pd[1]
  PIN CsrTxStrenEqHi120Pd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006912 LAYER D6 ;
      ANTENNAMAXAREACAR 49.5827 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 114.305 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 31.6655 0 31.7455 0.08 ;
    END
  END CsrTxStrenEqHi120Pd[0]
  PIN CsrTxStren480Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 60.7449 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 145.448 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 26.6855 0 26.7655 0.08 ;
    END
  END CsrTxStren480Pu
  PIN CsrTxStren480Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18832 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.43812 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 41.9082 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 98.0524 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 30.0655 0 30.1455 0.08 ;
    END
  END CsrTxStren480Pd
  PIN CsrTxStren240Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 60.7449 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 145.448 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.4855 0 25.5655 0.08 ;
    END
  END CsrTxStren240Pu
  PIN CsrTxStren240Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18832 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.43812 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 41.9082 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 98.0524 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 31.2655 0 31.3455 0.08 ;
    END
  END CsrTxStren240Pd
  PIN CsrTxStren120Pu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 60.7449 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 145.448 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 20.6855 0 20.7655 0.08 ;
    END
  END CsrTxStren120Pu[3]
  PIN CsrTxStren120Pu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 60.7449 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 145.448 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 21.8855 0 21.9655 0.08 ;
    END
  END CsrTxStren120Pu[2]
  PIN CsrTxStren120Pu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 60.7449 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 145.448 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 23.0855 0 23.1655 0.08 ;
    END
  END CsrTxStren120Pu[1]
  PIN CsrTxStren120Pu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.006048 LAYER D6 ;
      ANTENNAMAXAREACAR 60.7449 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 145.448 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 24.2855 0 24.3655 0.08 ;
    END
  END CsrTxStren120Pu[0]
  PIN CsrTxStren120Pd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 41.8661 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 97.9577 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 36.0655 0 36.1455 0.08 ;
    END
  END CsrTxStren120Pd[3]
  PIN CsrTxStren120Pd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 41.8661 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 97.9577 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 34.8655 0 34.9455 0.08 ;
    END
  END CsrTxStren120Pd[2]
  PIN CsrTxStren120Pd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 41.8661 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 97.9577 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.6655 0 33.7455 0.08 ;
    END
  END CsrTxStren120Pd[1]
  PIN CsrTxStren120Pd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18792 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4372199375 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.009504 LAYER D6 ;
      ANTENNAMAXAREACAR 41.8661 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 97.9577 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.4655 0 32.5455 0.08 ;
    END
  END CsrTxStren120Pd[0]
  PIN CsrTxOdtStren480Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 61.7226 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 158.802 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 27.6305 0 27.7105 0.08 ;
    END
  END CsrTxOdtStren480Pu
  PIN CsrTxOdtStren480Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 58.0544 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 144.663 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 30.2105 0 30.2905 0.08 ;
    END
  END CsrTxOdtStren480Pd
  PIN CsrTxOdtStren240Pu
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 61.7226 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 158.802 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 26.4305 0 26.5105 0.08 ;
    END
  END CsrTxOdtStren240Pu
  PIN CsrTxOdtStren240Pd
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 58.0544 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 144.663 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 31.4105 0 31.4905 0.08 ;
    END
  END CsrTxOdtStren240Pd
  PIN CsrTxOdtStren120Pu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 61.7226 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 158.802 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 21.6305 0 21.7105 0.08 ;
    END
  END CsrTxOdtStren120Pu[3]
  PIN CsrTxOdtStren120Pu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 61.7226 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 158.802 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 22.8305 0 22.9105 0.08 ;
    END
  END CsrTxOdtStren120Pu[2]
  PIN CsrTxOdtStren120Pu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 61.7226 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 158.802 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 24.0305 0 24.1105 0.08 ;
    END
  END CsrTxOdtStren120Pu[1]
  PIN CsrTxOdtStren120Pu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 61.7226 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 158.802 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 25.2305 0 25.3105 0.08 ;
    END
  END CsrTxOdtStren120Pu[0]
  PIN CsrTxOdtStren120Pd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 58.0544 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 144.663 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 36.2105 0 36.2905 0.08 ;
    END
  END CsrTxOdtStren120Pd[3]
  PIN CsrTxOdtStren120Pd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 58.0544 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 144.663 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 35.0105 0 35.0905 0.08 ;
    END
  END CsrTxOdtStren120Pd[2]
  PIN CsrTxOdtStren120Pd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 58.0544 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 144.663 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.8105 0 33.8905 0.08 ;
    END
  END CsrTxOdtStren120Pd[1]
  PIN CsrTxOdtStren120Pd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.19432 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45162 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.005184 LAYER D6 ;
      ANTENNAMAXAREACAR 58.0544 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 144.663 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.6105 0 32.6905 0.08 ;
    END
  END CsrTxOdtStren120Pd[0]
  PIN CsrReserved[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.17272 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40302 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 159.25 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 407.778 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 33.1555 0 33.2355 0.08 ;
    END
  END CsrReserved[2]
  PIN CsrReserved[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.17272 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40302 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 171.083 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 448.444 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.3205 0 32.4005 0.08 ;
    END
  END CsrReserved[1]
  PIN CsrReserved[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.17272 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.40302 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D6 ;
      ANTENNAMAXAREACAR 171.05 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 448.139 LAYER D6 ;
    PORT
      LAYER D6 ;
        RECT 32.082 0 32.162 0.08 ;
    END
  END CsrReserved[0]
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER D8 ;
        RECT 0.6 28.98 37.98 29.68 ;
        RECT 0.6 26.86 37.98 27.56 ;
        RECT 0.6 24.74 37.98 25.44 ;
        RECT 0.6 22.62 37.98 23.32 ;
        RECT 0.6 20.5 37.98 21.2 ;
        RECT 0.6 18.38 37.98 19.08 ;
        RECT 0.6 16.26 37.98 16.96 ;
        RECT 0.6 14.14 37.98 14.84 ;
        RECT 0.6 12.02 37.98 12.72 ;
        RECT 0.6 9.9 37.98 10.6 ;
        RECT 0.6 7.78 37.98 8.48 ;
        RECT 0.6 5.66 37.98 6.36 ;
        RECT 0.6 3.54 37.98 4.24 ;
        RECT 0.6 1.42 37.98 2.12 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 198.49025 37.98 199.29025 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.633 226.576 35.583 227.276 ;
        RECT 2.633 224.014 35.583 224.714 ;
        RECT 2.633 221.452 35.583 222.152 ;
        RECT 2.633 218.89 35.583 219.59 ;
        RECT 2.633 216.328 35.583 217.028 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 191.83825 37.98 192.63825 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 174.84125 37.98 175.64125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.36625 212.673 37.98 213.073 ;
        RECT 0.36625 207.513 37.98 207.913 ;
        RECT 0.36625 205.968 37.98 206.368 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 177.44125 37.98 178.24125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 172.24125 37.98 173.04125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 189.23825 37.9805 190.03825 ;
        RECT 0.607 186.63825 37.9805 187.43825 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.58675 180.04125 37.98 180.84125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 154.14575 37.98 154.94575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 156.54575 37.98 157.34575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 163.04575 37.98 163.84575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 160.44575 37.98 161.24575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 167.04125 37.98 167.84125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 150.24575 37.98 151.04575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.58675 135.812 37.98 136.612 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 133.212 37.98 134.012 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 142.44575 37.98 143.24575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 141.012 37.98 141.812 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 145.04575 37.98 145.84575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 147.64575 37.98 148.44575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 125.412 37.98 126.212 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 122.6965 37.98 123.4965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 116.2965 37.98 117.0965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 130.612 37.98 131.412 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 109.8965 37.98 110.6965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 103.9965 37.98 104.7965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 90.35925 18.1835 91.15925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 83.8965 37.98 84.6965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 86.4965 37.98 87.2965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.55475 81.2965 37.98 82.0965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 41.618 37.98 42.418 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 44.218 37.98 45.018 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 32.518 37.98 33.318 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 34.818 37.98 35.618 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.15275 112.4965 37.98 113.2965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 105.0965 17.4185 105.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 102.4965 17.4185 103.2965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 108.4965 17.4185 109.2965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 111.0965 17.4185 111.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 113.6965 17.4185 114.4965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 100.4965 37.98 101.2965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 94.4965 37.98 95.2965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 97.0965 37.98 97.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 98.15925 18.1835 98.95925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 95.55925 18.1835 96.35925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 92.95925 18.1835 93.75925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.55475 79.0965 18.383 79.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 69.3965 37.98 70.1965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 67.1965 37.98 67.9965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 64.9965 37.98 65.7965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 71.9965 37.98 72.7965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5885 63.8965 18.25175 64.6965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5885 56.718 18.25175 57.518 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 59.118 37.98 59.918 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 54.318 37.98 55.118 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 48.818 37.98 49.618 ;
    END
    PORT
      LAYER D8 ;
        RECT 18.64375 38.118 37.98 38.918 ;
    END
  END VSS
  PIN VSH
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 421.175 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 100.526 LAYER D8 ;
    ANTENNADIFFAREA 57.9223 LAYER D8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 7.4132 LAYER D8 ;
      ANTENNAMAXAREACAR 298.228 LAYER D8 ;
      ANTENNAMAXSIDEAREACAR 241.957 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 0.6 199.91925 37.98 200.71925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 195.85025 37.98 196.65025 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6075 170.94125 37.98 171.74125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.58725 185.33825 37.98 186.13825 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.36625 214.353 37.98 214.753 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 165.74125 37.98 166.54125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.58675 152.84575 37.98 153.64575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.58675 117.4965 37.98 118.2965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 128.012 37.98 128.812 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16475 106.1965 37.98 106.9965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 46.618 37.98 47.418 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 90.9965 37.98 91.7965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.01925 73.746 37.98 74.546 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 68.2965 37.98 69.0965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.55475 77.9965 37.98 78.7965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 53.218 37.98 54.018 ;
    END
    PORT
      LAYER D8 ;
        RECT 17.054 61.6965 37.98 62.4965 ;
    END
  END VSH
  PIN VIO_TIE_LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.35572 LAYER D6 ;
    ANTENNAPARTIALMETALAREA 0.58526 LAYER D7 ;
    ANTENNAPARTIALMETALAREA 0.0576 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4582999375 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.64087 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0864 LAYER D8 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S6 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S7 ;
    ANTENNADIFFAREA 0.16128 LAYER D7 ;
    ANTENNADIFFAREA 0.16128 LAYER S7 ;
    ANTENNADIFFAREA 0.16128 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 19.51 207.168 19.75 207.408 ;
    END
    PORT
      LAYER D6 ;
        RECT 23.307 201.57775 23.407 215.135 ;
    END
  END VIO_TIE_LO
  PIN VIO_TIE_HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.35572 LAYER D6 ;
    ANTENNAPARTIALMETALAREA 0.61246 LAYER D7 ;
    ANTENNAPARTIALMETALAREA 0.0576 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4582999375 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.76327 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0864 LAYER D8 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S6 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S7 ;
    ANTENNADIFFAREA 0.16128 LAYER D7 ;
    ANTENNADIFFAREA 0.16128 LAYER S7 ;
    ANTENNADIFFAREA 0.16128 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 18.83 207.168 19.07 207.408 ;
    END
    PORT
      LAYER D6 ;
        RECT 23.007 201.57775 23.107 215.135 ;
    END
  END VIO_TIE_HI
  PIN VIO_PwrOk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.552 LAYER D5 ;
    ANTENNAPARTIALMETALAREA 15.2815 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 6.8328 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2205 LAYER D6 ;
    ANTENNAPARTIALCUTAREA 0.0064 LAYER S5 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2016 LAYER D5 ;
      ANTENNAGATEAREA 0.2016 LAYER S5 ;
      ANTENNAGATEAREA 0.2016 LAYER D6 ;
      ANTENNAMAXAREACAR 48.9421 LAYER D5 ;
      ANTENNAMAXAREACAR 124.743 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 38.9363 LAYER D5 ;
      ANTENNAMAXSIDEAREACAR 124.355 LAYER D6 ;
      ANTENNAMAXCUTCAR 0.0688095625 LAYER S5 ;
    PORT
      LAYER D5 ;
        RECT 0 125.044 0.2 125.244 ;
    END
    PORT
      LAYER D5 ;
        RECT 0.2 29.734 37.96 29.934 ;
    END
  END VIO_PwrOk
  PIN VIO_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.674 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 2.82132 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 2.165 237.86 35.995 238.88 ;
        RECT 2.165 235.298 35.995 236.318 ;
        RECT 2.165 232.736 35.995 233.756 ;
        RECT 2.165 230.174 35.995 231.194 ;
        RECT 2.633 225.134 35.583 226.154 ;
        RECT 2.633 220.01 35.583 221.03 ;
        RECT 2.633 217.448 35.583 218.468 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 182.78925 17.012 183.78925 ;
    END
    PORT
      LAYER D8 ;
        RECT 21.4975 182.78925 36.1715 183.78925 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.633 222.572 35.583 223.592 ;
    END
    PORT
      LAYER D8 ;
        RECT 21.4975 158.50475 36.1715 159.50475 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 158.50475 17.012 159.50475 ;
    END
    PORT
      LAYER D8 ;
        RECT 21.4975 139.548 36.1715 140.548 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 139.548 17.012 140.548 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 120.68075 17.012 121.68075 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 106.49275 17.012 107.49275 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 87.8805 17.012 88.8805 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 73.646 17.012 74.646 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 52.684 17.012 53.684 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.338 38.438 17.012 39.438 ;
    END
  END VIO_PAD
  PIN VIO_FuncMode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2016 LAYER D7 ;
      ANTENNAMAXAREACAR 9.99107 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 41.3104 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.413 37.98 208.453 ;
    END
  END VIO_FuncMode
  PIN VIO_ForceLow
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.35842 LAYER D6 ;
    ANTENNAPARTIALMETALAREA 0.73307 LAYER D7 ;
    ANTENNAPARTIALMETALAREA 0.0576 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 2.46317 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.30601 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0864 LAYER D8 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S6 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2016 LAYER D7 ;
      ANTENNAGATEAREA 0.2016 LAYER S7 ;
      ANTENNAGATEAREA 0.2016 LAYER D8 ;
      ANTENNAMAXAREACAR 4.31673 LAYER D7 ;
      ANTENNAMAXAREACAR 4.60244 LAYER D8 ;
      ANTENNAMAXSIDEAREACAR 19.044 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 19.4726 LAYER D8 ;
      ANTENNAMAXCUTCAR 0.0536706875 LAYER S7 ;
    PORT
      LAYER D8 ;
        RECT 19.17 207.168 19.41 207.408 ;
    END
    PORT
      LAYER D6 ;
        RECT 9.59575 201.57775 9.69575 215.135 ;
    END
  END VIO_ForceLow
  PIN VIO_CsrTxThermP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.9886 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 75.7048 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 210.453 37.98 210.493 ;
    END
  END VIO_CsrTxThermP[9]
  PIN VIO_CsrTxThermP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.6413 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 73.360299938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 209.773 37.98 209.813 ;
    END
  END VIO_CsrTxThermP[8]
  PIN VIO_CsrTxThermP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.48 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 73.6287 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 209.693 37.98 209.733 ;
    END
  END VIO_CsrTxThermP[7]
  PIN VIO_CsrTxThermP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.0498 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 71.7502 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 209.053 37.98 209.093 ;
    END
  END VIO_CsrTxThermP[6]
  PIN VIO_CsrTxThermP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.0117 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 71.4979 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.973 37.98 209.013 ;
    END
  END VIO_CsrTxThermP[5]
  PIN VIO_CsrTxThermP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 15.959 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 71.2746 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.893 37.98 208.933 ;
    END
  END VIO_CsrTxThermP[4]
  PIN VIO_CsrTxThermP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 15.8158 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 70.5146 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.813 37.98 208.853 ;
    END
  END VIO_CsrTxThermP[3]
  PIN VIO_CsrTxThermP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.8432 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.8643 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.253 37.98 213.293 ;
    END
  END VIO_CsrTxThermP[30]
  PIN VIO_CsrTxThermP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 15.8375 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 70.3139 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.733 37.98 208.773 ;
    END
  END VIO_CsrTxThermP[2]
  PIN VIO_CsrTxThermP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.6724 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.0843 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.173 37.98 213.213 ;
    END
  END VIO_CsrTxThermP[29]
  PIN VIO_CsrTxThermP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.3055 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 77.3435 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 212.533 37.98 212.573 ;
    END
  END VIO_CsrTxThermP[28]
  PIN VIO_CsrTxThermP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.1745 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 76.5399 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 212.453 37.98 212.493 ;
    END
  END VIO_CsrTxThermP[27]
  PIN VIO_CsrTxThermP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.239899937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 75.8925 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 212.373 37.98 212.413 ;
    END
  END VIO_CsrTxThermP[26]
  PIN VIO_CsrTxThermP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.0168 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 75.2171 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 212.293 37.98 212.333 ;
    END
  END VIO_CsrTxThermP[25]
  PIN VIO_CsrTxThermP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.2415 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 81.3662 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 212.213 37.98 212.253 ;
    END
  END VIO_CsrTxThermP[24]
  PIN VIO_CsrTxThermP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.228 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 81.3772 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 212.133 37.98 212.173 ;
    END
  END VIO_CsrTxThermP[23]
  PIN VIO_CsrTxThermP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.1753 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.9847 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 212.053 37.98 212.093 ;
    END
  END VIO_CsrTxThermP[22]
  PIN VIO_CsrTxThermP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.2984 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 80.4418 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 211.973 37.98 212.013 ;
    END
  END VIO_CsrTxThermP[21]
  PIN VIO_CsrTxThermP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.4544 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 77.754599938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 211.893 37.98 211.933 ;
    END
  END VIO_CsrTxThermP[20]
  PIN VIO_CsrTxThermP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 15.6468 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 69.6243 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.653 37.98 208.693 ;
    END
  END VIO_CsrTxThermP[1]
  PIN VIO_CsrTxThermP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 18.0657 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 80.650099938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 211.813 37.98 211.853 ;
    END
  END VIO_CsrTxThermP[19]
  PIN VIO_CsrTxThermP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.9482 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 80.2359 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 211.733 37.98 211.773 ;
    END
  END VIO_CsrTxThermP[18]
  PIN VIO_CsrTxThermP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.8617 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.974599938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 211.653 37.98 211.693 ;
    END
  END VIO_CsrTxThermP[17]
  PIN VIO_CsrTxThermP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.684 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 79.1491 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 211.573 37.98 211.613 ;
    END
  END VIO_CsrTxThermP[16]
  PIN VIO_CsrTxThermP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.6546 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 78.9312 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 211.493 37.98 211.533 ;
    END
  END VIO_CsrTxThermP[15]
  PIN VIO_CsrTxThermP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.5681 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 78.427599938 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 211.413 37.98 211.453 ;
    END
  END VIO_CsrTxThermP[14]
  PIN VIO_CsrTxThermP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.2723 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 76.9923 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 210.773 37.98 210.813 ;
    END
  END VIO_CsrTxThermP[13]
  PIN VIO_CsrTxThermP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.2026 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 76.5698 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 210.693 37.98 210.733 ;
    END
  END VIO_CsrTxThermP[12]
  PIN VIO_CsrTxThermP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.126899937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 76.0991 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 210.613 37.98 210.653 ;
    END
  END VIO_CsrTxThermP[11]
  PIN VIO_CsrTxThermP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 17.1565 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 76.3459 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 210.533 37.98 210.573 ;
    END
  END VIO_CsrTxThermP[10]
  PIN VIO_CsrTxThermP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 15.7299 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 69.6262 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.573 37.98 208.613 ;
    END
  END VIO_CsrTxThermP[0]
  PIN VIO_CsrTxCalBaseP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.564699937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 73.3582 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.253 37.98 208.293 ;
    END
  END VIO_CsrTxCalBaseP
  PIN VIO_CsrPreDriveMode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.302099937 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 72.2795 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.493 37.98 208.533 ;
    END
  END VIO_CsrPreDriveMode[2]
  PIN VIO_CsrPreDriveMode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1008 LAYER D7 ;
      ANTENNAMAXAREACAR 16.349 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 72.376 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.333 37.98 208.373 ;
    END
  END VIO_CsrPreDriveMode[1]
  PIN VIO_CsrPreDriveMode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3024 LAYER D7 ;
      ANTENNAMAXAREACAR 6.2087199375 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 24.8596 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.173 37.98 208.213 ;
    END
  END VIO_CsrPreDriveMode[0]
  PIN VDS3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.0779 LAYER D8 ;
    ANTENNAPARTIALMETALSIDEAREA 7.00596 LAYER D8 ;
    ANTENNADIFFAREA 2.96654 LAYER D8 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.628992 LAYER D8 ;
      ANTENNAMAXAREACAR 373.687 LAYER D8 ;
      ANTENNAMAXSIDEAREACAR 131.142 LAYER D8 ;
    PORT
      LAYER D8 ;
        RECT 0 240.888 38.16 241.65 ;
    END
  END VDS3
  PIN VDDQ
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER D8 ;
        RECT 0.607 190.53825 37.98 191.33825 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5885 37.018 18.25175 37.818 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5885 33.618 18.25175 34.418 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5885 31.418 18.25175 32.218 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 193.13825 37.98 193.93825 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 201.21925 37.98 202.01925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 176.14125 37.98 176.94125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 178.74125 37.98 179.54125 ;
    END
    PORT
      LAYER D8 ;
        RECT 2.165 239.302 35.995 240.002 ;
        RECT 2.165 236.74 35.995 237.44 ;
        RECT 2.165 234.178 35.995 234.878 ;
        RECT 2.165 231.616 35.995 232.316 ;
        RECT 2.165 229.054 35.995 229.754 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 187.93825 37.9805 188.73825 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 173.54125 37.98 174.34125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 181.34125 37.98 182.14125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.36625 210.913 37.98 211.313 ;
        RECT 0.36625 209.193 37.98 209.593 ;
        RECT 0.36625 204.608 37.98 205.008 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.36625 206.688 37.98 207.068 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 155.24575 37.98 156.04575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 161.74575 37.98 162.54575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 164.44125 37.98 165.24125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 151.54575 37.98 152.34575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 131.912 37.98 132.712 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 134.512 37.98 135.312 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 137.112 37.98 137.912 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 146.34575 37.98 147.14575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 143.74575 37.98 144.54575 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 148.94575 37.98 149.74575 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16175 120.78075 37.98 121.58075 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 123.9965 19.46575 124.7965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 126.712 19.46575 127.512 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 118.7965 37.98 119.5965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 129.312 37.98 130.112 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.527 114.9965 37.98 115.7965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 102.6965 37.98 103.4965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 108.5965 37.98 109.3965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 27.92 37.98 28.62 ;
        RECT 0.6 25.8 37.98 26.5 ;
        RECT 0.6 23.68 37.98 24.38 ;
        RECT 0.6 21.56 37.98 22.26 ;
        RECT 0.6 17.32 37.98 18.02 ;
        RECT 0.6 13.08 37.98 13.78 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 85.1965 37.98 85.9965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5095 82.5965 37.98 83.3965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 40.318 37.98 41.118 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 45.518 37.98 46.318 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 42.918 37.98 43.718 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 35.918 37.98 36.718 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 30.318 37.98 31.118 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.15275 111.1965 37.98 111.9965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 109.7965 17.4185 110.5965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 103.7965 17.4185 104.5965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 112.3965 17.4185 113.1965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 99.3965 37.98 100.1965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 93.1965 37.98 93.9965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 88.7965 37.98 89.5965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 95.7965 37.98 96.5965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 96.85925 16.623 97.65925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 94.25925 16.623 95.05925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 91.65925 18.1835 92.45925 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 75.7965 16.623 76.5965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 66.0965 16.623 66.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 76.8965 37.98 77.6965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 70.6965 37.98 71.4965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.55475 80.1965 37.98 80.9965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5885 61.6965 16.6115 62.4965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5885 49.918 18.25175 50.718 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5885 47.718 18.25175 48.518 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 60.418 37.98 61.218 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 55.618 37.98 56.418 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 57.818 37.98 58.618 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 51.018 37.98 51.818 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.5995 62.7965 37.98 63.5965 ;
    END
  END VDDQ
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER D8 ;
        RECT 25.1005 4.6 37.98 5.3 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 197.19025 37.98 197.99025 ;
        RECT 0.607 194.55025 37.98 195.35025 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.36625 209.953 37.98 210.353 ;
        RECT 0.36625 203.848 37.98 204.248 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 168.34125 37.98 169.14125 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.607 169.64125 37.98 170.44125 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.8195 123.9965 37.986 124.7965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.8195 126.712 37.986 127.512 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16475 105.0965 37.98 105.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 107.4965 37.98 108.2965 ;
    END
    PORT
      LAYER D8 ;
        RECT 0.6 19.44 37.98 20.14 ;
        RECT 0.6 15.2 37.98 15.9 ;
        RECT 0.6 10.96 37.98 11.66 ;
        RECT 0.6 8.84 37.98 9.54 ;
        RECT 0.6 6.72 37.98 7.42 ;
        RECT 0.6 2.48 37.98 3.18 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 101.5965 37.98 102.3965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 113.6965 37.98 114.4965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 75.7965 37.98 76.5965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 87.6965 37.98 88.4965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 92.0965 37.98 92.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 89.8965 37.98 90.6965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 98.2965 37.98 99.0965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 79.0965 37.98 79.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 66.0965 37.98 66.8965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 56.718 37.98 57.518 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 47.718 37.98 48.518 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 49.918 37.98 50.718 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 52.118 37.98 52.918 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 63.8965 37.98 64.6965 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 33.718 37.98 34.518 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 37.018 37.98 37.818 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 31.418 37.98 32.218 ;
    END
    PORT
      LAYER D8 ;
        RECT 19.16125 39.218 37.98 40.018 ;
    END
  END VDD
  PIN TIE_LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.88785 LAYER D5 ;
    ANTENNAPARTIALMETALAREA 4.77515 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8350649375 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8529 LAYER D6 ;
    ANTENNAPARTIALCUTAREA 0.0064 LAYER S5 ;
    ANTENNADIFFAREA 0.016848 LAYER D6 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.559872 LAYER D6 ;
      ANTENNAMAXAREACAR 48.1036 LAYER D6 ;
      ANTENNAMAXSIDEAREACAR 99.5868 LAYER D6 ;
    PORT
      LAYER D5 ;
        RECT 20.887 201.876 24.09025 202.076 ;
    END
    PORT
      LAYER D6 ;
        RECT 23.607 201.57775 23.707 215.135 ;
    END
  END TIE_LO
  PIN TIE_HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5552999375 LAYER D5 ;
    ANTENNAPARTIALMETALAREA 1.35572 LAYER D6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.23577 LAYER D5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4582999375 LAYER D6 ;
    ANTENNAPARTIALCUTAREA 0.0032 LAYER S5 ;
    ANTENNADIFFAREA 0.008424 LAYER D5 ;
    ANTENNADIFFAREA 0.008424 LAYER S5 ;
    ANTENNADIFFAREA 0.008424 LAYER D6 ;
    PORT
      LAYER D5 ;
        RECT 20.967 214.321 24.09025 214.521 ;
    END
    PORT
      LAYER D6 ;
        RECT 23.833 201.57775 23.933 215.135 ;
    END
  END TIE_HI
  PIN CsrTxThermN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1313.56 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5769.15 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.708 37.98 203.748 ;
    END
  END CsrTxThermN[9]
  PIN CsrTxThermN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1290.28 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5671.1 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.628 37.98 203.668 ;
    END
  END CsrTxThermN[8]
  PIN CsrTxThermN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1250.67 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5624.81 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.548 37.98 203.588 ;
    END
  END CsrTxThermN[7]
  PIN CsrTxThermN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1254.8 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5628.94 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.468 37.98 203.508 ;
    END
  END CsrTxThermN[6]
  PIN CsrTxThermN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1257.85 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5552.72 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.388 37.98 203.428 ;
    END
  END CsrTxThermN[5]
  PIN CsrTxThermN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1266.2 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5684.67 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.308 37.98 203.348 ;
    END
  END CsrTxThermN[4]
  PIN CsrTxThermN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1253.81 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5630.41 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.228 37.98 203.268 ;
    END
  END CsrTxThermN[3]
  PIN CsrTxThermN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1240.23 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5557.29 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 206.548 37.98 206.588 ;
    END
  END CsrTxThermN[30]
  PIN CsrTxThermN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1282.48 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5715.32 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.148 37.98 203.188 ;
    END
  END CsrTxThermN[2]
  PIN CsrTxThermN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1234.37 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5553.33 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 206.468 37.98 206.508 ;
    END
  END CsrTxThermN[29]
  PIN CsrTxThermN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1255.38 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5591.4 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.828 37.98 205.868 ;
    END
  END CsrTxThermN[28]
  PIN CsrTxThermN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1255.87 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5586.74 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.748 37.98 205.788 ;
    END
  END CsrTxThermN[27]
  PIN CsrTxThermN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1267.33 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5624.33 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.668 37.98 205.708 ;
    END
  END CsrTxThermN[26]
  PIN CsrTxThermN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1268.73 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5623.59 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.588 37.98 205.628 ;
    END
  END CsrTxThermN[25]
  PIN CsrTxThermN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1190.63 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5338.32 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.508 37.98 205.548 ;
    END
  END CsrTxThermN[24]
  PIN CsrTxThermN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1246.29 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5574.01 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.428 37.98 205.468 ;
    END
  END CsrTxThermN[23]
  PIN CsrTxThermN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1234.9 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5501.39 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.348 37.98 205.388 ;
    END
  END CsrTxThermN[22]
  PIN CsrTxThermN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1255.59 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5596.73 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.268 37.98 205.308 ;
    END
  END CsrTxThermN[21]
  PIN CsrTxThermN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1248.69 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5586.55 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.188 37.98 205.228 ;
    END
  END CsrTxThermN[20]
  PIN CsrTxThermN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1235.58 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5523.36 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 203.068 37.98 203.108 ;
    END
  END CsrTxThermN[1]
  PIN CsrTxThermN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1243.39 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5576.03 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 205.108 37.98 205.148 ;
    END
  END CsrTxThermN[19]
  PIN CsrTxThermN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1249.13 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5600.45 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 204.428 37.98 204.468 ;
    END
  END CsrTxThermN[18]
  PIN CsrTxThermN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1239.38 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5535.29 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 204.348 37.98 204.388 ;
    END
  END CsrTxThermN[17]
  PIN CsrTxThermN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1334.51 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5967.73 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.093 37.98 208.133 ;
    END
  END CsrTxThermN[16]
  PIN CsrTxThermN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1274.83 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5674.29 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 208.013 37.98 208.053 ;
    END
  END CsrTxThermN[15]
  PIN CsrTxThermN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1344.18 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5792.53 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 202.588 37.98 202.628 ;
    END
  END CsrTxThermN[14]
  PIN CsrTxThermN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1317.88 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5745.13 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 202.668 37.98 202.708 ;
    END
  END CsrTxThermN[13]
  PIN CsrTxThermN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1336.12 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5807.04 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 202.748 37.98 202.788 ;
    END
  END CsrTxThermN[12]
  PIN CsrTxThermN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1302.79 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5665.07 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 202.828 37.98 202.868 ;
    END
  END CsrTxThermN[11]
  PIN CsrTxThermN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1325.72 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5781.6 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 202.908 37.98 202.948 ;
    END
  END CsrTxThermN[10]
  PIN CsrTxThermN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.001296 LAYER D7 ;
      ANTENNAMAXAREACAR 1275.9 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 5725.6 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 202.988 37.98 203.028 ;
    END
  END CsrTxThermN[0]
  PIN CsrTxSrc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 607.474 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2727.88 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 214.213 37.98 214.253 ;
    END
  END CsrTxSrc[7]
  PIN CsrTxSrc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 609.986 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2732.4 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 214.133 37.98 214.173 ;
    END
  END CsrTxSrc[6]
  PIN CsrTxSrc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 614.607 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2756.36 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 214.053 37.98 214.093 ;
    END
  END CsrTxSrc[5]
  PIN CsrTxSrc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 612.189 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2748.18 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.973 37.98 214.013 ;
    END
  END CsrTxSrc[4]
  PIN CsrTxSrc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 602.723 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2706.22 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.893 37.98 213.933 ;
    END
  END CsrTxSrc[3]
  PIN CsrTxSrc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 600.451 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2690.58 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.733 37.98 213.773 ;
    END
  END CsrTxSrc[2]
  PIN CsrTxSrc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 608.51 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2731.15 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.573 37.98 213.613 ;
    END
  END CsrTxSrc[1]
  PIN CsrTxSrc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4952 LAYER D7 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7355999375 LAYER D7 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.002592 LAYER D7 ;
      ANTENNAMAXAREACAR 596.955 LAYER D7 ;
      ANTENNAMAXSIDEAREACAR 2677.3 LAYER D7 ;
    PORT
      LAYER D7 ;
        RECT 0.6 213.413 37.98 213.453 ;
    END
  END CsrTxSrc[0]
  OBS
    LAYER M1 SPACING 0 ;
      RECT 0 0 38.16 241.65 ;
    LAYER M2 SPACING 0 ;
      RECT 0 0 38.16 241.65 ;
    LAYER M3 SPACING 0 ;
      RECT 0 0 38.16 241.65 ;
    LAYER M4 SPACING 0 ;
      RECT 0 0 38.16 241.65 ;
      RECT MASK 1 10.48325 205.5215 10.53125 211.595 ;
    LAYER D5 SPACING 0 ;
      RECT 0 0 38.16 29.634 ;
      POLYGON 0 30.034 0 125.044 0.2 125.044 0.2 125.244 0 125.244 0 241.65 38.16 241.65 38.16 214.521 20.967 214.521 20.967 214.321 24.09025 214.321 24.09025 214.521 38.16 214.521 38.16 202.076 20.887 202.076 20.887 201.876 24.09025 201.876 24.09025 202.076 38.16 202.076 38.16 30.034 ;
    LAYER D6 SPACING 0 ;
      POLYGON 0 0 0 241.65 38.16 241.65 38.16 215.135 9.59575 215.135 9.59575 201.57775 9.69575 201.57775 9.69575 215.135 23.007 215.135 23.007 201.57775 23.107 201.57775 23.107 215.135 23.307 215.135 23.307 201.57775 23.407 201.57775 23.407 215.135 23.607 215.135 23.607 201.57775 23.707 201.57775 23.707 215.135 23.833 215.135 23.833 201.57775 23.933 201.57775 23.933 215.135 38.16 215.135 38.16 0 36.2905 0 36.2905 0.08 36.2105 0.08 36.2105 0 36.1455 0 36.1455 0.08 36.0655 0.08 36.0655 0 35.4905 0 35.4905 0.08 35.4105 0.08 35.4105 0 35.3455 0 35.3455 0.08 35.2655 0.08 35.2655 0 35.0905 0 35.0905 0.08 35.0105 0.08 35.0105 0 34.9455 0 34.9455 0.08 34.8655 0.08 34.8655 0 34.2905 0 34.2905 0.08 34.2105 0.08 34.2105 0 34.1455 0 34.1455 0.08 34.0655 0.08 34.0655 0 33.8905 0 33.8905 0.08 33.8105 0.08 33.8105 0 33.7455 0 33.7455 0.08 33.6655 0.08 33.6655 0 33.2355 0 33.2355 0.08 33.1555 0.08 33.1555 0 33.0905 0 33.0905 0.08 33.0105 0.08 33.0105 0 32.9455 0 32.9455 0.08 32.8655 0.08 32.8655 0 32.6905 0 32.6905 0.08 32.6105 0.08 32.6105 0 32.5455 0 32.5455 0.08 32.4655 0.08 32.4655 0 32.4005 0 32.4005 0.08 32.3205 0.08 32.3205 0 32.162 0 32.162 0.08 32.082 0.08 32.082 0 31.8905 0 31.8905 0.08 31.8105 0.08 31.8105 0 31.7455 0 31.7455 0.08 31.6655 0.08 31.6655 0 31.4905 0 31.4905 0.08 31.4105 0.08 31.4105 0 31.3455 0 31.3455 0.08 31.2655 0.08 31.2655 0 30.6905 0 30.6905 0.08 30.6105 0.08 30.6105 0 30.5455 0 30.5455 0.08 30.4655 0.08 30.4655 0 30.2905 0 30.2905 0.08 30.2105 0.08 30.2105 0 30.1455 0 30.1455 0.08 30.0655 0.08 30.0655 0 29.4905 0 29.4905 0.08 29.4105 0.08 29.4105 0 29.3455 0 29.3455 0.08 29.2655 0.08 29.2655 0 29.2005 0 29.2005 0.08 29.1205 0.08 29.1205 0 29.0555 0 29.0555 0.08 28.9755 0.08 28.9755 0 28.9105 0 28.9105 0.08 28.8305 0.08 28.8305 0 28.7655 0 28.7655 0.08 28.6855 0.08 28.6855 0 28.2905 0 28.2905 0.08 28.2105 0.08 28.2105 0 28.1455 0 28.1455 0.08 28.0655 0.08 28.0655 0 28.0005 0 28.0005 0.08 27.9205 0.08 27.9205 0 27.8555 0 27.8555 0.08 27.7755 0.08 27.7755 0 27.7105 0 27.7105 0.08 27.6305 0.08 27.6305 0 27.5655 0 27.5655 0.08 27.4855 0.08 27.4855 0 27.0555 0 27.0555 0.08 26.9755 0.08 26.9755 0 26.9105 0 26.9105 0.08 26.8305 0.08 26.8305 0 26.7655 0 26.7655 0.08 26.6855 0.08 26.6855 0 26.5105 0 26.5105 0.08 26.4305 0.08 26.4305 0 26.3655 0 26.3655 0.08 26.2855 0.08 26.2855 0 25.8555 0 25.8555 0.08 25.7755 0.08 25.7755 0 25.7105 0 25.7105 0.08 25.6305 0.08 25.6305 0 25.5655 0 25.5655 0.08 25.4855 0.08 25.4855 0 25.3105 0 25.3105 0.08 25.2305 0.08 25.2305 0 25.1655 0 25.1655 0.08 25.0855 0.08 25.0855 0 24.6555 0 24.6555 0.08 24.5755 0.08 24.5755 0 24.5105 0 24.5105 0.08 24.4305 0.08 24.4305 0 24.3655 0 24.3655 0.08 24.2855 0.08 24.2855 0 24.1105 0 24.1105 0.08 24.0305 0.08 24.0305 0 23.9655 0 23.9655 0.08 23.8855 0.08 23.8855 0 23.3105 0 23.3105 0.08 23.2305 0.08 23.2305 0 23.1655 0 23.1655 0.08 23.0855 0.08 23.0855 0 22.9105 0 22.9105 0.08 22.8305 0.08 22.8305 0 22.7655 0 22.7655 0.08 22.6855 0.08 22.6855 0 22.1105 0 22.1105 0.08 22.0305 0.08 22.0305 0 21.9655 0 21.9655 0.08 21.8855 0.08 21.8855 0 21.7105 0 21.7105 0.08 21.6305 0.08 21.6305 0 21.5655 0 21.5655 0.08 21.4855 0.08 21.4855 0 20.9105 0 20.9105 0.08 20.8305 0.08 20.8305 0 20.7655 0 20.7655 0.08 20.6855 0.08 20.6855 0 20.4755 0 20.4755 0.08 20.3955 0.08 20.3955 0 20.3305 0 20.3305 0.08 20.2505 0.08 20.2505 0 18.59425 0 18.59425 0.32625 18.19425 0.32625 18.19425 0 7.696 0 7.696 0.08 7.616 0.08 7.616 0 2.9735 0 2.9735 0.08 2.8935 0.08 2.8935 0 2.8285 0 2.8285 0.08 2.7485 0.08 2.7485 0 2.6835 0 2.6835 0.08 2.6035 0.08 2.6035 0 2.5385 0 2.5385 0.08 2.4585 0.08 2.4585 0 2.3935 0 2.3935 0.08 2.3135 0.08 2.3135 0 ;
    LAYER D7 SPACING 0 ;
      RECT 0 0 38.16 202.308 ;
      RECT 0.6 203.848 37.98 204.248 ;
      RECT 0.6 204.608 37.98 205.008 ;
      RECT 0.6 205.968 37.98 206.368 ;
      RECT 0.6 206.688 37.98 207.068 ;
      RECT 1.08325 207.228 19.41 207.268 ;
      RECT 19.51 207.228 34.1415 207.268 ;
      RECT 18.83 207.308 34.1415 207.348 ;
      RECT 0.6 207.513 37.98 207.913 ;
      RECT 0.6 209.193 37.98 209.593 ;
      RECT 0.6 209.953 37.98 210.353 ;
      RECT 0.6 210.913 37.98 211.313 ;
      RECT 0.6 212.673 37.98 213.073 ;
      RECT 0 214.353 38.16 214.753 ;
      RECT 0 215.135 38.16 241.65 ;
  END
END dwc_ddrphy_txrxac_ns

END LIBRARY
